`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lEAWhwyix5jBGG66vdOS8nJpVNdFrJkI8qYgE8UK5+7avncLp8v54uPGoRWR36jLWh6ehDkiSjec
BS6Kf+NkuQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pIREr1/dqaPvd4j2lTxOBSnAy2Ra6DuJsnP63kEHv0IS6up5E7T2izznuVUSTCTOb47ap4dcNzFs
VunReb3wPh7pLPeb7xw5iV9uBkd/TpxZM73yc3k1Rpf+4J2IVlTVOAQ5OEjaorVixNlt8NiWGqzH
R/d96oqeazauoI3oOnQ=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DELvK5o++4pE4MCoxr5fui0H5JI8L1lrkSphbogK2GjTRYuCaX9esyobvkVAA3D3d9tJqaP3hGDO
abwxN4b4ezNtusv1gy6cglGx/GN3jUuKSbgskyfUxDvL7LrGyqNFVNMUu2E9m+BfM4Ntpn0n9FIV
ziDzomLe9jJOEfua5U0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V5WVwaxzoZCaNjBtQkebL2emEOYwtLrt2YC/Nhjv+maBGQv/B4iXQaCQdVt72XysdOqpG+W7acY4
LQoDKOXjpn3NnQIeXe5yNHpeBxy0UeQS9x3LKwyD7PTy2e6Psu8FyrhI0YZfF7izMLFdHz6hGOSF
AIMgUa/N0UmNtXEjM3DkfZLqoYQAht0o6JFtiqajvc59tPsvMZCCtiKwhXu7PlN11ghLauG7TulD
K2KfLDkX0cfwDA2TPyp16kT6EIfZoCRnafITvpKhHXZv+NQc+XN9PbcRpp9BOAC79WhsNkBBXYhL
PABV65LzYa8+x5tqKdf3v0X46IAMWJ1e3wS5UA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U33OFhvyDr6TZQknmG9CiJblHCnuyjNFktguLuIFzd/VYuPGNPUXzm3pNVHAmifAJrPB2CT7TAF6
SpBdgM2KIeON3LRhsrRAbVtPF8PLeYtYTgU5BOY8SIKKoSu1FY2Gr1zMrTO/nd+RiZegYkT/1u27
xI0aTCkoWlFt3amFg2MasqdnOSk77Lt/DgM2JPd9muhj3QoSr10ZjlsDKpO31B9RZyxGfIMIft8A
zXeFtxJQH+1UZmzli9TNedfnlc4Etx1ofsn10PXyAOJjpszIhUCVPKZIY14gmxL8f+2bLkbtbsCM
BVqE9L8J6oKTduRVz5WGnDuPWMDwM24T9TA/dA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j6YL/khcx2/CEaOFv1YeHhnfPBfzoLLf3YocgJW2UWv3fiNKR3/XVXrjS7WsQlB+PoA6wradLkll
gsCEiQrgYuwxUEkrZPREX1CG/XJwUl9PKDBg75CevIh9+3qKHJGSxr9GydBxI8A2Bl+6FCqWp+ji
fmjdmpZhDdGqO9F7NIOUIknT0jWHS4jX/6J6w3BhZ/5VtUKxAeh4CNotWM+2fGo67UsEmFovMSdb
AWdoeaA+uo+Nh0kX6bc0yzej6R0ECeV3uzW4Gr9HgZtmqiZ4XMox/30Qmatsy8mCmeKd4pCcCVaP
xJ2QjwO5By08VArjkqF+F5MjSBTB2AgEgKQm4g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
R4scO4k799ATEXO7Aw3hlXnkNZ0vVZJ7vYdnkigrFS/XylZpGTM7PxLt9/klyjgZEX1L5ZFv9rZ1
KMFH4o+lz7ErNdGOBRy1B+35QtOzi+EvGNfe6LXPYHP9ZOdxSbh8AxoarW066ytP8o+8KcQwoymB
tFnzktbTUApejpw5IZJT8BaTn7itocT9BpYlsUDml3sOVaMAKKfOQKrnJWtU8hB1SvIUxWq+QMgD
GTfTxlPEJQkN/Ghdxr5MgvvkvpHsXE8rkGQz5Wk3qES0yd0Nik5ISSjStg9gGV0LIK2dHMBJ6hsI
UVRi5DqR7MoRJ+7jbcYmVu3mvDNRuC3PbVTHsVlO24t7n2t4QSuk/3aOz3M6+QAZ3OUMFooGmpKq
JNeKznu+ctXB55jnRq/n1ZgQvGFtH7QuHErOqIUAIKZButkHYYbbCzYQgo3zi8c5K38Uqm35UAxV
ISuorraw4cC1wWcAtea8y56YoHuSwvDjKIcCfClAu5N5sbpplWfxgvAF39Q4gEtNPZkpjuPUiosE
l+Fx1udPS8CVZjC7f6blgttI5HwCkTC6g6uoZSXkFiAuC737l0KSzASChISMB8uERLask4bXyw67
I9iHPS/Gy7IScBoFoelVbfyw836aSs+L1p60wE3WC1p8vPKI7nRScstLcBjKiRKXnm+n5crxT/Ky
Krm6whk5at0gwaiV+zCbazb8EgYsbVikMk9xf9sZOs5zqN+PIkaCzCVxQfIRJdosvNuWAfFJVMJP
QMHKdUxNuvBK6Ywlti1kKyrL4BEfTZVWD6dCy8H+ssW0PFIxy/eYRzHUUUlsaOTO39gekVsN3PXw
88L0lOINPgghiKsEPIBl5sw3sq/DfkNpxhEVhKe6GvNl1tgW0PdT11lXOJAcAcx+wD3wbVFJew/r
nIi+2nYEROyZ02oUpPTNeNN0sRsYW/ctnStEC2Jxfd+ZjNP1NdrAw7eeayK2sp0EYCjMwYMcMQR7
FeJ18E1isdb5k1bZG8Wyz8oGUv3+r3gLiAuIluKRNgpQnONoNdQ//VI5QSOpw1hiUeD+A251b3V0
f9Rrkvn+9q87LtpZKKothrM7o18qKeSHiS0vI1Bpu8CTTSqDUPYk9umKCbDUHOKPz5O+1fclG0g1
M9Azhx+k/hlS/0oqyNXal1lKhdGzT6GIRU6ppffbc6b8gudB7pqCQ/Zr7WBv2GmQ3SLEJNHk+Hie
NAfhG1vjCXjRnamWO1jMr8hRXBo40vNaBFqZPSOrGQRifRyM64Re0ZQ5Bqu/dRvruIbReEJ7nOff
/4XrZsz3l/IDrEUln95ZUVZi8ysqXRdmwoR9FZcVVB1oGwii8Gl8ZyzZuiusxujGim6Pk+oY2meL
O8/RBeJDUpD+oIH4qRe7zfjFk/+TOAm2MZh7/Up60Y0/5URs2Nnd/UrqtB1bxag0jicxCLxTAK4T
xRjBQRQSM95eqe1AnpA2Qu4oEXaOseYz4WoDtSUU5fqSQuepSFewOLySOssPOrDydadxeOvNRYAv
u8PrxLqTPjHqEbgcqDolI0q2XutUQgtE/p+eL4mfauWGwaR2WGUQ0t/SZ3Ystol16ILmMJaY9G98
UcvqsflpkdG9PAhFUjwGyoZz+a5j+VWBb9JVgkvxUFdWuyIGyeAan8Ty6nA62GZz97IB4R9s3qH0
l5FetABc0iXdnW3TfciSONYQJxGG/x6BrSUaLnlumzCTzHdoVeWYyainpH7ziFExS/EvIItqxGjC
hOaPvN7LVB4IXCf+ZtwOa4OBiyFbryx9vIgzd/o7rBbtzSyBkcxJYzwgTykI5qc21C3El8M+uloX
iVn7DuFEZHlywCSYBv7s72SBFlcn35ATQlfxg3ii9Pixw3YLTkYsgnhucKODbEszTsmta99BUate
blCKL/F+C8vUVecarVbT7Xw6zTGixh1X2XG0fqAjG50iL3j38d1LE7YfXyMTLhbIuCyR3ohb1IBl
dvgH9KRlgDK8jsdfNfYIknEnrYq1RiZO4t9l8eHoCFw8UknOklQDvZoA0N3CmUMQzeL8gMFocIaW
dlRQE9r/XJEQeeZaOaOLhYls7mfsVBWzJN4rtBWiZ9xp9UuARb6cwTp/TmUZ6i0AZmz1qGR6P5ei
LE1PuJA5DYjl3/w+nqxbWXVS7zk14K8FRxsqc+i7njz2ZD6qa0+pdtbHKekMETWFoA6owDZG/SIN
97iAt6ThNzdkvV0Ltthdw8gxckMsFXmT1BBu8toVcA7EIxR4WpitfwRxOCy49nJeWmKDRKKiux+d
MEbDSYywL4ezg2IrPNPrFPxzvBTKJlvZu8COqwYTBPHryzKwv6BMy0VOi7BiJxeO7hwDl2xLvZ7B
jQ1NYEKi30wSaPyPnAywkpmy/6sZvKx8PMb4LV3ZukGVxiYmHeRYtzbYl9u8lMfznqnH1nyLroKH
U4dvQFh8P5J6RW8J7v8XaeGDRQscYBswlUocsTPKA1J8/ZyfSfJAELz88kChQi+PjrEOSiFRXdI/
UI6/BjrnOEapsvpngBh5glUgL+x5RD5KUzncE/zWVW3JM2hDG6nL/38v1CUFeqRR0z3fkYFeJF38
Nib6AxQbe/3vXsSYDELZjUwGlLtTUHl6tHgoiu/Kbfnaf4Nc7kOvGBq5jHTnUQ5UnfZ9QNIs3ovt
GIaI9lYMIVK9GW2+5NXwLJoP7s62dZTF+/bXPuN2N9C+YgWzQF/+QsZ0nCvD8NV2nFsPS2E7n4o2
DGgiCZPjgtPSpxrpydDdBxDdd2xNVFBYPLFLMUv0JXTusO9WrA40MlZ/8BG5v3XOZN8S38ArpjJA
TgYfstgFk+GLuqqfeaIJJ3vMli7nUwj/5msxwaYt9waXU5aT9Ci1JDJDTR7YmY4neTP8OdvPHBL8
XSc1NIgv2QwmF0wCeJBy/44ArJ4c4GWIa1j6TL3rV+V+l9nvR3av+xoiI3zekp6IUGZycTsMyCcs
eEg/YVPHawhi+ycucLPQwqkhG+4wrsiDPXhaGWbXX2v//QRSPsiZkp75F24TN+cDE7Js1vfdjQAv
fyxLRDDpZ6aAo8XXwOMTpT3SnNh73IKbRxwIty3xAraz4MGhQmfhT10hHrSxkqn7fP0kDyMISeCH
FlihzMQW76yvAUDZiY+2zXyhIoNoxsujInTkjuffd9RszZar88iCpqg4z3MIF/4v2raauIUQ7XoI
OZqrGQ9pOU/udBya2uwcIxySW/5gkQ/HTWCWhbwlxzxA7xIHiWNmCRRQVsCjWdhZrzle2mz0FuJN
U2drmeVgXvMA6LjeUhwlYmk4qYETfiC4II4YOHqGOmHeu1MiVDPEqBEZtO5FwfjVqrWrlm1zhUqa
NgwkrPkenlUxqtu1oqOAwAvW7slfI2OwF+iWBY1I0HraULeEPTqtPzBif3vNH6cPd7JPydaT0Nm9
hn2RbeALBESMH/vzeT5afD6xcImQUXhFQziNIBLPMc3dVFzTDkzM0o4DHPkthO0LXhTIcUgFtFM7
AYoAYhhIuEV4//8y+MFWKQZveZNjakItCzu76vyqG1F7gaXVZXMwvxxTVwKxsWyGJiLlM30eXLgt
XMvrMncSV8EMyMprhpCa0fY2bgYvuzXWwwXdIWSPBXBpPh+27pfEsPjH7tLHq7nd9FD7MtUt1B0n
qXfApP7VYKkjAiR/cX9a6ErESONAhW9413tOe+1xjAzAJJcqNRXnZwbeY39DgsqGmJFBpq50pLSX
H58hCtnd+MumZFjh32IrkJKzWaca3k3qN0Q7F3bE3PFnS6NSP4gO2aHPfrBWAzAcRxn0FKVXRYz3
9Lz2ub1TiN+yZPuQUaQYOFl+kPChwm7f5w5J5xN/3nSl9ajuYg/ovxw2em5ihxT+nLK06TcBjcAO
Geti2Cv5tqeuaVp/9+2SY3hmo4tNf9EeBrqBtHycgchuHoRb/zdbATKe7W4WX4a3YBy/16aaQhyg
NpuIZQAXItyCXfiH4gIFYEeCQNqN8Y+vIEAYEfVEyAZlXTN54Ajhkcjec36LXqG3NnaNPpkUQizF
EWY4QKlfZftesgdqURMxPCahZWU+YcEeckU/BbB4LKlP8xpacDWrUYbLFh607kpJ7m49Y4XmCeXg
hAGgH+CtEb3kOeNZPfMSVLHHCCqVRz/KiEn0+d3EwIrdM2+hDVhLLT5aglOris9FoMFB+W12hri1
ro0hu0B4T9Lqd2xeUyi66t+ouBmWSlEGtwlxe8X9KNSQBU01da5ShsLTC0kDCiCfdVrWDPtqEoN4
RUNx/hoQiP74QsSxiw1pyDWaAWyztah10PR1LZCpXRLw9JBqwU40BQImm2a7hnqxVcx3S7En5uJ6
QZgsucI6vpVBKcGhdHVcXypesxF6uhkz5l30hifuNjojmKCp4CeBaM3TzY05ZDDtNHnHLff/+yfb
/q+4KqcOqabeNquwZ3v52sypfhsA+mBtjdQ9McNnXB9bmaK81zTBC3bjlLIgoS1BJScXeHqtK/QX
+9TgWrn7DlqXFeCcwiGQ8P1wMjnPtCiSsjdR64wwj6WQn/nQzjZK0a7VuISosRawL6KOnOsPkf5e
N5vRl0gYbPGX4DkO5GSz7vf2w2wDmQIsDWdF2OIDZt+zA7P0YQAXixaB1Alrpyzp+IkMgT2pwXo6
url0l6Z746oo/UqMDKVDbehKCLtWlaZMolhU7O5/HxNS4cJ9NE4q7aXwjTGRv1jizYvaTuRVR8fL
2YhwG6zYwcNLlirb5L8cgthZpZ4/L44FEOnx7NkF8EYgyi14NHudua+RRRoT3HRr4DMklegbyjcN
3LT4xE0tyGepFIU0VU0YY41O++r1BwNRirqmatGTe8KOrPB5doGhVT37AjX+HA7toWXsPGEq+Kn2
ayM/OxgpQ+H/5ksgeGMDxPtDKmvISorgBTYGi5HDv8bIBYnnQwcEh8ebjHRUSTRTzr05nLYy3iXF
cbb8ivrW2uV0NUaMnpp++7x8HYHxolPVWTKyqZpR0S7HyeChnb9BdTSp9NGGbKPFBXaFfV0d0ZHx
jNDgKKBUnpslR6+jIypvzb7JBaQhYNjU2hhWr4JVVmAOtPQh6vmMMwEwxnv0N0DblmLXfEeEa0Y1
i2xQk395MBtgDyAHONgy6LHJJrIgObqACxG8DhLYg34JEM23dfHy+CEgXsuu8ttV/kYx+L5ieK9k
4kldgIKI431Agd2Ky1aFVeHIkc4maxh8ILrDu9C/KBV4tkM/AQ+rWT/IRsze7I/3wrNejEdKWRKN
h236PjgjlPlSHvp6V9KzNq7VafebD6zXsWr2xg5ZzlhpJSbdqCOKnhZ2Z3KHallgRB16+F6zR+VK
zjzkS1mPmSx1wWdhgUsAwD2UtcNXfk52FqsmNi3Dlz1HQ3/n1SXb9CKPnuahZX7qQhyggB7UBqcq
g2e9AbvVeZ63LoHqAEybadL/dDT3eEZblB0KOaQFFrCPSzWyTW+LVRh1sR8iT1PTQupSzzpcfQCU
0lIDTG3CYsIKG0eaTiLinrKNUr61hg7ZZcRmxrpvXy82PGuDyQvdtCLhSU1Ez6LKV1PcNQ4gVt1H
qP+4FB/rlfpY14NJjwvAYRjPEzXtQQinuA1E74ab2+2Ykyesq420YhuARYBzkDmWoz++SSgXKrFi
OyfeHeL7v7mmtm7ZVJZ8SJy7UxMxvdMBC7BYApKU355MBs6RomFgMhhvH1HmQMPiQI8gNegCbseD
rKPo+S01NwgO10kcbiX4gvt4licc2zMB1ysfl3jAfSXAxgColpSpz/TQEdfMTP+UrrQsehM5iylf
fIEQwUlDo6nWmtgGEt8kGz29Yl5VOaJSDqMalhRwWzNrJSqIUYrtbi4e0YWuDDbyU4GsNVt8Subq
W9ww34feSXHi06xVQuogpIiH2qccrXGpZIE3RjbcCKk7UPsKtWHHqFipkVx31lPpEKDfw6r9QB0O
LY4u4F2RgdUO0SuUkvBNpEyueayF4Ry8Ld4BB+7isupOF11WPsvRQ/Vq2ofQfryBOigUxQL/laaA
oTmrHdhDImA/30UYOX4uReRvwVT89vshvLQL4/I+PLuDmwx+CNc48OjDA+g/J3WqrrvNEXBOb+xd
t+3sIBRztIABruproWs+zfkqKXt2HV/Rz0yYurTVuOATbuGBK74L0bkB1Hp7YKBa5avIW8h/2lP3
wwYEgu+gD6RXX51dpSXLVIkqTagV/dYSjzileJRIiQKHTEvsH9czcVQWOQgIwDRYtz7gJBGx+DIZ
CKmNBGtf3tR45MCQiZxHOa0lOCtDejc5Gi4rLuPENiesx8K758VXaWAlVFPQOw0Y15/f/ZBCdlDN
niKDv3eeF/H+rTcehhMIA3DftgMONb1XOv7iVD+X3e5WxipdvLfMHPtIhBYZzdpiYV6YhHlCbapZ
ZjhaUBctiPemtNGNFQt6E28RWQONWDq2rA4+uUOfl5gidiZ4elLDVPVvxpPVBLmxqmgedpsq9PwH
+KmVHlqG4OqjVqyzLgODYjmXr6xAbcXoMaquW4m56bOB4lw3L6YWZ1oI+4boy/gOaN/h/RLmu2E2
+JLTYhZxAR4Mi5GWhIO718FoXx3juEDo5F3UdrnVUXHCnhqwxl6J5PJTbiiMU7o5gOTPR6qVxjdw
3EBTzQ6dIb5QA0Z9qv6gEihDzj1DjpiMFOuKiElKPdPMMX+id1/PJ4O4ABwnDn66t8jewLrgNzAB
wuRopbrqipxLsFHUKu3IGeeZyy3kykCK4VFksb9nDsLxKjUZemG1QRVb0Ukct+yVIaUS5s3MH/5A
XwZ/fyJn6JKWDJaxp7fuJNwwLzllE2zvxjhZ+tWjOfXwe5f3ZEnxzZLisr7HxZ/+psDlF/dGPB4b
c+14nrGyoe8K6XKsT2+1eKsSkteMdWHx81IOyCZn70NL96KRElQSW2/AGw2yLwf7El08DXExRMEm
DAdfX4HnFGXwwEFMMFjS5xXtdWmrbVz4ovggD++6aid1ejL9/v8TrZaqj3KKftIN31YoBv7t8vZl
DAArQOqeS2P7ZhmAsOIPfR0jDP3qlsFxd+uPT7yqkuBv7ChVnHBru150OXsEEQqW9st0cFPb6Cm8
yl/ek/lCGPHgrzDT/y19L2qheU+lT714/UiHCZoxGiTmyicnu3qhuIIXK3S0tPI86bS34hmNQ/i3
e/OfYvPCCABR8wlsam18s2z54hC4/NoV0FB08MXcJ0poTpJPQ0Fz5WyOYhPdBdtN0KK0iu1k9RWM
Rnf0Qw4dEpRKymk589ti1LosETo43kSBACsdEtcCw3PhJN4hBa58Yk4YQEqFow4Z7xiinWqOt7LG
wYc69O+H+hN5/ftJSwxjasJvhJRZU07egun6CJtw1r59DzS1qL3+owW9VEG5R48mlkManNHpxr9G
X9mJ38cuTUHoZvZIf2BPUYiCsZhCLRMKUq5ok4HgrZS4FNLKnZoOhmVNx84gVDIUQMbTHvO80H9a
cuUfclUUQLvDMp3uWKQSntPYQFsJQgBy6/qgb9yaMeWI0uky9FquIgjF8KD9DQ3j9NMUx2+VrOqo
YfbwNwfLJUXNPqjY2pTNpNVeQb25RCVDi8VR0wSBCFonk4adFGWRD+nskgKMTCxAPcfHvJgfDiRF
Q8tx29mML5h7nO4l0WTTh1YEq7048geJL79iEridnqLMUJmViU273LScaixTRQWTZfUUdYPgzegt
lz8za00zRm3EwhaLQDbXmnmsDYLeXuGJeAmGLO4wx/nhcChYkf1gNy2gDCzqJtzPNAK6DDNCKoSg
fUSIIkldlFZhtYmwh0hfaMCaeKnGyv4Frkpq1/Y+3sSM4xZVfvJbNc/G0LlKqj7OIoyQiV48YkK/
pjg19bYTqXnusjmUkOfXxdmi6eTdgXvlgVw3LCA19x3pHBOCzPUdMJIzj6pMRC8Ai8r/XpF/TPPt
hNazLY5HZsRSawG/Oz/oYwo212Ayml2djlmS4RUr3fFCw6+1x5K53/Fl5cvQwwF8Yaz/gccXhVqN
jPriFp28eulXLhAdlq5QhdY7H8J1LAOQUoYRPU8IrRcZxWkUupHQ9knglNS6/hev10FGOAkp/mN3
IaXEqRHOnF8V+Tfq8g/V4GiT3uUCrwsqPx+EKEq5oD6EW8n8dVbrmDdiF+VLe104f93TEEuJfVJe
s4VCv4LLC5EyR4+df0rtmhEXJ5M8vz1OpRe9tgIKlLhO3IeIrZNYMzPXqDZdZmTwhsyuu88jsxl7
kKBXGoc6gLnZtTxho4kpY/GqlXsQVJ7dVjSMLUbPynJ6jOWFymKfEaydIR4Gy84ryGlDYrmslDiU
ApuZwtPcK9EAMfP4T5tHQjm9ue+pFlVfAwzWftyOdLon9veRTMhp5h0TxjYCnXbhpEQ0f03Uv02H
aEcO2ohB1qi36+gThwsyLgLjZuqzB8zS2tCCyhlawayXrqTf2nwlMcZIxnUNI66fBXs8KJovudHt
Ar2RzKHNfyMCQgpZYQrLg7ts3aOB1QRsyWW+lkKyI0y1+sRNOwq7v1v/CBatnAguYwYSqU22BOhH
DV/gY3tOX9G2s4fWY9vl6cGjv3+xsDrxnqU4ZP2bCaMqzhz4vw2V2PoDFLuv4rGdO8RU5CDNPmg5
Ve+3rEh/if3k77AZzprZ3o9l5DRXLjM0/Ua2Cm1MCrEedwP60jrqdQRp3CZnii3dZdBfCJYrS+sf
rjJLiHQuok+G5WioRSwlS88izZgymjPaE5q5iI6iH+tp8Y7tYuuLUppYucN/igCEOd09Ke62n3/1
X+FVoJ1+oW7ciVr7OpGySEnuzKtFUfZKEmxXUIMKklnj20yMoEhpzuSDrgpZjPrrv9l51rBi1H2X
KU7KvpLHnFyebK8NqVKoMvwBnhCOFuITppMPdWB9REPFUJojQ2tQvYaG0y+yn0m7JPb2A5KMQZPi
+/AZnbVPvbvfzokAZsxCiejscYcVxhfskthSZSwR2P//Srb21DefYQfzqjgQc3UE3NIukto2OrRK
6n9UCpDfXAXNo4tuK14u/XWv3bbZPmN7wF99FjTMuzjD7s0pCl9tDdDhcEbM5f++ypddC3G+ho3r
+sGXydCbyLwRS0ZuTSHVbOxyGSAV7V8DRXBuhlwEywRIJM2LqlvJTbktd9+7TfM9fdCkJ22kn0MV
mlnHOpRjsLbGK0wXqGueqFN78KcVvPVQFSWk/plxKpAL50bCWzpugJpEV2QnorDZ7uPbV+tK30tz
yXD8hk64pLlVZA/sSB/LOsvwEpETy1cxwXg4Bk7U7Xj+hkqzyZzLq4U5uULoWwkUqenJk1py1/h6
44KtXo9fPBxMXYPik3VWGrQ1sgWQAP2eTXcpl1+gSPi2WusKdPoP9RSaoY6+uKJi7YSFeFWcZLjC
Y8PDqdo+VKno+qfyiWLFo+wK0RlYG79B6qhyPsrOxAMsrWQq4xaZWwBwvQS10HsgB6nXIG6saf7w
ZuC+EZi5PA37vnU6shsynAfs6cukEyw9wrJOlUz701+Ji7FuBWrztnn3cbkKD8gIUxUg/Ub4UrL6
/OlN0dWPT0Q715Cxt/IdPUwMFTLdEgOovKbOvQBdPNqNKcdVmtY2LoWIiJdJn73EiRYZdpZUt9sA
Yf8CxGz1OKG4W5MrTaEFHpCGBDJOji4KsjWHl3FIJnV+wpItVFNp+WGUMQcHaP6VpTuKAtD6ppro
nzVTNdhuLQONVJ1of6P9pkgmd8o2pN+Url9rHGZMvsW9ZwN390wCqLHfl7mI28Tvn9Bl0wTrwg5X
+48WbQSNi6OC1z9iConIyNiUkcEOUsUneiaAH0saYJYSJcCE4i3ooUnTd+Od1L6CT8ZSTAeRWmtf
lD8c4UQvq3NFNrXyTeiPz/WmUmnSstKJ6Yp3YNHmqzPt5IIZMiKbaneNq2mowtvuAz7bCyZYObPG
qiTYbZydf771IRCEz6xFMla1RQYrt5AiRWXzk91c4N4W29NoVV5PbCxFmFqU2IO99htTqr4JpmWk
teib0VEPFm0GHO6Jj5gW/OsGxpe96VR8clCV48/YAA/Rrfcc2Kq84xtxci1RTnVTDAWY9r9n4K6n
JWRxyI1gKcIrE+SiqOfXO5JcQYjJ2ynNcQwgtJXPR4p86+iXYypo9fvuYEPn6JVNVsiKXfxaa/Iu
8XGbfmxFHx4Ubo2Vt78Pyx99i5WD0ocaOG/+exb4QBD0RMux0bA2ZxidoGdcvdw2zllPg3pJtMyB
Qk0Ka7CJ0uFfemIXoa02jH+Wk/ZJdm6WaJsioxiRDJCM/ggOEyT7ntm7r6amSqcT5sfvVET/2x81
CM0R3iTqWjcrZIIMFinThHpX299hlywxDE8VpkGvVbg3mBCTo3BhvUg3aqj0bFYTLSwkbUcbMIUx
qcMBNTvzZvaZ6JM4vpozW3LnK3S+H3vXK348cHVKPAnCMEPuwgiLbG3cdJC/XdPiS/OMsDUC/e9U
EA7/4V3EyAuI1YKYv756hIiOnaPhPMcYziZbZxI5i860LEjDGfjtWne/WYJZ/MrPcMfqZjgMSo4P
nR29WnOaLAtV/WpRzJ/TNrpNc0n81hVckSxsxXfzvLtmC36IcGARFje1Hwd1L2vrytLVwSVEKtr1
q7GAnx5IVA78s5lFeCcl02KvSom6oaTMrWt1VFKttfiIONjir9M5pWkfZw4aclszZNODmCc4qnUe
MWUckfE1R8nBX+Hlp5IIHbCbRS4sGXhruRAHSc/Bm89+w6bomg0Gjp+OqnG7Lsb1dZRtaoKZyD1o
t5IJGUx6QdSzwqf4OtHlMj9xNc9x0VIz//70yn+6b4m7po8Fp6iUZua3g76BvVVBv/MT6+RpewA+
dnUfRsuYrZzrGlQii5gZ55NnZPXg0z92UclLUZdOUU+/AC6JdhGCwVfJeAY1zYJknnuZQAtm+mDp
fa/a1/ViKoeHesG/G0vt129cJDOAZybGGLvmjJDbaxKvXncYCrtKj4sBuywx9ZRDbx9Z/3JbbCLt
hfKdDWuojEaUZDK19hKqflxFDl2XIdEC6paq4zsBx6g1LvVsLo3xCld1t2g+9pCu8ANpzBKGmHGQ
ty3pVfC+E2pd0NHh2iMVTfcIBiz6tmLU94Ee00e63oWXQGrKogZ12b+/2EbQKBb2th4Tqsgj2lrA
DOeuTXDM0Yb2ZD+0cPfHlNG8av3bh3SOkiPjcIFs0sHuUqh5vothTFUb9CzQHT/ZdwkiwxhgVlus
ThJeUOxT6p92tv5YuZhMuURPbjttTKPK49zAEQXtHXag9CQLlohHindTqStsJBXv84GBeWYbFPVm
au2jepOhGTl5CY2cOhE5ZVUo+nepaV8K6kCrTfQ+383fu3XfdOa99aTw8ckXIWjt4LA0DpQ5Bxvg
lIdwjJba5uDuFGh3ANt9cpg1A4/l5m55O65AbZRN+Y4iwzum+cfpeehE6IPwGqkQXLG9X9Vy0Br1
bk9UD3k9UF1+J2FcO79qXMoIzIgwebmnqBczj7TQi9V3ZD6FUAWBodfGTuj4h0f4uZKW9+5Tcswp
wHnciGOSXqAZLLDpPXqh7uHA4EhCwP2z+WFxIYegRLLguQBykgLya3u9lwAKUp4ARnp1bM559F9E
Q1YVJoQOFSFIAMVihAc3EJ2zqwKcEY5pT2gg9hiE/YNmqPji4n2eWf/H+LExw89lFfcT91Exe4fJ
BNRO1XGudP7W2axupf2nrv7AdUxRs5EGq8j2a283oEii9/fhXAX6S4M6UjIhGSKy4cVCq20LjK+W
akfOK5bKbQcACASxZO+loP2AyE81mB8ycY85O8VP1qlbYC0OO1ovlh0OFKHKhjD3P7wgcxS+5WnA
0JcZL/ezrCz22IhHCzoPbpzy1qdlQcWhBX+ImE5E3aqx+EaBOs1urI3r8sE2tqFCGAm2rHpKDPc/
rlUJ/O+qatI7R5D02w646jJJSTDmk8jbik5qH57zl/6l83SZiGrFXDLNwWirLuETSLPq1XzPzXZX
VDXXnVZlJ2Prpw7zPftpe0vtcthYvhOx/nZu+GcZ/5TPBNVwlaq/QLZyQMXH9vx9+r87lXWQr7p6
dANWwMCt8J8Dg3ha6L9VYGXR9NW4ALKOKojeO7Nc06nvlD/ZbVS7/vY5qqaR/MmK9L8cAvkU0X3L
mNDsZVb8Y8Mfr8i54cyd9ELeodaG7rRv106AEvQIqDBdp5yMqlRsDceEKux+KCXjfMXIIh9WRKxy
bEjolgtnzRHvxIc+LCtdjxXzywGvrUba+sipq2vx3FdNB2KpP1uMFTT1ITDPZS88pHJjq0iLN49R
LmGGAKrKeI4JGRuZl4aA7rmrhNjgQ2v4Aps7ZoAHSbNEBdLVcWEVq5+Q+zPhKXULmf96Q/htX1BL
hxlR/UyOMUit/OrD17AaoOzF1BADzDRS+3DFJGXkdmFHyoVveMNck87esAKCKWbjELaL+8RbYUCK
dy5W29rTfgI4/AzPXjrE59ypPBbOH4XxUgm7QjkkxLTJi5+JtyO7zFlnn9jS4odqJlo0ZN5JMKqj
A4L2vZ+ZSJyVP4Jwan9VP3Z8br6zC9EqD0dhoKt0RsPdFwMmYsw8Gez/hUbqzjSXDHkxCccBUQau
zh8E3xyfA0JB+0gNaU9wzgJay/IGMXry6cGc1boBeTj+vgWadSGk5w36W5WaIcGzc5mM+KbA9dpT
oUUhxfBdU7w+dwJ89xqgp+BsS4/hrHK4IA8lReiPIpNBUOHUCAUng8BOoaQzt3bRiE1FYwlB3Yx9
G8YOJTPBH2seZ83ecmZ0o4uF4A9AvwzPbM/TeUN9sDx8UFJdIGIjl0K7n1OvoGtWqtZ2P1kUJO3R
tNE/efMFsNY9/KkJw/oYYVf9g9x/pZ9hthguIqWeyJkJpN9o+2Wuw857UFLoeuK+68OiXk+Jsa0S
+EMtyv5OWUIYCA1y8CNFpS1/FTbktrl1ZcUkFIvAz/lLs/fBauZbGoCKfexz3Z0CiD4hyPCnrKVH
9aydbUpkusX6nc2xbG/TEa0w4EimXidGtPAWIntJpLQwoAjVA9paqtgaAOc7GA6fIeNn/Swp1eox
DZvXQQ/rVmofqE1HeKb1k/bvr5U0SxiN7KYQItigEe/ebF7VVATJmtvF3XzEr9DVuq3Lj8xd+nnP
xOtb8Golqzrv3AHCfxVLwYxN0XePul/izXZvXFt/VxOvPjSIdO55O09/uufPGeEPzxwZ/WsPfPW5
Dt9qDuVrmcFZKVDSeKCbxkxCZT8qcQHr7JtwhSwCPynMNAedNJOL2+1kb14nGmz1o2XRGaeyx/SS
uAU4ZhM5ohjHNA/fwaAyXh/FavUyQpf+aXkxGlehuj7DCB6Di02AaYYEOEUbVvpuPAbmCreXR0S6
eoExWVC/a+c2UO+QPeROe3GttiFd4+hN/unsbbtmoAuIF9k1ZgxlZj/Z1c58ldNSkFZulvs6+uD3
9tG4jt+43a/qVEsaUF4hQd2OM7Ekwx/TXlz4bi2zopaKd++ZvMcj1nJqypJT02zq4zSQEy4sw7nC
Ob4+Ko7kkUmFgs6aqP3T1UZhBE3lQu2sCqlDcAR9fdWtV10rrZAuDpChNyb3und7Sn8zqrfaBpJT
PuCTVqKmW7kYIhqWgvNS67B4lSELtXOFOQi/30lPW0z/CkX4jgSmqz5IcEDVUnGHOgQcg5cYSKD5
ySKDoAQocU2Xiyc8rWCEjxftbLLEjwdz13zC6uRqHz3AF5RgNVh/XV/UVEPtvdPJ/nqR42Dd6X9c
2ST6LW4D8iQncAEw0Zryya69t75GYte16KD2l86tgXfUHV7FglAh7pMg0EtkdcGXS8ALiwJJeAhS
y5nVV3jTNdrZSPM8einJlvN1iGDt7q1IGttzdYyJrrPyatP882XlBn7lqosAPEOPSVcn/b90+WtI
vCGBw+D1JinMfYbGOd4TUIcws7JeUrs0bgc9aCPbAgW1t9UyZ5KI8x/ztyo2t+3Vp5u7REJ+CTr8
wvi79aG3ivq67BY7Yd0CNlFwfCJd03pncbeheqtgweowULA5WTjwH/D/eRBik/7mtaBdfwCOStQM
VegzFFkPSls4UvXuIfVYc/AoRN+uKbFg4G2v07BEgZVhcpwzQZlCf8wkegNP5QPSD1LL4bIJPmTO
m2e7OazgTCP+EbaIgj9kZMuRVdjxa+8w7l5J0luE5sx9ffHWHOmmB5qTuRbgvNYog63P9un1M5jK
7qF9q4i7bjvrnav643G3xKOzHKSuvieG+S3HFHd6pzR1aE4K8g1y0fhgG3EWRJ0h0TutQG94uYI8
Zb7bCZ8S0G241JWuErjWXS0c94o6xt/rCEIIeanxYNcRSAqOlwok/jF/xCyfIArpMV8cAh/ORel8
O3beRZEezqcApVqQCiwneLd2IMUZeGX8LC3Pr6sSHrQdvMyLv8NL0/aU6YjkZg6CjqrRY7+MfMhw
5JJT7CNo+loBUPXWanGvpZvzHuMXfMfnKygU7EntbwvJNNkK5U1dnnGlzW7Pof2UFW9M8ko57k0v
5LE6kR+pWhmgu0CLUlL7crn7+mWI/P5HrP1FXocmCN3FWhAW3gusRTK8IspyIBGOCGUMI4FTxOjJ
Dye31zJ19G3EMcwgWMlwNIXfKs/PDimh2M85lJS1PNeuSHkayO4EJE6/4bPIf2cO8UkS78OYZjjj
EXqDXS99Pk+qT5tWltIuustYZ3vEDlbr2e0vTGyKKSI6A0HY3Eq0jSjxq5juXY4tOmBFFVmrPByE
gX2yjXtBeuBkY1gPQ8U2T1BurgC7HgdSucUQ62oB+atouhJajvDhGjQi3ZsMztYe+coItb1xe5w8
mHJwmyGRgHAyvdWpQ26LWfTaQjZzCA5UxEMmjd85OjCuUFLQwHp8oTmtaVSTLPKtYXYhIQaTHryi
BCTlXybrAR21q6RZGuFAWSZcS7Lr5db9fRUnTaSD459xN+mrcNHeBL0b0V0xpXIIOTY35ZDiRIzz
/iXXtWYkE3Qd5mdqvluUNLgbxO9O6rJq2G2UeOi62BTu7zqpoS5S8US+ieZE/OmhbaTX6vlW6w6G
ktYxsLAGRSBmr800aP1EJHE22LIJgJH0IZoD1X4YHUUX6WB9ZCP5UJz8Myo4l2Hqp1R2AUWJlgG5
Q0WzJC6iXhZH7/RYJETWqbKpi8mEvRLx6io2Iv6F2SRrgoHOQO8L/R384eyy0s8VwFOxWJUUlxat
a5pDU6xXkyTXivdRGD2UMB7+iN4060NCCvOt8KSGr+moMZwflGBKRE6G9DYau1H4dVVMkbNdG0o0
eDlx7fqrzk7kue+gMgUqiqq0olynsDdwpTTkY82zmZ56bF22E288w+EUQInc119xgICVfLKdHu0o
4Nq9Ll7R2wL/pgn1J9BgkrrMAntHlF1USOYYLndRMJy2EF+a5fqfB+ziZD9+k+Ql1DmYvJQJYSSv
v9UQ6BGIufsAWHOGHi2ol+TFez3IezrAe9/qfXQKKz8jg0Pit3f/jsv/2e7sx7SMw1ov9kzQ6rZe
wXV36uf8MTj5jKH017J/22BFCyyWE0jhYJHDHTX55OB3LxOn6lRNxGJzhJUj04KoCSm3ygKVTY94
baWpsHIbaoDXij0PDgsNaaNIUf9K4NXwQbeFo2FfgqwujLfyT/iGNEb00imvhzjC2P2yxHqFcGVY
gXss+Za93Xi4x5DHdAxCsVW5in87c97seo7mm/gdHrXaJKd2uUMWnuOIQQuqalODGGP79tc/W/+Y
3ETUZHydY27rpn+A5V+Vsg6Xe6BLhcvFNjB/yaYmF2WFlGqhthX1cBKrHoZ0C/FAZ29kVGSUam9W
cyNZwv9XOdbKt9hSW8TgOyx9NL68Oz78m9F1fDFgLVw5zpL7TiGT+nTz5mkA4Sf7LMtY+Od6wsay
EYhj3Bryt1GSjnJ39elgjC2HZvdor8Qe/7I989h5mQBaDypo8cXJOgr4VNqOEvCGcYU0BWzRE2sz
118OAQdquXHyp2a6T+x3uu1v92BjpF8yd1lu18GrDtW99esBP811CI0AvAH2yNZXCf0NeI7kd2Pm
OX+Ykuqco5njb9aKdiHN52I2vspjTCrF0yipk7z3BAlkWbqO/9TARjrGutSGvuYYgat7TeHR7a72
uyaQijjQv2l3i2kCarI/yBLSPtoZ0+ok4TbYdUH5/4mZH34KthOuVr2rQ0AwMs9RITAjEDP3FlME
xTFzRgR6QR7pXh0i4F1XrRN1CY8QOcvPdHcdMh4pm1Nueae32BVGprXfw87Nr24qdML3xBaXvt1C
WsE+8pWPWgA6fgGULWc3exXr6lA7AdtWSbtsWIUIfCPGAYOARoqRzJsOkl7tjVHhIt0V9y9JM3iJ
9HMOlJvjivZyi/SCKijVunJtCNRwYhGjc78hCzzQAGuYo0WJdK55O6ujlaqxa4pGEl1EjkS29Wij
bfzocwnHYak0tV2SBYE5vmmSipYPzldgh3wx9iyEoYqbbcl5JidlF8JkENuyghf6XDMOVq9/aeK9
volsYbUiaKQRQOuZ/NYkNSydk3LfcchwNxMtx02gg17559+4j/G9Kb3CrRliSdqrjn/gIXR+8dVC
0/Tjk+B6JVnpkvz0Rrt7o/c+8ZiknbPqqPfd7xW8Xil5kUBIS3QbBrMQjVkBUvNRzjE5q99OVADg
EklttnIgdk2YqECoBS/YfzPPv3IriWcUCShlFEo/Mnv8UefU1bfeaHcWM42rMWYcXJB8miSBCn1Z
MBMEWDgbj3zN/gN7qtYhPWvX9MXz8T117gkkJgA9GIBNqGaiVhZuEbJsNJaOIr8sfn8Fez3vipeA
hqb2C2fSX6Gde+jiMz//OADJJjbCQlXU70S/q/yf3MpEIgrVJCsFHaKDzItMbJNc0JUxx0eKBbOO
MKEzsWPIXCRFKmOgEEZmMS4TbZLwiTcL5PwVlo65v6SkYfpQc/LbFYIx7iLBriOH2d4PNek0Vo04
8vQrLRO/qMMmfkzWWCb0KVttCWjtTCUmsomuffw66zSTfi7DDRJo1pwX0i1wFecisEShylzbRQTc
o7VxzSaeVrbrZgdqItd/FvBCyI9k4Hskb3jXDoL0TRvx43f8ixya63lfNBCV/Y9jpp8zCfKa1Zuc
VIgK2om4yT9HzpOWKwIaKMo8KrSqY1gOA3tH0w6cE6yatkXz4Gcodho4V75Nl9VQ18gKfgXo2pES
2jOb0QNStAlj2Wkmg8LNCkIQj5bLIuFJw3rpNEtqRmXZTTL/FhHczxZCt1vZ55NT+QPSDFzg6nAT
+c62HoSCDo7iihLPKjZEBd73oLY90mwRnyfpyJJTe+Ig07snYlsZ7P+fEIjobIIGtx0eVXlxJ04y
2ftkjXda38/lNRA4F3UYfSOmJ+kTivJEHaXy84Yek/Nkya54YMvuk784x7ddBm1DhQRAU03TNfW2
pVLf1/h4sp9/lQ9Li2Njw0A8xrango3oJbLbDAK8QrJxVJ3UvMTId+q+17hWqC6MqK2pVqgaz60s
bJ6VpPIlX8m/pAIP6qoRT1KWCsumNn3ujH6+Q1e8ZIdbJEmxrhODySVLB10PHNClQeDq5rYtpdfz
kZSKiCU4Qi8CXJGD02Px+691cZgYP/EWEQc6L2U+Q3aRd+mITN5toKAnvZ/iAQHg5/JYeKaPXed9
eVaZPv2ot3Mh14AzBtWUuWzBzYw09iRYqA8XwKwPsiI3r/QbuaJlOlfaeC+hSax3TiNLbCI9qou1
IuY3kRgqiIHFuew5Xw4jnp8ds4rMpnkyTCoyTE9F6DCzAEEQUq+cG1STgr8ojj100R1vTH7DYwus
QE8f6wL90hVPXYqra22xCGPDUzeH1ssXKLu7c1iOzt6PJ38oEsBSmKTl2b8oTa7TrP9cJ3AZkDPY
eyKtAMAIIhYCxfebeU74r4FYyed9bZhqZCqctIeqoiO25RiVokFwl6h3e/nxKagb7MiE3D9JhaL8
tfzRmfVoZJGxNqU4Wgmgd0hDV6o7eE+6v+Y7ioxfzZY7xVPu7SAVNK4sBnEjjD7W/cLbrEvKkBr3
uo3U8PNqxSbVxf0h592IpUUkx30BrxE4q9li4YELIrwZbQmTig/Xh4lu/PuPturiqI+QRVlprKdO
/byhjykS84Eb28qXg+2XnYKEdpvVT8zTuYECY8z5HnKl0WLeA+nJ3nt61x12dm7xIXTXot8WsYeH
JDkkvszOZ8BYgxZ9cqmItyBNtL5Lw9EzqCyfpf+T3zCyl2y2tBDlqe7M5AuJyE46KDYtBidMxJVf
KIleBugJTacyR6CPNjRmkN0THTmT/m0qpOmf//bJwpb2w/XQXHt5LbkkIBozxB7kx8SyC3EY4x63
l8xgOyHCcrQK2zcY5T9SIdc+WSUxwEcY708qC7SjS8WGf3axXxQc1FDoWi0ndS7yyPqfL9QfoI3B
xMadhl3iLlnB3+ipHeSoSrH9u2tX9+eYyge+WXXOrFRLYnzQL3qgSq/KRbiZx+yEclu2WraLbPVO
qU7LDHIFtzxB8v4WLugTiZWSDOusdgXE5sGpc1ldrwMfvCbHauwzMinDMzVWrc+86w37Iy6T3kdG
JYqYQYlNxL4/Gv7blPtPfLEUqhf9s8jTnUD/rv6GyzqjIwlDCuEgqYZdNLtDEN6CUBJO4PLzoKEi
b7m5Hj07dm4cWyQKLDRo+ticVl9JR5ychna0pu8HJRoJqBtiQAZ2O3s80ql3EjYYr6OJAojA7V2i
MLMdC61gt+Vtt2AjUYpudclpIF8K3siAFTc6+1dR/N286pHaWq+zsHsPVJt2w/dG+IX5SlSQDkgW
VIm0rBe2BA+NdDr+ZHQn2GPU+a3nK4slphapw/h+/p6hldyFJ6iTb50sgh3fLtDCO+cZ3xzxTLY5
bgq33MVvjfTFTNuzn0Av6kV1FlGxBZfRY1RcVRGy2T6vBZh2k7V3h51bItBvDRiZl79Hb2iVKTf3
crFl5RWfD4TGvYt7pfKDUCy3EcdI8+HFq6FhT9n8u4wo6zfAWyxQO0tFVd5aGGGPWjjwyZ5R8ihO
mohY3kYlEnb/RH9QUvYh9CxudXAf83CYzBQqdAj/ExY7frNL2OIzg14yiWbubBvINqqtmO3I6hdq
euk8Jnb9pMnptkVjjeQjTjcS3ZQHn2t2M28nisYzCgB+/ksFB+HPP2DXHCcs6wyJ3FFK4n6h1NPV
H04HbK54ZPB7g+Srcq6wG3wvM1uIQRXsQnREO+XaGFepOid+4ASIq+e1plGHTxg8g0d45MQrIs/V
jBtMA+eOnAKYuiWt4uXe5zopdEGVxdYq7RZbxMjKTPW+fA+u7nIDUVyKCtAWRZV3KWjticdiVtvX
huOuKtm2W7R7+HLYlI99TYt6spZWeFKHS6QMGgT70zwWwvetNDh9CtRlpcVJ11HNuLN5sKpMyOhi
TufnDuOkZ07+rlTCzdkc2woXMNIS6Unv6U2N6p0r31Wc6BXmyNvXne+IstT0H9Bh8SP0Js+tKOt2
HnTz6Whg2hhnlNBiTXz0t/NlG/V9vYKHxscyUUBmjjceHH8ba9VmPmidqITAFNfvsHnXE+r58CPg
NdyUhHM8/B/jsI7AaKFWOW3ryMVyQL6jGBYBSdKQZ+9Ia0UTZ9R68aM2ziP5YIl/7ALHF00Hlr7U
cfCPCz2K4hjU4W1ET6I1Jnhw3Hi2Alc6BzUxQei1pkvgn8MSXw6aVXOzaijkymPucMWotUHM/OQl
dp5ger7iRonhjXL23G7q3Wh63ua58racT02IXpC+vBKhtO0yqymT6MY5DwZ39BfNJOyPfU2xZq35
Xor9qkxCGI8cnQ0k9H04A/hTm3g6Ka39QmvOVwJ9akzsmeSy4DRhSYSQkYQeKXoQ6ES0YPg3oPFg
eMCRGZ86lD4PnSXurxAE5oLAdauFDRlbU9z/7rgNR/5UgDQmbSd+uTJFuqJxuAElzverU8FpjoRz
XyQjFY1UUW9yW6rlcJuN+0Bf6m2GfVITzZRBACsGF+hegeUTu+u3eSQsBcSen9BZb9TP58HUrWtp
WSc6X5GmNU/O6NfguTk008BXMYVwT+fHKcmTemZuues8xElozANRuesG1u7M/9tQ6p7SG2BjBr6o
XczPvcNOr37T2rqCjtWwOJALXqxzv9DlyNIWtUnbV6XtWWc4tn/sRC57kG9nXnJhvGBGApg4IiXe
JRBSi86TZevW4xKTIUFG8pCkh0YJvmkRXU60E592t4cpU1XjmxPD/Dpyqk0CyVrr8pDsMciFJgqU
7rGugyJ5chBjIQEmkt+5Z5/tN35azcjNzhzCI9uYhbOACygg1J4srZ4vf9qv8Re9hRT+ktGXnhIN
27Ov089GreI5hIl2eKRP7VCLccpWgCmtbvZfYetuyEgKPr0LD6OOopk4/hn8z0voMBdYo959B7yF
2OaUCNApu9Tgjte9p9e0ES6GbXIUv8mKMZMKJHNDnvYUgvZ6q4MKQ2TdYncvbZ3BGuayyot1Rugg
1O73qQIL0ToCxSSr6R9inXlNQXsq2CyfADbsur7H4wAH68yaSiVX+l0TCrG3HofSB5lhvbKLjW98
R2ypOZGEoSSB0xDed4hxTMk8+5ubaZj4+kniu6AKiBP0NJ1tLeKDp+wbSpu5I3Ex9M8uZFLrB1sl
ci2wEh83Y3Y+WOJs+iis+rOvowpINGJzHXBnY+xZtxwcbWCNcgeA62oCYdD7MSh5DAi76V0+dhRT
TCYI8NCnrFZU0QZ/25/aAlcMznaYB0htHMgT3XncijQbWtma7oZxaX4tCGlSjpJn445HmQlPyQZ3
az2762v8FBfs1kpMhbvtr1wOYDPctzTafT8/LQyd1Lt9JJ+axvWNpElRj0wE53JqO//CJZyuJzZR
b7vXASQ9AI/u8QJJu/FBqn4D8otnaQ2MKNNdJVBOI1lYsUClRP041LXNmXUt+mZKbWHM0iC9lg1V
xKRQHXg8BAjiY47ZPNZ/oRs11jkzRJx7gGU0q2Sy7uKYTNfUmVTzHzXUlbBp91J9RqYlDLoFSSWU
wKD0aNebcK/c3XVdX5OO/PFsQbldkDeas6MLYvyWjeL7UC2ojhz91ZFs98+9gOJOfMnJ0qP+DpxZ
1PIgO1M/IdQn4QTAo4s/pztyCso3HHJkW8L2m/jiUiNWLkh7s/i7045J0j5NsNlRlnyrC2gTWNkU
/BoV0ToTFbwwngGWOwaPGagrhoIw0WxlSXTmTtLld0n+WBMQBh6T9t7czIh1uPYASpA/kMhafhPs
J4hNlpLzRXZbzPYMFtQkYgxSQzccD+kKHNDBvNjjGWvAHwgjm7XKyQ0PRslRx/wOYK/hw8uKwTqU
9mQ8JiCK2RQdKNvqdsQKXwByNPaNZSHfDlwiwKzvpMW0QfLHgy559vVzmzt71fnr5R/7ysCK8PCe
Ifx18k5ESFCPMN/zuidybjlIGMrFZv9rwJPDsXToyFSFd1227zijKYElyS4z601wHQjCbbNLpUqz
pdoWRDsedr5ylwB6/x+DyMEqxrZQrU5D+uHRb2NGpw4tiq1Qq+D8+6RZQ/EJ/GxxX3IlhTC3merO
0nRQvLzWArNGe/RbPdRcKXRdx6uSy11d6ygYbB+hiPU1rYL5qPMmSIsPGLPoYG3wHMV8Ad4XHfB1
iqDvXtLfFa5klizZqHVz6tXWRZyY0ND4t2KBUBKE19OBdT6MT7vLy9rR3ZhhJ78rexUjRT+6zh+a
trTqPYvNrFqmtafpxKn/NMx2CvJUcCxWW61o2oFKGRGJ6N3KiDY8WFzDc+ko+NHcE01g1/zZX4od
MUJ6qv26fE5qVcBizzqrGsHwIPColOfJnqvrfEpxHjtZLM091e3V4vUiTKMYyHEml89KUramun2T
7tZ9b4CUE8mwz4AWau7fv+oA57q5ZiVa6EIArwVyY6NjSiCvRYf04q+KhGu4UV7CUfOEaYIQbhpy
vytAOVCn6TwhBFzuSWNVKKx9xQfkDcPdxSXvjY7fXG0quvfpvIpgl/G6PYVy3oVjAmlEd0EHesOg
qYxZoG3zz50oKgP4Tn7fiuxxerxzyKMSarYumnYniZWfG+OaWvvvYk2AP0K03K8fEk+aD8Yifw9g
cwSdk8TQMOSOu2eMDWA78aSQdg3Am5VFzV/E5xcQtDGJPtfz2cLR0nCoih3VHBIEFalFWjwjzLgB
zRmc7RoKR6Sz25k7RWbZIB5uZT3yAG45zAto9IRwH6dbWAoOZ8hVVzuyiqrgzkakrbqx5GzjdFwF
5NLJ0slh5Oe/WEaN+Wp22z4pN42KjtKJmzHzHxJYSkzu/hcHvG770NPLbR7ORxIeMzZtNARKSiSn
GRng1MKRY/RDbSVE7qZn6MFA1FLTdUdBQgafjiQ0rf3+YK1YiwbFj4+UtmoFLedEQu0IvUOVQ2QI
Giq0LtkFP7DAMcQy0geBNmFqbeX8/z15+/UJ12nOwqai6RE9G0rVhe0SGyWHAXGp4u4dqa68ePDQ
PY1A/NNLtbKBL0mhEXpG/VgGCBHd23uTTZqT5HOJW0+X0tV1Q/f57TuUf80a6KTiD5g44n3pqL+a
V/S3JDMXwBRFcBUErctL/jY04lPIe9601YPxNuR7ZH9NW6GlOIHThJ21ZlVjun4iF0goFVsCptAp
lmGUfxNw4OxA5xecj56LP4pAm1vueBYozjQuHkfZJR3VzlqKDZ7aGq4YDbBzqdFLrPAZ9lONXA60
jV3djkYLaUi48rul1YU9YbkrCQxlV0KP+Es3WGitKufYdRCAtFoa5mcAeoKRvvYKabXxhzifRhkB
Fo28M60BKjM8SBFCX/aofBGZBvRXcS4RsI78s6WLoaCdRI+npdEpVS5l43TQJ75hqOlLeblMtXU2
By2AYRHKbqMsglT6uAdKNgxww2PlgSfGiWzKT+oHaSZ9H6+Gs7xSO9ILKdXTfa3d0GQFP89odsQJ
xsanjEz4uKyMT1dJV3NMiIt2pBbZ19m0kRJhXoK3o6xVCdfZfUxoFmAzbL/8h0T1it3xs+QS+tuD
uCHHxR7OnXo5G3ERm2IMf96deNGiQIgwadv81xMVmhoOnI59nl46s5sQy56v+kPkeWQpyKG3wLs7
N4wzKnLWljqws2r6uaOZHkj6t3yVOLgfGWb3xkxYpboiMEg2s+6oBkfNUPfg4Tompn77mp/S3f1l
+li9YK31Mh9BGUBI8lYSMqO16U0BBopmKk1twbiZVWisSSF5QNGno/+HaF6tGAKYrlEkh165xYnc
bbKCc/21QC3bvKq+TJMNqDTTCIYY48EMJ7rZ+rcIMpFuVFcKffnKk/+T+pxTyhVA4bZbskQGFSQ1
+sqIHW0U5ydDh+lqzbkiVp/mNOkgxl8MP1EmN89UVCpbuUcMgFfnfh6y3z2gwtwe5wGwT4E3W2H1
OU0LDfQP7iO9u+ClJ9TdkBQQdF8u0BJfFYa7SJkVThx7Zc2dxoebwZKA5MP+8Dv07kja/aCm8QqN
O3V29d+4tLygdrt6vOWvnw4sWZZBejiFs4Vv8PuO2L9TN4SYiJgjffgV6Wvt/kNKcluVMpXRDsfz
nERVLMKd8M8XmlUVz+xImwYgjxFb1TpL3+27lL3yfNJskzOEe6YJMVqZf0ESE/7S3P8WU1gM5Iai
rMOKbYVGSjQ1hp1LrjkiBYfbBZFwBOzhFGjiVgc/3dqkwtKHgnMptpYcxh8cIXpMAJ60M9NHUvyO
9fm008pa2s5NwXu9wWC70RYpP91kSfYx1ERaCMpnevU08MvnM9DoReAh43lIji1RVWH/HHV8bsk/
o8Cg9GXDCotVuinQBQXB/2GFhEZUny+uHsw67ZzbF2HmZP6uhfTDdVQvQQFDK3jSpWOtsJJcz1Gg
tmzQssyXOxAXZZnf8nxQxfFvj6i2kNsLmQHQ+gOzfpErPu7nwsqzOZIKiv6sD9IMdKth63wrX3Y0
ZAAxB2PGvf0rw2hBTBt7YodLGufR6fVvBQQv0KKkdid5hhRpDohH2q3R9MVOzv5DKml0WF6IoAFV
dpPt8eiTuCsQbtYYWQ3nWaKFqdGJmFUS4dnvDKK6ngjvVBNNS2nHHFYDX/zHqQaKXJrwgUUKhA/G
KOswE/OTAIvW+p+yLdr9fAasW5xvgbttLjx31DCYfKgb/Q5UKLWyKc8CDuEleYA/dh7kKrYXfB2c
vTRocKR/plNPloZJDEBPfZFuirEV53b3km4moFJEji54DT8S8II6SCANbc6fdRjL10IKAs57aHZN
TfbO3Wwxy06EBrc/hXJhcZOcEVqRrch4lxMXH5OZMejX6fQPqVASAyph0gpmdDF+rT3U/3zw8cHF
TFKcntqCbpsVelIezaMKFnogJ3EY0t5DJ6bG6DL76lOAz3FQBSSGMRt5vVQfAjQS6fvMRum2HBMl
8o0aMEqeqCe/ZAicsUt9EX1YGsfZMWIGbvkUoqmuVpt6fNIDdFqkOMzt306IYgZTYWF5SpyfrkwN
qn176Ow9zZiEmx+T2bB6JBunDNeGe39rGZy70JgKK2r+Q/+5g8rkFHQJNf6BMqxffYtVvHjAXYkc
Wq750bxnhAgKAdETQyE6Qhgu8vFUNiezdqS2jCb+/5BSd+wG6hVTfzVKP7z5IjsUrN58Mv5UJV9F
LK/vYAe307vNUmYC4zqjE9UvpGdxiYcjlILRKbyjrpN4ZIalIMeCUKYIEeULoLrye/zi2KU+7N/a
g7ftbY+XYbYNa2F+y+bu3Kl+KOBkURj+rleZNTh/LRlvd27vHShtU7biH8WUGjcyH55Q88hTomRf
OdmxPFmmyZhbtQXVKZ/0BvbJsxSeVndAF1Z/xbuDuyzBB0dDvfmbmkZkGX12k9hcuccORYCAuS79
eYITnjYOkex3wA8h8K1Vg04eGf0BphsTHFzxulVoWsPHs7ZMbR7ylfD8VWywk9W4E7ZwxVdinjmk
hDzLgB7r+idWFwuvZTKzaPTomDP6jn2yloiPnT5SyA3DdPdqRcSkwtm8LT+eZy6vb8L6oR4PqqRt
uC1QQ908iYhQJHYwuRLOcSmdkkZyS/G+aB/+T11PhUL4fb4Fr6Dy+N6Vax4Xg/Pvr4aJP+x2seCi
rczXW476xwuq6R37qvlPN3wN/Fws3DfP/BMmO46zeLWCrZtTXgc/StokSr95ACqL+NfzD5+wIn1g
P+pDcvtNdtw6W6cjIeOE5kD92xo4ZtDB7k4ZtACVdanSLyO0bmVq0JA0TWJ6E/56SZXSNfBHxOBB
2PmPHWETJjs7mLO8jmj0rFqcGsOppnklBGz7dLwXn0k4+skNSXnhyOYPVTVB0FP6b5wbbme1b82v
S6WGlIz6z2jLj8n5p0sBjp6RQEgRfPcymuozQ5J1LvVHE+wvdq3GRS31vBpOPjCRD4KPrqSBSjg3
wRWtTWB4PbBt1eupNHm6UYAcT9s4NkWcMKQIAHt/H4NzxGcUaJuO2/HrvPGDepd6b5OK2bB6gGdq
55Imsr2VLfcv8JauPm5nA/CiQpKvfkVf/5Js4JZX+1jRfMRhn3GGGPTw84m9tdSMhsJtznoFpWFj
khfFqRVxVwvhx1HDW5kER1tNkTmgyGGasBea9kMPf/WERY/hhQFLPBfJ5U1VwYS9W9TyhmsqvpXK
mMvEXI08S8Q52cQjhr5d2HZCL/P8nmGjasnI9B+FgobnEiWySNAOPOWnTulA+0LxNPF3y9YCFdUv
YbhPp1+vRS2y02RsdJt4PlgLt09nRShh4iiqltSGa9P69AMm6JoZ0Y77hGTaePkbXNIm66izWbE/
x3xmv7MWfmv3xq1ZPSxhRWjumtEjET3OA0klp06m58es9Rpv4bayDi7pqnKvbzrJ4In4qYvb+cij
hXXgRm19QGXfgt9KAJu9ofJaDif+Dw07QL5ksqSjcC+xyQ5b0lDvYO23Uy6wtZk+XxUkMTT+Uz+0
yC3sPSpud8uVRXeq49mSN94OYYxgD7FnM7cZmxpc9GLRsLA0P9HCC3NZMsimO24rZ8pCkfHM+0dE
ugS1Zgt/NKMy7pun0AXYw7cDizk44Ce+9GGdEjF1XdZGxdRLru5Fv48u/Nnwv5JpiPE+X76mwGtA
ivInpiLtBVbVAUTTuD/bxhjHH9VrqMPmtpMfJE2GRTBhfJ3rgQZ77O1Yf5vTH1RkUzogTqYaaisJ
a1K4s20cqqvY0sElFDP9OHSo8hTgyTFYW+S9rtqNznKHKh3OZ8aGpNGhCb98PWx5qg0bCBUF9OEw
GpYn62QvMlqd3NpxZYXDA3XWs1KOV6sHFsPZcfP3RsyDPz81VYj/Kn18eTvbguPw3K0F99owhtie
FX4THJrb0ZIXZYfe4AVqb9+SOJwQA0J1oKY84fzyurVgh62+IiRcBOXOOsSjm9ZQ+DAVLL/P2x6z
SCseKZ/PT/rfAtBnCH3nf6WO/qipprHp7561TUmQ5AO6+Cj/p7rPyZNLYPDZGwpW/AL/9uls7EB6
fkGX4CZbsw51hcpf/w2Dl2afNL4iMBVp/kkm2q2JYlyQl+bA8+RGqfRPD3OtqIpudbklgC0UZhdz
a4NNG1CYumMhh85lKTDQonQ0aYp+ApKPdO24DTIScnrvFqPi/J0Zvf0ia/yM+8LlrJVfLetzGV73
FLIBLjcjjPV/4jvK23kyeuxWMU0Cf1MEhP2S0nedT0l6nHPQdvU0R+XpzVt5CEdkJA4JFmtw00It
TSBRMDVFlfjrPyrsAXU1qR0mf9/mFaImiuU2542i4tti3vUz2YRZa7DL6xLa3drBBYpDprHcBQgf
B19mXfN1fsnfSzB0OVR/HFPAxDy2ezm/t5qSkifqvYohpVf6LjCcJrEqjc2oRJh3DZIF9MYNaZeM
hwNrZCHsCVGaeYOv+J5xdH+AIjvTgDlj/X2OTm54H9uv45CClFI7NwMAdKQzZG3uyWp/8E27II6V
lEk/LdooJaaDNptXtDCfE6Jpfmsx0fhzxRAVFjWblyuJsaJhSJr0RrTY0NeavCrxP8JWH5ozysfv
lYO0mM77DClsAWMk+Tg3VYtDF6h2GKCWOiJSl9/oVFYWoE7F1f8n9iJjg1vEkWiOwxPESHKfGrzo
h+obCO8jVSPkKX6dtO7QaDRn0D50udECwfVaPKCghRHqOMFDjoFLeWvtig87Ww6vcmPFW+8Pv9JN
fJNVW5SQUpHu1IknZPxP+amOF0mTnix9ylODI7Ck4K/XcY7geRVfSFAsQa28IxG1lNNMbp8Anzd4
Ds7lqlqI3yZ8e6e/jgBNjlBvu56faEzYqCeSwX+8lwZSb3WUdPPZyllHXu6tC5XZPbjCRAvqmljp
E9UpjH/0dSncOI54vS5ON0apxJPjb6SFRDBv37pSvAu8r1QD5JGF8FxdrBasPgDdhqR15q64tt6J
eZZG6EbJTeWVFAdnQXurJIfk72MhXeCNYiitfuVpp630gQwgYPB0tBks9FndInGih4ryYmJFCSTj
VUvwfj4oEldnqrKvp3NOWkrcY92ZP/5RCEvJX6UTxmSClfId2IiXMB3i0JIJqFXl8+rvrL39rscK
EKjfm7XkViWO8OTHQUUnngZCZuGmYg3tjz5toMM/lh9z5VAb+ILVxTcipIKEnV3wWpOJQAk4c6o5
Pl8JmABRFPrdKQv173Adygp2tE+wOD+fyQfxG2LhJWcI2KjfItX9HnwjaSo7WhTb4JnxjRtn9clE
FG/O+2Q3TNhGiMqASzSsxWvEYvOpEQX+WaE5cY0MAyFdtuZrNR679BBODR2uvKwmccDfBew4hpMh
GXVroNKJxIy4r4d3YU2dD1B6XTIvfT4QaMconWfFZl7btWpn9H8VM4Kva83i/gbsEwiyMaShUvaB
3kzr/TPvY2j1sSu2qVcRqy8CXkO8s0YLxoUyKCZz9bGC7Mnb0W5gt/HGl9mngDmPAtbbS15ThsZR
hrknUGcWs6/7KDRDrHxupIjg2jzcDFDkWwqP6Dsl8Q/JK5IPaXexknQ2oZhsbP2uxvZYD8aRF98s
6cM54rV0433I1Oy+7AoDhVBBkYXUiSwNlEk0Za641FSsYIm4nTwhiL4DzMFruXf2hkT9Q9YKcYZv
We1TJ5sC7DuPcuQP4S14UZq4bmFUxbvLbD25PAYeDFu8A2ljA53XZgeHxHbt2jHU5TiBDpS6MtZ9
ZtfkiYzJEO3Lw0q7xnvWiWxnN8LbyVCGZ7yQlyqnKrgyM0LhqcX6w1xAf5e3SBp1Tr80RsllkJJC
19JHJqK6XEQyqDJGD12+CFfZS/VPWX0+Xyku93j2XOv7ZcIbAacm64EA05ovAXoQbJPyR3NF9gJR
2H15ePdpjLBoE1LwrGldJZX3C9GROemarxvezAgX7XDVIrIaDiiBKZwZzvTggp0716VcxPtqoAyi
u+WpK5xZaTCpCi7ITYAwl1JkP+X2zrCNYrzCON9wEufyELOYUOEKRu7ns6pXcVrVF6jdVY7EEXmK
3WwplynhtRIfGry6YNTkMbZSZkIcg1NIcRhobtIzZxWZoP2tj70NLlP6MEdZqlxRHyVu0ou5nSSS
tfk+TfurW0HMwEQb7/BtLaKGZsBV5Jq+yDGq/mkSDqkXSK0Gqwv8pV3JMKCfUjtg287A5C31GYoo
BNXSXBJlQl4zvKd16A0VFhRF4a5g59C920hLJbTrS2/H6sDALHKAdRqnOANHPyU1ZQS2mmjHY8QT
3agV+V5VVYMd7gO1YuwXokP61lJ01/Z5vSlN4+Q8OY+mkthSmPuV5/sKSqWYjNkQsWKvnHRZ5C/U
agRXmOLDjHTc1+7UB2c7As7DxIQG3Ukq1flnVX+OmblQdBK3BfumMOczifOWzHgWrYpQdYulfizR
aJKXYp2MjO3BPQA3PijxbUq4kMWsd6aqC/8OUEeBSv+2oNJbAoJnsQMKehr22l+iYTL0UjsMS2kJ
/yCxES4Lh8GPfvBEqTjXwlOEuIB12hjtFzXCaaII63MJpQXZF+J3kS3Cx2GsEopJuFHz/2lgaFCb
XgC1dv4aycSSc7jtWd83CJ1mVtiBy6J61zDy0caHSjR7GFIEz7mAKqGBXmkPN5vqPJX1GcWCelIQ
w6qFn5xHLbQHUO/jbuMirDdZcD4ZbRPx0Wwf8FXamN20HjVBLThP0CnG4YDdlZ11f+YbZ5c8xre7
3WDCHVQQvEWHdMem3KaZDO6JBTQ+MWV3Hbt6Q6iWjoqFpDXUVcM6gm2I5zocipksiXrCA9cNQOl6
sNzjASK4YnnROOUIKgKNoIHS+JJB9Bh7wzR1SuUPX7tL8Jey643hw1d8W2rSQiRJRC3klR718s2M
5urd+LY33D/pQtvnc96WKf0Oo0AZyWdEyrkcwq2Iz2dtCT5IJTa1x7b8GtTE13QtdnESFwnQo/0u
nGRf3wQPIwzUh8zIhrK/f7NxkbbM2hYJg9EaVmmq5ZMa5RAT8x4H05Z+WvxWGsiV6TFIW0XQgZmA
OIcyo5LdktxYiIkUWZi3k+6bNLTio9StiyTS8Ez1O0IoEMEYwGOryJ0hlba7rFxlRk7QfJD9MEhz
NUKhSniF+4tgjwPU5i/7/5MI+e9gnv8xsO3GgSGHgUIWSr0bD1QuXtTh3zUQcWlSwgchAJ5mBqOL
J1NPp4uuTYYLo8eykLcyOtNAeK1klRmlJzOi4qpxFPyiWPxCFy84VjS46D+msBQ4c98Na3d8vPHo
ub3rV704p6d9eVSCfFYhH1jqAgB/ou5XNyyLCwUEj7ORUdojHavJTBUOEuPZT3thX5KZJWTNpTgS
9dku1cx6tTgRQzCkYCl3KMM0YVBdz5o1wMZ0PmoBSFXVv5a8Q5h7N4S90BEzoyEEZncgOrVMp8md
bq/T+Dw+gf+FseiopUFIUtFxTc1CU9sVFZ/JnmC6UjIYnu7ffpzmX5qbAFyNfudQ66gMH9m9cA01
eouwkkSzmXRW+JT41p4WFRmQWAQ3U2I4tc+wCRuz+AHGqVZl2vfCI4Qfpc677D+Qk/sLXz9npiI9
OopFl18Va2gS59SNkp4a8Ba99OXIaO25iymCNAvJXeplOKE6cdH118NGbR2+m2HWOGvYy+qIBzUF
MrKuOzAoCU7MUl9ax+UHurX4ECWSZBRYn+tpqzPT0/cwSbUqg6NM6/9JzbK5nielr1r9i7dv5+PC
OTvcbjlXDK4Gd4jCOiMhnmvTzOBU7IjkJBMwUE2ARoPvAqRfVbP56dSHFD8VWKKsT1Q4mdLd6/7B
scSV53NItm1sAzr2YwAAe2WG1Ms4ykl1BjR+TQNIeRPyGHuGzI3Ap2gNAPPL1ogo0AaiZwKZBCnz
Gyk/AOeldEiRxzpQssyWo191ZdaL22d+5aC8uZOwmxKKQp4I/JlpW3kF0OMNGV3oPxRRpkePJM97
xMHvaosturEfKRcmZ02d6DA9sLaXyrHHoB1ryOAgGR1AKDQhMSMH7Za15sH6Yy8baXtrJj3EdtdO
fLky4pxm+ePW5shJdawzzToi8gCDDrExVefUfaH0j1BXPafgPG3mwabhnOnz6DOkc/ybtS6SMKVx
hnaZzrUS8AIkq2XtniGD4oIAG4eaIEeAYLyNLdY3M0RUhE9oL4HmBR8z994CqZS+s7QAbVxvSzwv
JG2eqJaR6FQJWPMwwwuz0CKfY65SiWYndEGgF0vl+Rtn0+dN8k3gEVUyPfsWVFVEnszc6Ircsvlw
VlLkyUsGofxt3MwSg3RjJBYmM1BscCaGaIQM/gHqxs5i7VZvAFX+FJjoFBKxp9Sw8IjDsMxVlR0e
CZllsoaUK/uPitD4/WwMW2jOriSn+aETAbZSWKgtEtx0EPE/HOs/zOnvSiXF1c6KRW5LdkejERee
Y8kXfI71wr22efC2CWTKMlGgTo61+ZG/VSaFNHBedYR6l8NiklA9ccqqHqYkYWOmgDXHiVX5Su3Z
pU0EE3wqX+pm3UyC6CSmEuAeysO3EHWNOv69mMNfQnfkzHMgQ6XEvx+Uhz+FTmClm2rqrtBRPnbC
qORqJWwKJOCuaathTP5pofJHN2mb8oYqznvGBRrP8FMPOAzudnvkVVmGIPIfW+lZ2uepaeHzm2GT
4JwZQWRpIG/yELxd2KuNGYHLLGsDu2f+12YYwSd/rYuVyc/OYBGrFuQq30zkvHNIG4zVrJ3kARDp
SlOCyJpI0uPty7om2z9eSS/YTcloyP4WGAQaiZw1ZSOAXFTaTpfZrQOBZLYXagqnBMzIfMS2QRg4
vpyTRqXzCtmQvHCrmTp9gjlhlKkOmAcE9SPn5UYruxrRXWm+2k5GbFlTn+v1yqlnBzlnrYusXkL7
HoGWCpQA4Kosn6yGXIqWXzjKyVJGIhRPEEjExrdWAV97bF3OrF5goXdflXV7A0UXGadcxSM43bRk
Y87uu9vWwJf9zZM3U5auHybYWWIc+hLSqg0tfe5nAkddSlJtazjBum/fJ2LQNZWertj4i4E5HMat
AtDax5+4UB/VVK0NJPrFHF9OTTMbIGSSC5SBXupJXADDwmCO8mNrY1N5zoHaKcmdqMhpbk3b6XgS
RhszWp0Stxm4MJt2tCkXOkjyLgsOqZs2e3lc6bxUbNtKRduXT44YlRYTeplOVS3Mbt7DpjUQfT0e
U0nXllXCh7v19Ar1a3nX68W6k31gcwK0T1dO+rM8V33zel6gUzuEMy5Cd5JluZeVfoU9OI8woUTL
v5LN7BOj6azFttzPZsu4aBL2YGGkodyjEr+vndlIkl5OeIECLqDylZDijAMnPSv7I1MZTABakxhy
IdFWNjk2mEEbX2JCARKh9cEFq9w40zuVm0jEJaodS3eGsjk2Beh43ZJO9yE0rR+T+/Fj7sLsUFC6
VvOLg65Sy9IGhdyiRsNLiKPn2df/awi2F2bhcy5BIczRusIm1SwMwc24o0s1vxCSukkxAQtAyx43
jD+7TVIwNUh8EzAvifxPE2uYd43lPDf/zrGWYQEZiAtNZVC8amFUQTvETuGyHU59Fl0Wqw/unqKW
letqIkgOHQGztBPnebFoNCt08vEPWtgiDJBszvUxFFKjgzf4Yot0s6LLKpR48YxfjD2grFQtJYwJ
vS9Y63tXH+4DXlpvkC+0pDRwQaRKu8Z8fjV5ZmIFFqatKvzjOZGrJ3iVRAbKjQmeJmNXV738pU84
47VomNgLTiMtESRmL8vnerRBGWqyyMP29i/gW6qUkvfbTjzUY4Vn7NVHd55zVm80Oxdkn5g0C8d3
YDojvzsrwtERnPKiYCJ/JLvXtKbW9/3SNBHWhigVWb82jpe3w0jzjfh4C5xYZCv6HtLe77c5Iats
aGWucHRIDTOJZ5WJ5oFViCtcaFJesfhzLykDEIAYnAKvbU1X2rQIUHdJfiGy7oTQA+8iVX1Q+xNV
qbgI6+3/gysmXuQgZV4dwP8Da1SB6pQkL0lmeRfgAr5dmYooHzcJH5BWnJlqejO/UiN8FOqNGHl6
ASXLqr3Gej0Nak5Bu+wqNC0mLVl6jiOpSgLghSrPtMu33Lt15OcSYQglSoxtclsWHyw/HFqX4wF7
RA/ipyC0spp+L6CUg3X+OArjJtKPla8hKpSm37QdXWPIO/bBytpmHMpJtMmHFuhqVZrz6ZhVDRrD
VL6yyGuejOy4+PK8VEv7EEN4T3AYTGsdK4RI8/9OUP/ZGqS3gsrFvdFfaE+M47wZXaQsoE+U0ANp
ZrCtYKzbnYn5EaKwLvx5Atmw5oSEFwbSkfB/PBWrggv01n/KqI2wHpJMEKJ7zMKIZz/Xl2XU7n6+
E0tSmaIyp5kEK/t8rO/4+YjydNY2/adZte3B18ncfkoJuWH8NgqAgGzA9Iyr515H19T/s3U/Xb5y
NZZtqvj9MmcZgEanQIVqyicXYjB568a+W1eFuKoXjQfiVursFD+b0gRbVJE6nBShzWSIHZlvQKl6
kfv3d2FL5JMCm70DUZKN8Dig1LBgLqsTrm7K8icV08mnx755VcccnvcIW0G3GLSmu0rLQd0XlFIu
JWklPJSvlVkGfGiv5P9zAauTBuaM9wlNNTgRpJ2/CBNiBzGZGeHcq/Yp4lkFK1Dk6cnltV36NkSX
1MnkC3+X787V7za4WCqwSdwI3T42+U/ZX8hIcIR1zlEALgnxhPVKd5NVNCSTDCLmTSfC9Pk8d4k1
mXDAS2Z05LPIZQMEt4avuYmWNkyt9auF5GG25Ysi9ROP4AOdQDpNOonW30pI/l57jA7Q+VbZLS1r
sGW6NlHNP7i5kdnEFJ+lcpSiWgql1mcNC8n+s/vVtRNz0yhC95rFXq5kkR5KYdItDog/NRfM5KRe
aNifmgmi4ZExMafmt09z2eSsPgY3rw1zqtPY9nfvRuYLNbgnHTh31V+KuDdS1m2w9PvoS6wnOoO4
4fPVZuLxnX6OZK+SOvEYOLDzo9pl0lIArvvOJQXdIrwoYJwiMj/QtRdX4Mvyo13695kWOt45TONl
ilmfH2NgAXfHMzlUVf0XxQN6VIFaUoVx1XQALrZP+X3uRHOIn/N2okPPIkEv8rIpusnR6lcsW6/h
eHPyt89c2NLZ0k0c/AQPEub6fhJ5yTjHtPwG/tA4oJK67W1avczAIOdLTp0A+DTNRJ5FKmADyML/
hvAK9wjAB++pwWfBquU+WpGa372HgE8/Yz0ewmk9eQmoH7QGnahV6gpFzQcvl0H6PBfgQMJqtPFt
YdQggeLSASPK7zobvubdbaDkCjLwOzDLrPXpWG+C74bEZ+1zRDoHU1ZNyH9jEh6LI3Gl6wrGOoJ7
PkbUHHqOnW942ljRv9AGDl/KQ/nDDYCGsQfeHO+aEl1copg3tBg1+Vr5IW/GH/6kHYIeI14m7wzn
e4mW9ZYcjh8oJjAqrQu1rswTg+pucVZw/ZkRxfQkBp9MMNlyR8nMUdDrSPI10D0d28m5MXbgXNSs
jezMOM6oQuf0ZZxgEMt/pSzNw/oJrd91pTEq9ybdj9r/ZCHpbdQctFtmh1uvIJWivpMQZEEEZpSB
nfRkQF6EVGf3CBpClTsJhsnlyPQ/3jNgOjcE3ysxNOgn7jYG39+EhGjZNKGi+2xtpcd2tYkwK3ne
7rYYkjfrMBWdl/Z3mhreY3ZOIOvLVnjh4fJ+8RxYJx/vtmRHuA3IoGKFbMuXORkAEtQlB92SPq3h
+jRyPYt9cVCWn0vXvPUsET8tL7LYF6N5xix5H+QomFJDvOab4BW1zL/BuHHn/IV36rHCuJelN4Er
RnmicLroxOG4ZaqBnInEHaXjzrkxmWArwsyClPYNd7A89loM424w8HgAChQSV0v1r41Xq3SL/2yo
5fenGII/77fzz5mIvs/+q/jWdEkdvpyqIqV0sWG0PpFjhh7WTTrTKYrH/b1CmV4+z5ghleYCOj5k
3+lKzDtdI7HT4WMMAapdB7JypBMO4aUrM3sGu/lAogmLyaJn4sgwpD3jQZ9VycDWrYh/7QXBrAqv
GX2uyh+TbR8WzKbDAEJosM1Ekfeb/Wyh82OMuxJGz6QSJyAkloZLlND3pQxjyqlRZct+nZn0lHi3
7f1eZpoYHG3V1l5A17leLvoAs/WBNmyvcBiCRuK+SBZtLkj0RZrmWpD7KsCN57h2lNiUdtRNU3ww
jjyycuWg2fiFRhexUgvG+wFLb51qRCZtWHwx1JMAFYohGNy3ADFbFTy7N7RZvRnl1B9lO/HX8DWO
rX9TEs9QSG4lN/7Vh8TbY+U8Q/eEyC/5LMYjm8YrVM+GNBtXiDy/tKLu7/RyBoNHnR/eu2XvwNp3
mpywMYJFnSwDa6Ma2RPY6goRrXXDAIznFo4DJ9T7ustlSqzDruGqF+Tp3WHhq2ilOrLaFFrHvmOs
dmI5bT+L2HKv9faeZiRleoKOY0sUJm1S5fqazy5ihLxjuZWZ5C8fc8niH3FoF4sctcH9NC2sgzYN
WE+19KmOAIcl1Gucp9PobImZkkF3W0sOpp0TUdKKmS9GHcJ4Ve+DrL2DlKpQtNj2/2sb0QCZ712E
7YjGG+rjxkY33znRU1knLnGWq7a8locsCngvMhkgHcw3dHvc/ZeivlBThC68Ae9TzHQ4pK4OKVZs
XTveR/O9Z28cu/EnNfzUZ+fGlUn72yhG/50ZpAv+veFFsMhZjO0eIKmU9mR4bPB+W2XMh7hkZrh3
uWs4FIepMQDGcsM9DcFmjQNlD23zodzHLX2QVAyEumNM1+g7RAb7CKpE9cav6tjarO83mNlCii0D
f7qhK5npuXe/ArV9Ydzvymkp8pWpnvyNx12Em20HI2DSBkRPOuaaFXqNVAlp4HN5lytgPrems/I3
vTViUoEJafS/CY6eRWFgyJ4pOEmZ5ffKvUldyzxwbizmdSt3CGHP34+Z19UeZg3+I8JMRtIPAHx5
QG8VFlZHk5BVbFsDv4ZsRrhLlUmw5JHwZtzKQFBMoNUmR0jkuaqwfP4IZP/+NK+97H4egeMfmfMD
NH9MR+p+jzKPbG8dYUvGBJgfQJ0Ou7nRbiEZ3ASJUqYzfd5tcJu3GS4ZJ45M3IWMqKMk1MHoM+T6
X7tpI35eRhkc1zVgVdnaEiVwbtv974OOIdw7xzOV3UPIOyo+GUN+3g/zMjvjtduS4bkHGFcjlAEk
lxRaIDWbj8cG5V5lStFq8lDqQrYiZ3u/6NMnjD4y/+J1aFPcGWQH77pkTp6AZfJLLnTiL7kh08bG
+/wZKxXbDlxpXcffWCe7RsxTJDtXUte/fYdJxQg02J6u5WrTTe0CixEUYhmd43ktiQcYp4bFSKaH
tQRKsPe2nNn5XYsx2Os7Bn7A1r0gRZQFTf8S1/VWAt84Hwu4kVPZRJia6K+g5I2nfI6BabnUHFoV
L0vtmOksJRUFPkGevT6UnjamEC9MZsYxRkBr6WJk+Ud4XkpsIy0vnCG+I2v5/dWh+wAGpyNQZB+X
95s02aVnWADUQD+9e+lA+CRcfT3tKx8JKwdl5WYCMRJswSUYKfWRhRZo37ZEbexOcm/FQJqdI+Ec
H1pJBeIdcigpnDHJLrqp8d3IN5/PpaZLdXPRS9I+ybQkH1yk6OzolkLrRwrDQ3oq7phIgrp6zwH0
1WPNZbTA01l7/XhsZUdOwmbiBiSxmonOC7Tn0O/DqO7qt/6iqvzgTIGdQJNtdA+47lj2FXoxCu+6
og68cfQhmKaop2brGqRZB9aXkSfSsFoFqGyTqjB2uHiefo/OzNPlXG7Cz7Sv0MkSVwEPEkKSneie
lHog70YiBQWLVKF9Il+x4mJVxFU5gWsGrBD6Sth+LlV0MeJeBIarUdyC00Sx4GYgair7SneQCyJS
VXxx1junZYgY2zVWXCbWA+Vo0gJpf1500a26bY0nLOxkTA1dett1aDj5D+MRVe8Qa8tUkICBwwl5
A2c/yWC4EHDr+/0JjuY1CqT4ffiCoYjNryWV81VS9LL1R2/gPc4r2jAZP4Sbp9eS/Jkl0xN0EffA
+HaQRcDO7pgwolBke7u7anMYsXNVw/ocGc9e+cLu1ZUSvO/UA+6pHZ5KDrsQ6cvEwQVqbfQgmcit
jDw2WCDL3ybV2E6nCIYYitBcvX500MMIJx76CBkw8Qjyx7VqiI7Yi0593SbArW9+mWB0SQH+lkam
aCo0CdMGjO70jjjpexNFbu1AwgJfcL5gYbBWRdOOAvxghDTgvwJPGfRejynLcWS0Gja74D5beVOa
g0aJHka7b5GJJt6dJaTzT525ZlC07q7UBwc6G+qL5Cq0CGU+mepuFpBYhxKAxtWKjXBkN6XED4gm
F36s35TnbM+CjoEUBNX5JOdqH1mI8Y1+ilbNDAJgMadzdEjKZ0KgRrW/QfPGMudY5iMz67pIZK8B
tJaKhqCKd7ocDjlCG1lGw33bJ+IaQcdqbOWaVpLMv7UAh4XquZikNjxyP4/SQ2PgOkiGHjTdUwnK
Sol7o5FJ/bEAWtcf3o2BdibvzuX1B+HN60vQWAZ5ntmUz0dS1kLDlzEGFJT02Mlhl5pM2+Ya59zQ
muh8QtOZUbnuOZKKyt7TcKo2d7TwEAOswZz+HRZJ3F7HjXFGUmgx8VuKZNFlHLP9Q0e+JRBm2azh
ECBuXG2T+S1nqbBO48BemVohDSM6363lgQrHKWLogiIMIEIk76Rs0LFy+Ej987oXaviA5vV5oaoV
j9hfR3WAHQBhnBoHPADV0MPPWWRJB9cTxIJiOmZk0G8CGe+SofS/IQYuyCded4QENh8py2olRcLB
7KqYxP0g3jqHwtszD41J/L0wUXxkct39YmNwTsKSYkHrvHooOIDW5XNX5/Stz2ux38sfkZHCQH74
AhoAkjrxjGY5YVddGx45ibHqZFuC65qwVhq+zWjrVEbJEjeJqSCYA12nnvEF49N8n3L8vMVYKJSx
ER2O2asDb0fUKrynGEbYY0d5lGSanPTd/XADI5Jd5IWsPIdStg3zm3FwhFXnEsE+sCIGxcY1jZap
FeZczdF55hdfBqpkxBwTQriRf1n6wvVqVysfGC2148cgaVU+hm0otqACjlxSd/Ti3OhZ8P76jtcp
TEhx1lNgD9Wvi4SUCrBLtYvagThVwjzN9au6iDY7FfI/48Aa9vO1MEB1uNUY65RigTGvIKQaEutH
wsK3vJS4QYbOtymZrl1hGArJmUrZ8NVY6Pf50UhT0WoVjLy5KIaRU5orcOeBCz5kRNYI5Tae3apQ
dTEB/QGL2p8LTd9OJr9Ei/ETTmhFWiTf/dTBAYpVxDpSZ+l94sn6kPLrnqd/xdceDAQBbPcgFtd2
123bqoVSOZ+jn0Bc0r3QdnKgn2MYFwJgrPQWW4PgsN0RfkI0YQA35fVgqck+cheOpVRTUNpaUaHI
Bu2FfQOysAFkpgnEMdR0xdUp9VEj/4vfGuu+iuCvqfdv3dk3OwpkSRT0RsgN+zeInf+T09Q4kYxy
rz+QLNLRro9WcDsOM4T17r2fnS7l+3tpBiV+VYjnn3laYTqBdm+4QJKrPpVWFNHVZNFAaVSJBIcl
4IV548NeQHPiulpjsx4+27cbkCHdyZycnZyvCoPF4i42dJbLaWBIRgVwP3FeOfPBx6fyKlawC9SH
5cUldZbXpfZDVQZePL4VZYxFL804uFjv3K8oW1yztnl3v4HpWbcnAgzZ/pbqWoFz2rTRQqR5qb3G
fKmXH5TflpT2cludqz+XqFcSmE8h0rBkvAUpFAib02uI2pZzIHPxHYyB2ZXY8rxtgoAffocJU8cd
cOx24umBgtJO5byGs5cDvWPU7ljCzoeKQYSO8Vxr+FEDrfg7dcZ22ziVtqMTJ4UaKd8KKcEjl+fk
YjY2x57QeHWo2/AEZXwXjtmWW9NnRCqGtN3luxPtSC+EPxBL5fJsWgmqU5uuIRnVPkujt8JHArD0
aGgG0NcsKS85Z//O5A+3RpV3aAH66ISnkb5e49xAldQpD5wHZbwR707J2CMIYq9QRU7KBdkYL1In
sHOnXj0E/eUOW3n3dxwkIMgb71ZUQc+Gku4w7fN0/WNZ2mPMDejHAwu+MLoK8hfd/S6sXNqpo5G3
11mjWpamAcGsyQCxBbEzDz6HXl/lJx4ETi6icJvS0TlBXnQdZWB/prmibwuWMdh6FbxZ1SZpWTQF
xyHIBdqx1fZFjhwFFXcpZ7Sm4UMlpN4mQbNlSxAQFt+SvSa+gRtABfRaLhR2+919W5DJimoPDzUL
nM5OCDrdFhizWdwujyETLfz5sldxpAZAbfdJfdehs39BvRp+ebNE+7Wf6bmrl46LOMOHQLjpiHcg
sdUvEyhm3iGXni6tkZYPDo1aW0NwP6kXf1YWaJqwImqkKMzDdQjdvERH3tmY4JX9r6mkEOwW+FUg
qrBdmSzzJopRIIo4pDkOsw0g3QNzdSDE4TywuyxfFYwtHVi/GJyGZgJvKdtqGFJRveaNLf1kqI28
62zhubZbumBL87gHacY4YAWvVbAxBSYjU6KK0xENIpAZ4Drzc3rXAC1VW86wfzeb+GS71po1BApq
EsDBc6/amA/CZ2GvvF9p+Jyt/f4cWIkotJlV6mjWugCiYsuA22hMA6LYU2NhtpW7TzJw0np6MOHu
vwrWpZxAMRQDYRUl+uhiQ9iZ0UyoQSux0S2BkJj3XqxmSe1B9xa0e6K79UM8FhaxprOzf3GM8yDn
QE5OwNDXVkef1WB1IhchJoEgAjwBgW8rv+o3WmY1LNar7DdJW3e+0G/sw6ow2TGcsuOo6GHgVGR7
lVoyvjBNh/uL5TpSroNdOgvIFkwtOQEIT6swnv+Fb7sB6zEO3BdBgjxRLNjOiHpnNc1F2so7eAys
H4xh08t+OT19SraHF3os7Dp+UkCcPVbyN1AOflLMyBQQNjM8MN8D+ZMY47o9b3MKCXi4z58qPyhu
QciwN6WiGnXt9u7idRvs/PofA4Hg40tSCmAPRMSmwKH7d7Qf7q3tgAAKlmvjMS4FxaYzJZKtwvAy
qTXoFCXTwfThJq/pyoMOtHxlvnhbwZvSCWBUS7WUjUq04RLFQb2X4l53NIPr4a2PNsqAlXwubJra
NWLTrmCu+QSo4BT5ia8WzFFXbdzoeIsoUG7bplxQeq0P/yil2Gg+b8jrklFF7mDa4RTRtlI9Vosz
VE4/3sew/SywtZvEps9cja9BDUgQnsG9wVKOuv0l42DZOJistygXpo5hYaS7Y7TpX85Rhf8c1CkN
4ryOwLiwYODviEycPO258b94H42LTbqQ50Rp3M/GIHz7nOwzaoOHqWKhsSxzIl27RXPLUwXBzGzT
bw8sfLhtaW8ep0jcfDPWj7ZcqAiPy3l+HdfBh5FBCPLuTpmts6I2DKtH21wPe9JOYithA/7wS3XY
DgbpoMLwRMzw7RkRN+Aj0mqArM7eZW5x3SGfXw+ldLEvxhoytOh2l/qHPztJgGM4G0H1hdTCI85v
vlNZCCFvHsU7UWn+If19TwuE7OwvHCDjL0llUWtOftWOoluQ/nCYVXIS2c2BTp220SN7wSfjBZ2s
3FkUsdIZ/STHf+37BdyrkD8I20SgIyqdy3+ZEKQP44o4X9Tc9oAFv8DuxJq3vxCegYHODSq79doi
ImLqL1aOfHwCT9uHoEafDaeojHlYCFE4EOhm1iMfNCgyEhVfsj3D/J+LNq1Dp9yFRb+a7Y9zZvdh
77SwM8G7vTPhjwfyq+daveM5jaGuSX+3KPSBNrRNXa2Aq4qZxZgh8cEHUMW/K7aboa8MI71jI8uk
xcYePET5MFQPTEuUKXI5FZxHN5ErMLoo4FR0u9++H/5Woww4vO94OEn0tzn81TuSZvlqa6doBWOS
zZTJBsWQpKhuGgnrEsVEw9WZuqEmzNKhcDsivqdWpnozG8PFxU5ZVjSEuW0BFZwsHTxiWJU9ECVw
jrhDEIyl1GXWYSg0+973qC0Ii3Ta1qYGNR+oamX5DuF/HhNujICdbendXnfnNc58kEeUkplfDSJ9
v3MS5K4djl2bWv7sQuHYfTuDa6nTG9VvAkucaGRxAhlMndMqukKTYafqHUHEP8CGUxYvABOnWlF6
FRELQBpYHdTf/JuRuFJPTG+/Z5oQK8F+VAD4U3gBQYxg0xJ+p70R5pa1c1xGYcxFTr2kc85xfdKB
oHI4E4C4mfHuSVlr49j+pMkVLfx+bXQYPLF0pqodv6Tr6lDBC3UVec9icyyowEtf1em+YysjxITk
BUs1ccxMMVFRaabgE8da8KlTshcHx1x0pB2GlkFj9ztTpa7wA74OepNzSuTp+naqvJJ2tNDi1Hm5
JfHgxWSwBbixAaN5mx5TYQaQ//eu1Z3y+sh6PHNztJDQdjTm+/cu3pxKROadjFQAK9uIZ3fq8XvW
tw7apMxriWqvv/cC0Qvz3hx9Vzyp59RVAhtSQ61xOPH/PDGeDZu3wcC4/fycFcERV8mOJ2ME6Jni
iBIISNFXeaBGx9MssShdnGKiGaiE++kFHA8OtW8JbqbLKIZO+PUw9fLlQtVuLmlVyaXFloRWqbWw
Jd7Y91LPUZ1nCKTmTfE6CaTS/kvdwCcYZXW++iv9q7AUsjKdA4OtR0pYviV/chQl11oiMYe0I9N/
o4GIZJIUkMzA/VkCRmztzRtNKHOZTFTSLpXFM50NHnRWnijoyNahZSTsGJL0G/lzY48z//j+SV7n
ogOnpU4qXpYwJMPvQtLJNzQGHy/5Cd3jUf/96l3xCJ+Gkgygvu9C76jrZ80FBmRw5uLOMGSbJory
2Hx/IS6/Pdo2LCMfor3I5KiCyd3+wuXuL47wizMEiyKAXieHBOnR7OGx4GTfsy0Is8rYcPHrQiOq
16u3mIYeA3DR6vxHwrYuZ8q6DGnNAcnmodGTKf1OSPH6l0RDAtXKomrEVCl6Utn582q1mkLNuCS9
n/+je8jOSo577zIgGbCcF1lbwW5VbkI467I0sEvrN262J/d6T9bNTEA9akF5rPnZVpQvtQxdqVok
XhoXbOfeirYv9g7LZIjIvVstqCFtoJUyWA0b/LINDgEB2XwfT5fP7rYoEPhwwiS5+mpsW/MJX8Rb
pxaufhEZS/flywdkw03oNw90d0U1dGEnSuo6K1Yqy7ebz5c56QcBgbU3m3FXdMTIeykogl5OIJJk
lhjgPWCPrQB/HTcPs+TJNex3iDHlZQMSqB3PxcEGXRmZP6Rb4zhslFUS7764h4578AgggabwuBQw
FtRT8MBoz1ZxfpPvWcNUEWzzq/V/GFqQLRxp40Ok/prU1GgVrQveeqV1OdaDYbyHraMAdhjBhQnU
EY6uj7BtJ0cVYS6E7OM202soKZszhuuCHyno5jCJEv02BRxPhf9aJ/szhTd1idY0/wxZk7ZoLjL6
kQAnQYvf/+px4eQ9y3v9StLTPIgd76445UhRORlw0wcj/RqxGgUkgfwi8PkcECz/RAomeRYkz5jF
Yxs8NbAFX/EnAWKmTrEkfkyDC8WaPKbq1J2IjCS80FEXQucDQIc+1XPBV8icjx9vyjGBvxixos5H
Vl925y3eDe5xQIeI1Gk1Jf6ZCVsuyxTbP/r7ILKUjrnt5+xtPIsEV8kaQRvlAZ5zhJ7jOmfoVMVF
8u4UmN0u8RmzheTF6JoQNiO6WiMPNqXCWXPZ3cBj1W2DtQsINo8pnIK3l9i3a6Dg848H3qN1m3aO
NGn+Y+UKm5a2t83i4oxjRcXk30VDq0A1UkeZndNRoRVrMT3Ws7UvnxEXF7qyDDEmlC/hld4+rNTL
AmNATuBMv2+zlr2XCVYhIjd3ZVLrl7A4R+JbFchdPRCm+J3eCJNJscQPj8+zi7tJQq706zE67/+o
YTMxxsX0bKdobJ3c3nDe7xv/21SEJQpFppok7gmHoiRh2jcairFEoVjtznaGQJPrcsIEGiDuJax1
pwdQUyKmmR/kJIze1SEMzFUBhzry9gpbQluc6VB0i3+lpfNBOPPZc6lOQ6JAR3ig5wNsoXJs3g/f
OnPwZbpEPd2W6arI3+9E53/l0ZOgc6JT0DVTnyByMfalrQ5aC5/BfLf7kYoHOU2PZ2i6YfoLL3U7
br6T8bQmV+u+9FsPKMmwrpMaW/XrWljSiafhg43J7bhw7Dz6vNKbjPdY+d1HsCkafrugYmVA5xDx
Z7i5mpKUHaufXtshw/Ay1xoy1/do94or0VtoOALad+uGjEODy8GG0z3YJHrntLQ4GDbUPTNTX7yf
z2icHoXz8VWCn1IPJQy5q3IFt4hizewSbCpKPWrJSja0iHbBIgr/DKj18ClLM9BNtP90nP+qA9/y
ynC8jc9DotwvJf/UXFa5FAAl7QQo6KQT7IaDzbuyzxDRsHk3wpOAsctSH7r6p2aQP5leI7gheIcG
svhpPvc6qR6h2w96iJ9vkBF5GRsh//vtHZTmPyDENoiTNEOz2ce9B0AwkzH3nkJXLiOkg8RsrRsf
/hldoEX+ENoDovtXUIqhLMZJpHtJOwnMcS2GxR0FEhyNQH9CQfeunWOgWXBBBn4Aqm00noZPFIKg
zXRBuB/kPyW4EJxN6QooXVUxh5izmtr0r2l4eghz5PN/DvThifqEzY/v8Bdfps/vo9Wz7Paq549O
21kuxpFHSAKyamlENhhrWKPbOQ30tnkKRL40m1I88GdGGB98Pt81uhjUYsh/MF7GWiH3N0pLUP3F
29088qdDvyW5nY7/sBknlUPVBXDAh0Vlw9ITQWBMiGHxDMJO7ik1Q45zP5G0ovZonsFSRWTOe99B
LkLmR7ZY6Xal2ZYTRQPK7Op9RE8ieIMpCO2L8OGNPbzRRD0GgXhSZmEkx7PD38EFpNthjeDuxNY+
3HDnaTokgz7XxzdeGLakKiphSxiwIdK9n/mXIcCx3QVoeanZpklbzgSdQntQixgkw1xAlBeR45qC
ZkbRQPgEBd6VbG3dyeSrIwHatFBnftDLvA0jt49jlTHwSss4+dNoCr1YG5Q1tzrteHrijFlQJtuF
LjVhPvOe9APcJssox+F7WIKKd2SVticy5MaqZkMeWdn4ZXjR7afi4cRxuYM91CN5Eql6NJnb7gyf
AQyhvjJNgMoFetVUdMHm9lxURrcTQwcmrpX9KNUR8+cCyc94mn3xF0rMkfGBbZaLqyx3HBNsibov
KF9VwE8Am5q4Y/uv7aAGNqBdPV/bss3W81282klrvS/jWSMD+aMxxoJywVKzR1dfca0ogJbRz/k0
+Sc++0jNxQJJr4luB+0aPII1lAgWpw6BtAng+W9zr6/3Hcm57JrtprsUkoDRsxWWy4aY/3UUFfEw
KfCrNTYPGYQgItKT6KpcAF0J4YSAjpntW04zbx49m6ywJMXbIIjNDzvpvbuMgjSI/0PEJ6fx+2bW
9paQkl934sbn8No1539FIizjVycquc+xrhURORtRH8AFJZchYAtbTgs5DSS7dm6sqQK1GjRIWKIM
VOA8N00s6kSprvstDJT1l+UJE7f2EvjSyr1DuYmKbS1iEo3wd9GNo86vjMf9q9tlmDsvlucZrGbV
twrI1cxhZNFnub6weVhyt4rMC9Pbrsosezw1qzuSfNGAfqTjQcVzVlpZTioAa3+Q9MXCvu0BvSRy
1SwOsKdq29TST62v8lnL2Io62h+mFOc6U51ENcYwhqOKXA5AtFKVsM37Un5BxlZgVRHXks2effa3
5tHWyagRwC46FRROiX0TbpGe/o/VlpZmVmrWNXeuLZtCSpYsrHCSVvSJh1Wa/VYF9zaJX5I2z5UG
YkiTGnnaGvFtqXST8fkc9ZyL8hoziMnLhyDm4LIMhstOI/FIMExBiQZ5n/5QQkAQRt2I5Vg+Z5XD
1EI7WuIlp++JT5w4TA6qqLtpipJPXdqwwmQLKIKXb6ej8Fug8vDmaf023i9muLOLALGd+Y7nS+S4
tj9NmjiQtmANLq4Fp25vT/bpFjAYxPIRiez61NIFaK+WeG8wJ/Q5xWNbtOfVu0bpCOuDyY1pZYse
qHkjmj0OliuQeg2+ubEUZ/R2X0JrK+YDHp58YOwjUCF1wCv0TXj9HjJGOsHTkkJB4WGcLXnyaqax
ImVy/eCDGQ3z3GADxKK5Vtwr9dUjd4IYCmZHIc37Ynbz7rUyQYkgd+aDq+gECXhGc+lKg3dHDTLb
MDRvoz6pcT+A6nfnF5tkF3fA5IpQtsDiov0IMaHXw9aG4SqWr0exf/FvMoPfdjEYQfNqgDimTuRE
1LgGFosrRvaeow1B4dtxcb7V+9ysF6spWfIYV3JZHwQaW00x9ZZKMw+Yt7PQxT4s6B/EvmXNU8zZ
wJLS+frdgC6CE10bkN7iBpaZmD9jFcdnSuqi/OiApibScRhJhc/YQs8HwNuGqzF+i7HJv2nzFGDR
lUwpEe21n8ZJNSn7AGq8MlUPac8C2jfG/oqxAms6Wc+Bg5wE76z55R7JTkmxsWW9sEDF13wcW2Fv
sb55/56TOh4wlc6FIknHcHLW1qizVEC2pfgCnJhfBxT2Uxnou6lF6pn2jgz/04ba+LNqRiaF7CJk
gQjsU0d6W3kxw28ifDK1p4ynH+OqksR3k2F/u3iEn2zI4TlKPN80r8r0lRY47Nl00Nvl3wyJUujr
gBvP1+lhB3RSoaQWcUReri1zYAmlFvxlWNbVMoR1V5xhBvtgIAGs25/L+gSL07UB7+Ku1/JsA+CN
Y7AADsj4U01/b7ydy52PWrlHTs8hvgIICfp57Z5WVKdD/cnDKvqlDrgo7SH4gwrCRCcxGuutD+DI
NyMZLfmmqc40/o0vAZpa8uWqKLpyR4n8ZZ3Cbdk5QFu6u5plt40CWJXbAZSu9bND5rJSWfWAo9gT
QpnLeZnmpT1iGIt9XuFEzmNbvhxOokfHvDuKVIFXIGQsVEnT/jx0nVaTdt9mww9Ww/yk/8jSxczo
Blqs8MAcRxUrd+su193uBkM978nM8+w5tQFQSrqCP5LSCNWygDDAwSY2Yc3wbO3vtriG6RipvTvd
rlN4tvZ+MtVnHgxOIhqRzVve9CaLgRnFcwI5HmK8zW3UQreYGJQ4g+kxo+xQl0xArt7iG5eYGs+S
obcI5iIEee5myObIsSwND/VUqqiBk1nC5NKzzfQhh0u9Un90F92MfqEL7fOJgv+1gWT7ardg8WTh
6heaN/ZAqxKAUW7c54yynylSMVR+7WAwrwhbdBH089FptPvBns2rrRmf2EEgR+AIU2qTiL5oK1do
u2xV23tcQ6bPLF0xHjOZRlfFwqpP7tgvlVXn9qKMyC/uvVLbhcGqHQzNixemfDpEU4WrvZ1MFLq7
H4VQNu4qR5lTxgKaIyLzoWJ3+lXT+xmX/eeAUFk/trfnI1n8WoSbIhJif+XmXPJB4k1eejluQsh8
/+cQ1l0AVQ33DVcar+EE7EC8DqRtCg2BEr+vsb7uL+qnsvv/j3L0j9kyjRMywrZccyu69Y/lnDlq
ZrhIOJazEpQC+aIwGML4x0hS782yLgot07RwAwTQj59vXBxl9448kKESzcDLSNYjskynelIPhQXG
e+NqjVAlvNhMe1v+YQRAE6GJpMGQMXhY964VGYuQzGTtvCslwJgemEM6jZLvVHtzyAFju2avIlgx
Wfn//Vwr5y6VA30CLTArg/YeVNvpgXlfQsZ/ISOIrvqiNDEdyc5qkGPH1b3efIH99T9KCb83bcgD
NcYUzHZ2rTOr8Y0ftadwUx+5+Ri+qGVLB5pTo7DDiLT0uJqgOkC91B2jF9n2HYZWLVf2MYFbMAOU
EkE5rU90/3d2Dl1NO/7bPb674EvEX4dXq8OSdxkfr49L5NogSN+LQjX7MgrIgox5m371I4EcMNTt
CrzWgYj5Ll/uIINc7XqyYSvxS6EadSZKX23ECS6kLecFP7KzH2Sl5qUffPy9J7PqMBP/yO6QCB+b
cIpttaRbIruziO5kQwUyYXAsIewdrjSm6JBKFkSd2CuAxEVFpzUipMNfQvwVsgpdG+AzzDoVDWik
b12A43VbAwRNmyuTp/8UsZ+gdMEhLanI+jnNNXxot9Zt4+oKfkDoK5Rso4MDA399XO6Z9YC2ZFzb
F+kLZvTIYCQi4sPwYwJO0zKADW1DH4epiPG5/KCO0n/v7C8nIAFuVXHuVB12hOsj1PC6702cd6bm
14R7XmJ2mCCGmEYP7Q98XXeXdcItMmJAFXVgvdO1ajFF9z2iAc2NG76ypXWS2+ET9sFLd0/r0o/S
vcCjJMqvBLb6+eTd6Q40ZtK/h3483z8LQZDmlZF8HOzCxH0u5dn6JXHRRS0ZCs7P0ttpgYppj0ZX
jsjIOSWteN1Hj8TYoQ8xLXEzmF/Bvl1HVjYfbQni5nS/nziOob6EuRHDyipsuGvRABINO2eUyf5M
fPZ0lMj+26sX0aBg/7rWCwn+vAU9rLWjncrmeaOit/YSjK9Ks3N9TJOwjnjYz55X+UqHBE8saxUg
qTkLSM2FyHq82rrgboXKT2Gpwm3rpf250oYfJIPRcOwKF2uJUHn+b5J33LkB8qbK75JzSgzOEpmZ
5rAlBSaPtZHVo8k7Q2YVvoFrWNQiQjLTftCrjze0o+Fjw39+9nwgDdVLULnHaGABvip312V+y9zZ
7T/cNWhEI3865dQJh/pnlKAq10hELXbVkIgRZ3xK1ulaTBCyKzZn4g8gvhFldcsgQla2N25ovnyc
LAQS1x5KazbCOtSi1xBxDGM16uoQYD4m4Y69o1tcRjy3DVP4sJqjRfxdRZIqq7K3/V/8d6q1OFmp
p0pIahyEvIpTVtX1gQKswV0yEdPyZN7nokLem0LXw5xLXMe1yfQNFbS5eQjsQ/9A+S4EKJcHBKUg
vrW6egiOtVRVWYl1FplKuPfjp9d6UMYGxG5nTVfpgPG3UFqTQ2elVjaoe4h9QobsQZWRwjLrjdp4
UvxllYLpRR5ToOoOsZPjaiUm6hV5GFfzAp7XXmGYKhnLjcB2Yph2qxnOhy3gQdB6VgTswrR2zvpL
lYar0mTaR6Gy2DjaY/mWgxPK78NEKgsw+2DJAKjSy3CQKpMg8eQuLQ5lRu3mKKgMWr2SP06fKvKK
+N6CNpSirOFI45EeS4lAiBQ2loFho/I9iHHbu89UFpdykFJSNTYbw4yN2B6lZ7P+Ts3MxprvFhhg
r4PNgOkiQNUjygAxTuweshdHcYo8rnd3RWpJLH7Aj8M33TfsKfMSn9FuxKda5NwLFxIUGEhxpSqH
2DJKj8ntsNI18jr7+x/QFmQzAB+w0JsqxTHm0RPST9IithAATH6YTFKckwefJ8PXrPkbVIb3doIx
tTzLeK01RmWI7FnAvCVTqPLSblwIPb+B4CQP0Da7lJeavJMY4EPIMIsDo1bE5gZelbI2+s00bPES
ibiqOVSMxqZX2xu6I8LIW5BM0W/ais+5SVYLcRQK5qVNCGSnnIC0qG2plav/QEpU6IXTRa7n01d6
F/DHhW3Jel/BRI7EwwPx+ZhZZEe5L0yFk8KN9I+P1WL7qLcC9wCnCnWjSk1fS1o7jnkZyYHGlcya
c5LBS4NX4x3H/YHtZiYRF0u/+lEbcfuWKEsuArKC1MXdl5ykHxSGX2AencgleSj9ua2sCFj8N3Zk
m9Au6aNw7yyJVCsV3h+fKnfATBYiy70bZsNhiHn7ujnYDEYSQzBaWtAFlxkyNYKbSLlWqZpUm8e6
j/lS08Bn+9x2vu3DhDh0/sjmFg5AVTw+UHnIm9BwGOhMftCyVVdgyJqpzvoWAAH9pZmEMX8w1mZw
XoRPgxK3u0cmkJmoxttows3ZD+kf76hevq+EtejMe1njhDWgjUKGgBNyflovtMmr6I7SzP+VGp1W
KUyhqCmdJchI5rR8zIjh30zej4Jr5SArVaJwIdxwkWJt/Q6nzvpuG2HbUs5uqBpqeF9VrEjY07Vp
whV58ifAYIf3NMceJF5HRz3bpHsxEiNXe+LlUDF5T4cI+Zpvr1Xl9kEVr8T9Y90QEWKW1eKS3X75
+ZqQnQJgXQP1VF3Kb0kIwpdwgF9tzKWRglxH1FZaoYSUbqoPPfImrKHFApXIuB76ZINqIzjEOBl3
tkcZIr480obZjLSc9yfloEIoQgJtJeKZVTx9cpwI4cLh4rshYClbbFh2wFA23BUOaKeBJa4khvgD
czt4+9WQwpnUH7t/Fn3bmwKU4Xup9mSGhjh3gYxLJdmZPct0uS0iLijflnGU9x9ivh/gRAw9Vihv
7qZznJheECdHNmrIfri2qcbGVS/dyBZ0GrtpSo7TUg/EfhfUXImWALFhqLgqTcYhVesHGmoi23S+
EYKkJ182k2StjLI/T195DcMI8OTCeNQr1hrUSWD8j6HiPsztTydhy7RlCEuv0EzldbpyA6gcDIhj
otYZMVkDSxx614VHJOjMWRsmoSLcSQGo7vfXYbJS1N2G6La1NYBIyWfBo7Id2URXXM+16MzRKGmT
1nAgCrjGxhRFTZuP884ty5xP37yWi2invUtkWQm9vQIvrHnwc85lKC7KKbeFWKFwhbahqqZ3uNQb
F3zbhE1KDyudgB80TXvcBMJ+AmM7htEHBfJOTyR34hOpjAtKlFuEosLdNqZg2R2gx/6Yy0Ws/AqO
2/fp4lac+JvXhsBcW+TcA9ElnqXVzE9rwuMO5s6F2eHcJ3hPYMyEzhWdKx0DjbYAFSyWnQGRgwRj
dJ5BH2+mYdq7PYemihzLU7bvOyAbVhhdFwyg+/G2ZGe+6a0LtidZ4QT42zpWCYl03csKUlskuEVY
b9VmC5Y0epHt+PbSeo89+5wMDNVR7IQGlaeFBYchVdxPciySrPAKz1onFdxmfUagP/IqOF66FOIk
BiqC6BrDvkLXm+Qhq6mYC1Q+fMWlFIxx0QJKkt8qbq/OwVM+p4zMl6dL+BacjFmHB7lwzhx7xZB1
WiowULSTeEYy7PSLfzON5QvOw+ppECPnfzHXd+84mbR86my6coLUG3FGHutJ8Q2iEdwLr+r6w6lS
QnxEkrudxKabPFXAf6pue6c7JpQw60471K2AQzVEnAogDTuvDu13dM9dsuTuy+oSneKQ/kayenvA
C5UHy9/pSjcubiahS7DAOpPAwmtNum9ZRYLrhakJlzEJ0f3MttZ3INCVmi4f9/oCgOFKWyn0Yrfx
xR2sAwTW5cIfPgEGDbmZHo4uVufWbAuo45srD8h35mG6AToUUo1/Xq6dVgFz/AgPplw20VtsPki2
jvsmFt7GZeX5K9w6Ondcw2qE9pA71MdEAMqe1aKN0/AzitGlAsiz9RsRix38bcoEVPE0dLfGkwGM
jMkwL6MSCyx8FsabBSwry9eT2xD3jg646j1wDAwT4F/67myYH5TT95jWgiMjsxBqYVOZTe4AFkG7
WUhjjzgQjl/fucYEa8E+NkcBOyMPcovq6ZyELc8FPlsIDAgoMjJFqNWPv8jjTQw+/XeLc/0aC/9K
5EVBKVnQNuV816lfCP612JYuEVftzgKHbCg6WJoBCLVyaKgjNfAmmTdr3+Y0u61bV8inKDAtsAzs
ZaMZX2Q6++D0OJgOn/InoT2KqHWTzk4SRydCj4n+fUV67lhaHketOTtyZlox6AaBYiwP1i05S3x/
Kkb/iW71PKDk3K8DOhdSQ113Zw/w5n78iVgc5pks5SPc6gLDa2ypr624o97pRDS6/LUWqGHdNHWO
ZXMXE2OChG+xSfMjV+TQrz8609fiLadKSg+7Dj8Ecwx94YUMiroyuWWX22qqzma8Fo/ZkjSq2sq7
UxnMKeNfj0EKhzfyVyA8XT5GMXuS+7uOGW28L+N2cFwXcdOYIh8kOCKIeZu0a56CnJhhK4sEvV7m
LHzC301BWf48x2N8Abk02b8Ez8C9wYrAY+iwF4isqGN32KxH7zScXybrLI3wREyfaAgQN9TN7PIs
16N8PRjaEvPIvWWYGcENIurvHC+Xy5s+mv91j1ncwmjydzkm/JLPo7620vREk4LX/20Yzmt+l5RU
c/pl3h6pEkgiXbo818Gq5cfclzfclnPXtCGXBrozjr9QLBm2MEaSeDztQvog9ag6whEBggNXo5Kw
eZwPV3Xa7uY6NFD2eSV8m9/q5nt0YF65cECK4TB0/yP0Cd9R92uxxEZM805oaTp4qkyMV/kF+RD+
PK4I+wqYJyMfFZdEx29EOpwZ4FqoDxBSDdYizhEDbh8ZdfF3mq/VuXqVPSIpNLvjQLDuwkw67XNC
GkrOVayb1u0OtuyRzXel/laW7QFDf3hw+ZNNBP7p6dWZyQIBZsq7cM4ZeyZaXUXEp3aeatcDxvm9
smJCPoRDy5/oLqTKo+O0pAMTsmDA2AvxXdUT69LCAqqAjkRdJGtVLZT6DUeK+vd13NKJMt/Lj+9z
WtzmAJew7wihnU54nPy4+kl3hLd+4KRQvYqM7rKOE6fsClkU+qH+3OUZC35g4W4C7SxvEVLbwGdW
lr6WCSVUT7fJI1rkvV/FqTIGX/oWRj5bQtn/YjgScpIniT1G58xdKUkemAls194+3be9TinDxQFx
57x+JiU8RaxHDiltmT13+NLDWQk+hEKoDbNbEtSEHP8LSbLksGitiTZcM0Q3M5OFlDuGxkYK+Y5g
wAqzymQ1V0v/j8D/NbERVE/Rt83XyBTfIxFdv3967P0elVAaF+gfD0NaZnFhiyEzWzzVHfEpMVM6
+Yhq8Hv7r/edfAbA5/3sbIdYQNOwSCZJOjeFW7FcYg28+ylE9AmDgzozEHD6iqf4bGDS9i2GESVV
LMfesbHPbgGtmpXxZu8RQy7ptmdcfn0uhrFrX/mtvDtpU2tEOATrUEYpA05exdOGPVVCbxsXKEkL
uYswNTX5Ra5MnQ30HVJNIvn3Y0d5jTaRKdVMTH7iJo8/gFsdIkXFC5JNsp1IY6FQ5USbowCl5wrc
2FEtVJF8+QAKg2n/pVnuXdZ4BWNv90FaNTDHNAasfPWrv7NuTvUQjPJNztCyVhtBDdoGm6B11IxW
cn+KYZKo2hbqVIxVtK5z5iRPh8MUBCbJm9y4/Obuo4JljryuMmBa4xXAjub1t5xnnmn5G/uC+qGk
usnTvqSUdnR26WWuQ1yuaOgGD2rqBBS9E3Rx/9VpH0w0fv6ipgQOKZAyEe5m9+bsWYk2vSVcVR8o
qf5euKXfxSADODWLRFi+PFgaJ+DGOHcD1xMNFnWHksr6Ph9C/Z1bgpYeXGKuBKLbs7BnHZJqlSrZ
mR2WLn+pT/cU49O1NepTWuHUYimw7YHQn6ofxFICO+BYnGEJfImUYhsO+Ng01WFteBUcL/R3AocE
GFZpYfSPrb80WMG5pBFtpGLogNr6Zw8QJIkqXTmMx8MsO3V2uu85Pjn+2Bn9ORwn1KUrtlAKeixx
jp6dz8j9OyRD5suXtLW0KHktARMWxJFvih3pwTLOmICaAmJxMm3Kn2FSUeyOaTYBLzMbAC7a+wn8
sBxiCdGPrQUZaqf3fMKDC0WoybP1omVmWGQg2SKZIwg5sgzvnKfLQTAz1s15jVpmBsNP8K3nilm5
Snxg4a74JPrVjQwJd0aP22n+4KSjCIEStEYvG6zCZp4ItpftifPXmz/OmzoUPZhjJr31H7ztrlEV
70n5M5qpLIxw62Jpa8SJbTtH3C4sahVJFCjY65qDF4R2HSHdxRVd7B4aCb4+qqf5DqA7roePn0m2
RipsMHo+bQzBSjDmEe4fb+1d8knF5GSmm5rC/pzmalMukTN2c9x60F/jRVdEwkcw45VxOBfNs+qb
7IAiuRUUYdd3PSPHsQgygD8ddPokHAis5HUyF4OPiycQO67jgIW8QmUlwhQMQZOaIewhe0lqldF4
vd+y3QpVNbQtFyH5E8sfALVMbxNkgf3h4D9ZXjCSmvAVQ9z75breX73R4JaZX155P7FJKQgNhuKe
+Meqnq1Z4U4XBWvtxakaDinpwvmfVnBCEjh2gmlkZHplb6WI6Gx1tTedj5ziXiPpFYsRLFLiisLI
3uo4SXh0AZ9DoA2oxq82/kAt4IqcNzCeHzmWRUlJW03iajZ2TR8f0lRolZs0oUeT9YAp5swmKgMV
H6YPG36+1IRHqpyXh/OuAbkV2z5bGU2/v3TVToNPDkNHo+4i4Z/nzPTcvWkADAZB62OcSoof+d6w
MzEdBMioEW50oFM/6cS7xoC7ttVTTvHtASBGELPf8zA8Kg9ev7kzf/3Q/ThOxLXfB+YU4NFsbK1q
pRLgEsEo9djwxR/6TuJTwST+HqlZ0WlLSGB+AGjS8Q2PVaStFC4q2pL9QtECgCF4b7kGIP0yZckt
C/L3kjaerSuc6gPmgA9Exz0OnPmGRSVrwSk1tsXAXNyZyPdlEXA/7pezsqAly5md0wKXTQhsKS4G
u/C5LLEKLibaMWt2NEgR+zXDZmw5EgludFNUcbkxoFoKzt9g9xTQLztz5AKu9yVfIqA72J6AdqJX
sKIhzIvVyvHERdOs7YAFvfeBp2pPGd3og3z3uGjCn37x/r4cVAi3ReOvj3K9arojMadyk+SmeX1f
3xfbRpW3964gmwZzJDUZtv888rWWmmPnNu3dZLqOec14AuyUVDf7+oCze7z/08Eu9KYoyRp13xUt
hUozoCgM6qOdPTDHpHR+dOg9c1sJccKCYa4eiMqIrfrBfbCtPSfUG32SLO96puQTjVyiTSBEGwTh
ujNh91h0ywd1u5oiLG9bUKycRlWv+BGgPP3yGeE86QffX8PmL7dTVO+TNIXtoovTUc39mBogY7GE
/tBrcqCMPoG/rFwEMB+kU53FTMP8Ohd5eDpIZ2j+duKnc1/LguormtlohTvdadWCESErxQQ9QWfY
+ZfQevJMd5W1PWDGb1VwSu0LOa6tqSbpN6qqLTIjz0e+KjG/1wyjGla0qkGkWuI34prdBMHl/eOw
/psKHhpbzacppwogczWHiMlr1E4HVfjX4r6wGdEzQJFnpnjkXEEgyuvfUCtHLKbjVC9e/APBSPdn
XnP50/tNtaPSbUDuDzh82AdtivLi4FNOLC3h+jCwc8xmWaUaWVQ2btlm5DwiY02Sm4vBxvzIqrwo
F5ww08k7NdvlVmnUa/62zjGopHHS0WObO1ICI2OZiv+VopWkqhTuXjwvuj+Kmrblp+XZZFNmKmmu
BtLW96AIUycMcPSOcJxSBgjtXqqhD0eqZev0Xd2PpgwQvvMGvpsvqwU5sgZeEs6uirYp9U7ohM/Z
za7VOrsrUHSyZDDE98G1MywKSHcZ2mBmnx0keMKTXtEjio3ijj6uGOi4fsx5saFAQtMa6Dlehybx
lJ+CkIjqWNyTqNLEIn0Avd5k+huHg8+oA9n7GAWcT+6Bgh+UR7h9oUEqWPdSt3LCEofHKYapTgdd
3WbuJOFnlDSvJhTOkEOwqzq1hMQY6zuuYML2UsM+QBDd21i6Ta+LGJ7opRAibC5QP/s/ZM6DAImW
S1v6Xs4UHLu0Ud5X0Uhe69+bLPzgvphhERd52Nvg7lVNxkuj9UY7CT+O6+vHcZQsLf6iUneaDyZ2
gNyCzDkQreP5aoJeSis7AM3FvFH0eraiRPZp+UwtxNhZc+gJcwaq7tiMsxzpVTqBfruAEVnKhfhc
uFVhJrHHsXsoUiBKKNQ6dBqGZMQ2qqRq+YP68aNHukob7RdwAVRcS1PLltbYwPuJfJyQJdZzBqAK
UnyOzSTbH8hf4GOjD93Sk5fOs/ZguvYyDqZjIE4BJhw6naI/moIC+tJXpqBIb3+fJe+U6JBwEI7c
iBix8zJREYEUh4oK6c5kSX73MQM1f920gYUw8QzneVGiqJMGkGCZadwhdqpZPVETj1Fn0jJaDK01
YAUi0Ng5xqny3iIcwF9PUzNxXowiWtUGZf8nW/nO75wtAaYohrD9GTfA4l5nA0YRj/joVxtHcgeC
ifIaMim1Of6lpaMYghRnXYit+qAhJEjU6xc9Sqh7SScSHtkSQLgBkbabKTbcp+Xtlutq75DPtmKY
eFUer3V2eOZ4eI4Xqp/Qo+PmyEDyXv+7c+zLWmt+F/FIvkEu+2SBXEPJaAyWHmmOWIWb++ei+4qq
OoIRN1jEQMzcCk/luBZ0Y2OXjXoXCwgtKL6MG6IoeRbp42PPwmIuug3we5bf3Z9u7pjfYa7/26KX
Rlkw/eErx942HF9Ub7xMd2++JFKji0V0f0oC7oCE+L+uDCqGJ4Tl61Y68Y8ZErrzo5g6Oz6mLfOp
jnymeJK+Ibw/QZtzJmnaDtM+XZpWj4Ydic2wbZqQa69yErxBqqtik0/2/4/s7TRLNBG4K86H1thP
dC8mfnUApfUHWaApYgEDqaxqNEm5mQ2tbitNh5f3TThKq1T6xP4N4SgDYtJNa2Jl7QgupEWdP5Zh
ubt9HR3x93pbhGfE+SWnsdVToi+F/Whfg9hTNHogERlvg6bknwzN+SsFQjMcgvuaaXg9q6uD7YeY
GareI6rh4Ew/fq5URlOhstGLki/XwuzKJc7n4q37fEWE7ej/5Gq6wioTsLmMYBN4Gx9R/M7AVyH9
WMcverChEwS72yRCVesw68Ly0dEBoeyFDM5COdZpIr+NLgffMNvmVNnn5PsfySVLABmQo4pBEhpr
+jwQe7lvOWIE/OR2Sc+WqI6dvu5bV+BpjLC/Xo7ARdertPSskffx2sKzPF/7lH3KWTqOJ/RJNefF
2vWHZsUEsioZ4xEpeCs2ju9Ecarz5JdHvAqDqspVikzS+cDrhE7ELoYi657/vAENNXZQNAsyS+y0
Ge2Z+KCRbyYSl2WqKtlXxZKcrrC3DjgFJjaK3NpSyEbi/WHpx7MMxQVZj0AD5tNJlEjOrQ/4LN/D
3ujtcHPi7Jho2VF1SCrFZvwkCZRNCi6g2tI3iDu9i5VXs+vkGKJGUrmMFTtfdlyCUhijZF1I4nVw
hco1CFju73djvTHLSXUQm8M/sK+TE97T3YrZjtkm0nBAqgBGw79SX06WL+PL9Zg/OsrZufNITpYq
Jy42JuE4cxPpnz73RVEYYZ/d49/8Oi2SOx7gc1hQryuzo8iCyYwYAFrKYWp8CmQKMOjsMmu0SW+n
Pptm2epSf8kfiTbrIcFyhve4Il0w9bYZhxqXlSmRKlq8yiqpog6IxF+ImVU7+rduOcBx/wQmkggn
e1ONne1JGOLccSmbhk/iTYfWl3KuI1zYhfC+kOqMC2jLNmEuTeQAEoYhWEbRP6udyqccuhzWTM6y
6v4qdeX4xy1CkcyIUFaBo8MDa9l1BFhvbzev8C/Brd671F8Asdso5SXyXXA1FAklOqJiXb98i+Fb
QDbsqn0hSnR8cKF5W3h9TvebwQeWq8I7Licou7XblTLvm792PHNbqxa7REJnPil9zlmkK74E0mf3
jrqaK5WbfXYDQSklSaiu9Vg6GicJEmI4bs+SFNeKr/ObFcTsJjSucPqXAMUCerYxO+EXQTcTvT88
G0/wDJ+13EIlQ34PxXs3O4uJXlBghlihFxLmTdqdjfria58S7nSBTafhlUfXzOkExtLLVJ8QZrG/
4ka3WLvNcca1frpf9osmNBLJ3na+pkHY/Ha37qb14E4pc/OozQF2qyCbepX7lzH42ooxvxIE4Qfa
lyKWpxTOkTCf74PK7IUtvktowpaAGRgB7sAaGKJULGI3osuwkgA7/x2G71rbZYHeRTZxAVZHb2tg
XMXGthcVcVYYXeXXrJBwDGmn66EzxHQg5lTvzkmBKeZpRu9kARXGPoYBP23PXpyHvXQZoAsh3O1r
9jfuLrZB0Z2IuLuNJHLwJ2Bkqa8YtMJ0kN7+57sDFtzh/p1KsVMpect/SMdH+IsVCiqcssg1RxWE
JvP9pZf99STCw0vkw8n0FO6UPbsA7IsH4Xpz4LHgFGf1592rmndf1cSaJVcuCNSfH6ijup3CPlh4
UFhP4mDzmKk2R3ONora4khGTuGMb7oFmfl2gJ/OIcAF9dNFIIHJJcogsnl1P53efQEUMg5zg/206
bxlc0kYuO3Ft+wG67FgJZtQtU5hKfbYRFG3/UelaB4LUiXkGUq7qau3w/0fb77WbzQEPU7Um3bDc
GImBHgq8NT4QdKdR+CNw6cUHTWyWAYJb/cftCPfQ1Wqv/gVH5fDpSJDpDH/XmmA+U9Erz+187yQh
xlv6/ujzbd2Ii/mQ+FPUfkLsjwKu7JVg1huOKMbfpmohlauHIkiNfbnhAtPyQ/XCDLIRI2XvbVT/
W/l0awBz7XlWi6BrSgpshqw49LOvGaHkfeTXFQx/8ul65hSeVZMGDRQEBmbf9j3as+qr+8DHKH/m
xjNcNFPqJoLqJY3jE24oCbGr1SYQTHOVRExTcmGcDVwaidshuJRZBT07FdvFcMLP8Gfrxwq+Rdw7
kYlKYDvufgRTAHzx0ZeWQp2yFoMq2qgCi7Gj9Q5MBLQS7gp+is2OayMnxPwu8+FaK8HZNYAQ6UVi
EGEH0CbkEDpp4qNa63Bl/cx2voCm77w12OSzQNKQhCzswd3pe+bXRIwLrGYT87y0cwUxjlOQYYxt
mpPiGIJUw7NB6iUpxzmFP80QxIlOxBvQjhQ8trbP1qafyAkaGZOF6It2mkIVQ3JfASHYNiQ18S5L
gFzX4Ls1KURSN0izKgB+1wzETSVnwhlPZ/TKyt0w5kBhcbg4q9mty3hfQlldDbOffckYnlcFdJxi
/B2i341G3PFtY2f/0QGKaqG1dgPZ0DQ3/pvKonuVTRkcjYm8JMQmSex9RLHzPyqc+X9c67RrSACo
Ts+ltPm6JcMsk1D5DsflkX3WC+e9D3+NfbJ80j4370IQscKE2LI3qR0beDKENYMXQATb2WflAo9/
6cucPF4BxUN9jJxsmpFJS6isy1vWZwBktVHyhkpqdCTgcgClxhU6btcPGkYr+BLGpP4ncLuM8eFt
qss5BYUZd9WGovhPyNm95OtAOLSHz/qII27r9Hrpk+Jk5xxIVHrRt14JOHGpI/JO53Ul+hneSGeT
O0V1cIOEdq9StycVjzHt+SuMFy7gcR0Qp/X5PbtJNiL9njVSyHPH+S55hLSqWf6AV1ON8fUUIvMm
Chci83CTNXZ9FPnFGFCoqCtp+yBKXXRHBFQdl2gklDKAKlFUy97dqZ0zCAOw0N88An1e56ux0DvG
D85codC7m1Rg+CE160+A+bm3lV52V+f9YqKSqssVvV/UDn/o9XBhJSakrQvOSymZImmgj69z0GgL
1hLAc5vwpeLQKNG9Tn9/e7BlNUrihEQuWRJJC93kfkxlUq1ku/Isl2lTSyCu54rsjOKPqDsFS3XY
cDIes0MEeyo5rNLJ2FBCfo8PWVDzJmc97VM9RkIZxZxODvBFmNjWXA7vxpzyNsUgbQEhDqXsbLu7
E9Y07i7HAFDjthLuGnRDQO6fz6y7XqXg2Wl28TYXszKRj8AgHrhUeLRCGJbsUfkel5cGdoKT4EH7
8YxnbXzUxaa3Pnz8kYBngKvH3SnS34xhNW+Ew2f5M7n4G7UQb0jbF24W1zSXQ9d0vuFkV5sjw4zS
bYeZGinYQMpSAcPrp17QdVhjXOeK877Fuypufsk50d/NyfIH42cwLbLo0Uq+7ZowuGbbvxf7ToDs
kQRgOSWV6MItnOhbfqxL/DGCDGdkwDJs7Gw31i/VwjrvCxeENDZu/B0/TzLsw6ZghiONuBDsV/Gq
UtYaLNDhWzZ0ybEBKwQcqsBL9UFdr2fzf0A6ijFPGMPH/md/QdIW88LZJn5bsbSqJqW7NF/AqMee
0VwjIkRd5NUbzVgAaEiSebFA3BUMMcXjDVgtCBf66c+p0CZPTpBta5MJMbVvtl24HZk+Y/P2pDq7
GTk3a/p20fv2WO4pypj8W0/aPz9/jHrWvperhrU5whB70SnI8zXyL8o6/iBbD/urNYbqcnIRZrh0
0kz4VbXX9lwylhVQvb7pL41umpPMU9gnAeG66wdmuc3Xe7/7GQlNvgHcXdoUtyp872Hc1gygjJeN
llv2pCdVxr+zgCXujEi18jZ5Fe9C4lk2U9fyQOxmQOCont72WgAPujSKN3GPjSPsOmfEncgP4eIg
dRzp2RIZJpTnVOsP89m6uGHztFoqY2u4dpHqfHN/+BFNcK7BfBDPFjR4GJ3adR8r2moXc4+zPq0/
U7jD+5IrVVi77iEowpE9I7rjRSL8/PW8Kgn/MK3NiKUKAdT70nGiKLBWf0ZF9bvaZVuOievnnO9W
fRJkQTYrTw+s0ZVlq283rygXRJOgJm460q2UtPv8JIFGhBSeQeZUJQV0gBoRVH90TMT3wVPATb2b
jLCDfCdnh9Kbq+X4OFlxqnjSmtJI/bjgkAstGJq3dMTCClo6gfWHGQRiNxF/48fGQeTqQ7JLkT59
McX/+D2eFLy5k1z2i0FnmdqgnwD0/H9SiOCZHe/MZvQulfFYbCunicmmMW4vzxVkL5HbPV2fOHyo
1qirLgppE2j/LAHaOjNGYq73ciAPze7Se86cMCOX+lAw0+vhwBDsPx4y/NzYwdq3L5X66W/4q958
eUHoRsVT5H1wIpOSdqNp9n0d92LJwiQFVDC4HIhEz3Q3x30Wt0RhsCQgDBRPf18S7sTEJGjSbv2g
LHdlv8AjaYkDh/PdV2sFfMwZK2fdsL/2hVs4ae2DAgUs+UFcmiJlMESR2J+tWMNi2vQoHFWZxu57
oqHPgy+WloEw5XFQ8ZcaWy6aDFoOT3yt8jvkdj1DDVnSL/eK11wLb7EZ9jqYGDdAZFZ/Y97hlTtM
MRwosbP+RSo1P+weL+hSyeN5QuLn36BwObzzSTDkwbxuB92j6OUhAOSyThVt2kR/tfQ24F1qTX9E
W8Fw2E85JdzFx5W/r63s28eDI/5GW6M+hHHUBT9+aWNvy6FVOw5LFUPSYXLDeoqhpf1v0yW1B6t6
/x7o8Un+EqLKD3rLFd9uB9zWhDHUDJCBTBU0MWOWSTAtgKw640R6VnDgsxVl2mdiYR3Oa2L2J+3C
MtMtqs0iKe42C6+JJDqUvPsj6IfyzlXKpUU4hXPEbnwGONQsr50M5KCKwRQ9LNjN8ivfSRw46PUw
Z3qNdb/ssUDgEqPt+jFPBtqK7JiI3rSkozzwxrLG/04Ce38eMKfdZqkzlqGI+hzjh9LNf1KPUrXi
zJIyoM8m0K3ufOyTLicPyjUzCesC7rsZUUN2eihupoZhtqoVcSm1VzttCMlqpUa9gygELL7KKmpa
789KVdZmd6x1kaIjz3Iv+JM6QH9h4VqSUVRc9u/Z5jD+QdBL+Wk8ZydaPHBWhwG1+8t1dyCoZJrE
GNXfsQt0Nyd3LZStJcRPCwBGPGD6MsFygPfJC9AiLUeK+Gspsoy4yJ1hlZJeI5SBBlIy7HcSBbFt
hB2SZRHv/z6g+Fy9Nmdr45aNv7dWmbbALTPRPMhsCiPaFLQ5F9T6sb0W9c64EihPkemqimEEvQ/F
9NdLnalEWGtmdlny1ZYETXog8aHDYQIx8oqxY/LU9UyJoDwQmOpXXymaiJY5Pj/DhwaIKeKS3QGV
zoFesIRPUwnEv9YKIPXvUkmweMbq3YAimWfeSwnCd5yaw5+qOnTAiH6WRmKQ+T/kT8VJ6/G1O8sM
nbwP1xq/FEMAKSX+btlwozLe2zGoLw/JU6rF3hO3Ab9LfumQ34L8l9ibB71mD8E1Inu7iiaX6MVS
Rubesgzx7IRuB0xC1pz8G0oendRF+3D5yDRDURjywTH1Kz1SuPJMCUuYcbwDrESAuzNtriBbtfnP
cWd22bml49ptF/xbDCQFc9fpf7QKzp81/8GcKpYU5yTyCQCp1NDQYjo5p9urCyvVkZK5Ncx8z826
6Mv0P1ThCb0j7ak2/K1sknu37yFsGlQOIUjR3Jy1uSeCK3r8dt+TASL/JN6mve+YI932gYim5aRd
3ngokP97iRL+K+uAycFipxRI0ogaDnDUW0f0R2akF67lkxvAR+7Vs2miriE2cdh6By3EENHTJAeF
Et6Pvj6qlr0ynmLvR/uHMsKn0kx5rqUGgNhY5MNx6iZnOG42Ol4MY/mnSn3zblvJVFAz77oYugxt
UuMwkM6SExZxf5ah8Q0NwBB4TRc1XyglfULzdaf1+tHoF8Q/C7C47XAXh2jWg7YRdeIc2VjaH5BU
cPRlTw7V/yEeg0xTg2Cx9/K+ZmvWTCwTINZ+V+Kr/dkTAVRn+Ey2nSU7wz/GcKlK/ceRwktBEdRH
xWlVflEM82wFkuAni5SKjbb6eq2ulGM4yIgWDk0EQ9xv7RMEBHiBrToeJyGCg9WbzWKJVH008EI2
LiiZYa276BOA2+J3xqtUZ9g7swlrOBo2cOh8YWVb7QwFnOnfivP5lSpmwiTKCC7X6jvDRD92rg4a
5/w+vuDcDQ3h1bKBcBDYXbM3PICkSTFpE6uETAxCiBJhmG6zZEPFJDURKzVUKacP8DbLV/F6WTu5
u+uehH6mb7t34kgWo4+8tR0Ejc/QgfJiHeyHMU0je6pc5nhso1YqACqpwKccXAeINdMkzywXKZfE
0iSmqtkU7+s7IFWq8GYtNSf439I43WmIyf32be7LIpeVd8wMThisvFSdV3Dm7mbXPJdhA7K1W3R6
zp6J9JjbnLr17lA2/9FTzasIF+C1mq79ptqDAJheRUl1cATov7cH5AETKCLMjewi7YzTH6xgLtIu
F0/Mdh57BZ/vSp8YZjeL9OD+MNRGITQreHf2R1urzgEumnFiBaiMHhNBEQlLkkFKNwJsTeYKUXdp
gSfa1a6DtlPAnguDZ86S3o7L0BnefeIYeIVIUI3D7zl/vSNhjgQVi6MW9dJA+ODBep5gXnLprBMI
ya5mFihEUTINpBWgufg1e2YkEIKBUp15xOpn32mHkk1ATUlgGU7IXTXGXDKNFx6BlWZO+KrY3Oso
lRFq9nceBFNjcht4ARplWrY4uElV7uw6Wx66/DZ0ZbGWfvFoysC3nG6pmq5TR8R2TLdFFvgUKb8r
n29DTdlnnTL8raufholm0UW8K7Rsf5pKe5OtNN2PNBfev6ZpHoXG+E/u/Gwoo+48xpt2rI1xFrlL
VzppNaK72ZnFcHdI+rkp0KeFD/sYJ6wWSgAeMCEPAgYqzRK49K+HmGjgysuPasv+CNJxNYINfCkd
GHgvnVqyp9/Iinapn7QgrsvuUdfIpTmMPpUWV1gTSErMpdNojyaKPILzEXdsunkRpthtSV+bjNvU
gGr+vIoRGo8Uq+qdLwlqyoGIRMrVf3UCgOiY2TKv3/BWIhG9n0YruGhQCmD6l4bOl15Beqk+u5dT
6KnHK1dHZqPXhy7fJn/ytLxS3YYysKnfxqhHHiIwmQrh4edLWik8zSfo8UCJbIDx/onFti9B2ooh
M4r3u0r9tZQbuJ2VFLaEHDsjc57fs6GgSeaOZ3MHv8p8JD0+MsXyGwt42blOrg9OzjDTzSaw3a6V
mc7OfWM2UaE4b9i+44o7vUb60+gBt9Qdh+9Gde8zxKw+8BbEYHN5XN/0Qra0QQixCeqDj6aKuFu9
Yz4PBf2VSkIzXwcc+vEO/sQm1KAy3E/hiGkyg+/s1sBjinRTgPSdWfSTVlyo9x8uXecFV72H+W94
p2BkFDaQmqvDTsfqhuoo7Ern5gma9h2EXEyqmC+ecfXgjRrqA6qnIss0OazKVxq0PUOa8CbzNAqu
p4IYeS2VFnVpF1EYqty8vN4nKuQGIcIyt03x8OdIbB0wBz2aSfXV3CxFNktPh1llm3IkLtxjyTdK
KomXHa0H16xXowX9em5MCJE8TCI83fjeQhdTvFuBLP4bzN2h1D8sr/kKbZ1E+cQJofbzlCQ92eY8
HNQlqXquOJgdbvrK/Yh8rxSsnZsBRCoEajeMLZsJvfu6omZTTiX5p7eqOFvt+GY21wqWhNFOoHSM
hTo4fUTMlMCjsHvCDfDMxi7SSVsmG9YL3wy8059Xcf9hAyx/qGPf4w3ukqTkI8akAJGJ3dqvjSno
kBNWhzhDqTDsV68KGqi4quOG6fo9OwK2IcW4POjVhm7+FEvo1+UDT2OPc5FuA4tVQkS5eqh6+bqv
vlLl+uCAAi3N4pV/kyyDtBEm4tW0kAICuXoZvRjXACGvDcxD2y/3xr+yVYsD/Eh4n5YcrSlaowUF
uPSJLegu5N/fU5OcHLnf+y6xaiSaaazytt0wrTvJM1CUsqwdm/V+VOIeQ3bY/wy202SwPsS5kW3l
NgkzNWYIfKcVjLnk0HVVCJUN7Ep2vmWCSsEKrxaYy4OSx/rDIBEM3tLrpsXKER4V1dILPhwj1Tpz
nBtLNcji+JAkPNRZfXhaI1n+RC2PGhnlQjLTz/6yQp0i5G3026VziKudSM8TKGQAIOGm/4dyhhn0
DF1G7b9Tg1jzErNACDkrLU8OwAyu5J/qhDV+Mvv2yWJJQsmGrefQD+XqYJEkgtn7OfBmD+ysvwgS
ZpzNZKyo7XVx3yc9cKYsIsOhfSgi/Z8N2UV82lskrFWt258mY5SnV+WD9OI5OJOe594h5DTztKak
DmGDMZQSr8eq1TMIGbb5xFCvpH9RoD/p8cCvq/fBDtvGTNe+midgfuLW2jDys3Y+x9bSgWj3lSSk
K7hyoA6YjTopcuvnVacG4keiZ2kYE9FbViJ9zJlA7/AXx5lDzmo5bdz3a5mnYfYfEsU7P4276eE8
b8RPKDIM0gi+rWmYM6jHXU0Wscigh3v69ctrnIv83viRgRbC/xhiKbqStKGfqWARueVPf1ZZpRam
P7bWOHxA6fOpGWMqyblOQMBqwFyqe7H9ZYsUPsthKmSW/6L3jrooneSi1cXWhIySD6pxPqrF4pbT
U5VJwsI3wBQLBpEINWRx11XfgASCYK2zdcmB8aMYHLkjKzCNtyoMdvy9VaEjC4xego0QIlAksy72
OF1/s8/8ydyrmp3avptXACby7vXwk2lM+hmUj22UJXIypOC+uTkPh8/f/TfIM9Ibupav34S0uLUc
J9f1NjTuUJd+RSqeSjUDONJBB0REnMNlQCH2imxXy/E4ndicCcarx1hE4XVS+LhNUjhzJhZ1O6Yr
jZah+4Jokcj3h/vWG/aJtJO03W4VzPnBex6sH8xB8Q9qc/IP5vp/f6vJX9yjKPi59E47T+3RFEOm
GRZtM/CMbqQrUcv7apeFSraBMU52JLcyKEJn14o3ZXU8Ie6wOIuywwyurMCa6NSnKngD8kFti7gJ
ZY8iCIDKebnp42b64lHC7iwRUlsdZycu8Q5B30bPWdFwbrt9O5Kv5HQYI+WAzjJtzXt8lgEzkCs2
EUxzvl7K9jIw+GGkjVQUvwLrdGCeXJryEQzWJpgQKNbgilgmDOK/4GNTgoGfhSGonJcgO815CJsa
muWOKHcInXub49YpIAfZ5HL5a9ShAXUa/unhZ3sNjvmhP3EKpfoCUIfNWADNzPNe7s75GQrgNNl3
qpGDWWeywfqacNC94IcOlWOa6YTMNWJL/wmT1Ev9cNPxtbbf41uLH5UUNgt3mk/IHbI+90IPZi5Q
6jWLritZ8BUkc9cCTGZ+SihfebYdBcVWupQitBnVehQIqm+xjTSo9/oQ2YM46qz7AgqDCHLy3PXE
f6dMtuu+klPXSSpY5W7p/f1Z0Px2Z9gEyalqSinGM8pZsEkr8DDXfzqpQ/YTy6MKpILQhTuNlo0X
jsejO2x88ncQNQbAHaNbowhF0pZzxOvcbip6bWGyUS+Ke0bn8qa4ZYwpJdY1DzBbIfJCgJLWn4gc
d2iEdFDmlgf7hvVI3TAljZIemfYIjX2v6hNyUbQCajZ1oden70NnA4u57kgvRBxdi1cCh5iAYmWg
aAtsHKSj/S+z5leSl0/BSW0vKuSEKmPzm0U951L0MOPGqWNhsH4llv+Iu6xn8NPzD0f6SgScl/tB
VZiqD4k0Mw5yttQsZMurX+7LRYAhofkuB1D+dlwT4ibEQ39SAbmJS1uK+fUf46ZS5RuQStqukCPl
JYuIRTxvGAnEo8gGSr1CIqe+y3Eaww7IEpy6R88OkRBzW90Fk4bCBJupGrErRIDKE/3gaaCTj7cS
Bz9AfKBGTdA9eyGwjwIv9NhjlfLlQs6xUwzBz52p88WlQMmcxhoaW63MVRUYB6chdunYb37xpQcG
oFtVWF/Z6ZNfBhhGjAukRjMtfJ+OrtNaJ0htOxYiHL+5Jbl0Qzy+J1E+NQjI/jFvtBv3VcjPiAUQ
CiW+xk7RnScxgUlWy8Dniq6RZN7AdbG1/X1gIOaFEdX3TLMhN+jVANdG2Ngs24EPJaj3pTwwwDpW
4B80JPqtm8JA5nkjbzeBbSV0uPh2ZAzwWlx6rAyXJ1q4cO8mboOhLtE5VVJ8WNz8F6Ctyvq8KIGi
C3RUkdVHUlQsXu+4LcXjkyka04fmZgxjQy45UuUP40wFOEIbgymfkaHAN8RV1TJYXaFeQC+0Rpa2
qFstGHoDGLd2C6zw/pIwi0pTDaavJPl/jhkoR8H0jIOeBcFvaFQoZrl5jYAC0cD86UZOsX2L/YOK
4tozmpgL3jh0L+Nj9g/Bu6KQwJkkz+rS1IVykMUidQF1Kbiiq3V2lovGepH//Gr5l82YZKC3XRNe
UOEYgEKTEPiNtOQhmDNqhgObWkUUnSVC/qcPCqwA8QjHUOCbh3aHUESOXVrdDfae/Ch3uCN+AhKZ
NGVKFKEbS0oPOCwiCGtdeoP5kqCKuEvameMql+qOldU4iQZ10auXLBfpF8LkTclAjUcynR5it84/
+b6rsK5Zbmdokbw2hkcLZepLnE0F/SlTbrJv6Wp6aYOnsojZDef/yW9nFLi6J7HrNGR8alQYDTVe
MnEj5yQoEshVJ57C4mZ2vprOG86y5Q1CynIPmydYXvbmQPeaQZpKonfguRSUZs54f/MDPk3d9iLR
JH6rLzeQkBGxLAzpCe16jb4UF1DG0HTzrJUBKVzbETwEdSeLeYX6pyDWIjUrCLIaxRQN4s3mKfUn
z1L8i7QkOOEL1g3y5eh5vKMAjCh1G01+0JlFKLRKZJQaqum+79dY7ccp7tB2OunHOAg85D2cueM4
o2Qw0XmsriRe627JO5K5C1b8lfic0YH7yHq7Gd1PbShWvOw8n9fzSOPLmzHKmZFnFnFNVmhUVOgj
8qk26XlCfOQMeyQnWABT7IOqGOmsC8xQFpWGx1d07Tdtk2w/CAy1PjlxUoTWkNq7BA6NG80X5vJ4
ZB0dKgILl6WPrkAfQy7QHCgAMCv5Vi0Xs+F6rCpFovbMihMT2VDgxBjiyuRuVRNLefv4Qg0Jywel
IWyaC02MUuYseYJdbGamG4iLMHtnB3N+sgFYUHZIHnxZ/Vuvkmve5iSMoDl0dzYfoHT9u8kvwcL8
OKATmMoPlzU+el9BC6/2Z/vmuQJx14Q+3/OxekMcd7pzAfOKbY2MfvVjhTSfUgke3rcnQ634Y9M7
C5MvjT8uqPTdZg6/sn2cKS8zsl++zgSkftBN+CeDTxAFBnQBT9ELhX2NJzWr3OZ5VZk6hwnNh7be
ls90qaNqPBKotl64SirVERec7qTOze+sDaPwQ5Z5wn0diZ2KUuROCQSJovrizbdddaIv0OYxDlch
BcCdMbdhXbRdkTAk5mmmZUiXduHxRa8GIoSCxj5G7gPazDQ4FxXpaT9IZ/Kd4cA50LVdZpnMHsda
VArNmE8f489lXqez9c+e63mW+TpOM9PqONy4zH1ufjrj7uxdexrQWylyJ2TXq4efz5RJgmteUU8Y
LT18aXJFZc0vjXxxt8hpbiEHS0WmHoNQgGW89e57ACmIWsAi0tE6QljLHgMGAXQ+5YfzPsDr2n0K
+Sg7rQxeSylM77V/9W4GDMAgGJHf2kDw13PFxVKpHd0FjVX1VJOz2OJ24mz5H+SeF8iywMG7bDBb
VkRmMSU6HPXKTZcZDyA9K9TcHpMMTMT5SXU3RxH261M9hXfg15xCNmUfE+VTaqBH7caX9RtcBLiw
zTRRxe1rvpWt1MteR4bZ2SO5fhNYCl+jGMqMA5VOWI2dom7HSgU9qpAO6lEhEvk74NhQL8CaVZwp
j4wGcdc8PSbhs1tDyH/4ig7n0l0oGEZksjsxsPGDV2gKvJRG4tIx2TZ0g4egniFRblocTWgX3PMr
6o/ZM0h+eoC7E4T+EnY/33UQqEg0YBHHZj2mvxpBSaINuPjCZ4LLVEhtNA8NXH1lFYdH8gM68nYm
SjojhXOYanWdwenOz8ZKIpePeYBeKOiVAH+CfAOS9ygSqNpw+uZG8DkZJrESXZJQsMh/5yXWxVHr
VCpRkgqdCsHVey34H7SMagO7K2Bnxs80S4gWpwG8L/g3epSh1LlyErNtqJLTWXEIRHymwypZvWz7
SyJVmxU4jNiodY8NxdkozzU2AOiRvHx8fQbF4Q4udbTNQMIW4/cZW/TsxnBCwZTvJGUQllR+DCC0
A5zqhx4XSefSZJrYLPh8e23gh3vKdb+OWFoTjr4QdsA1QZEM3nA3eURCoywA3d5uSB+iimc/tY6V
9eXNGCqziUSsT2Ecua+6HEZmrG4qv+UPgFW/JcTyZVnMBJe27Ig0At3eJalBvcGo1l3tcQloOhUM
BZ+5omR9YKtCm2hjD4yAan1jd3WIDc2W0/TZvrwPO5WYIW4X3itYZZY0tGMAm5i5jJrQue9UJsKJ
IID8PYuXDzA1/rUG6f4QFtJfOslCtAFQZridcH/fb9UtobY461EOtU5sugtysykvTcE5+1NGoZ2e
gZMOzWTTRZ+1KHWVcwXsZyzqAz3QCe5kt+l6nf2Aehw7yd1ncG864SO/b2usMRpUI3fCAyJuBXG8
k1kttl0zdF7tLhz41s0TIh1Qdsd+L6jcWAuSX1iq2mra5zEi5ZkOB85YZemdsRDZx08QcgirDXGm
t+O6lwBI2AjUUWxHGmZ4mJYPE8vVg/0xOgInxoUKOJ+hk61wB9rslqIjRrhzkJ762VjhBEJDb2sp
SgwuGUF8QpHKqlforpjFUjyzAj7JpcpDLiIFX8xyu/S9Oi4dMtIDi6UHI9qQ2ilAnudLymodzhAa
wk7H5Dn3QcFzXm+0Yn+MNHWUuvVKtTCS4g1HCpbO69PSEI8zhGoQwQgvbgdkno/tpRI8/4AI9dKP
6TWVqbFfTu+Hrgs6+TFJOzIvCh1I0Heef3OCLiX0MUnAY72MY0nnuqJ8DJUkLAHN0dKR8JbordHI
HvLP0+HJZiJwqHZ6eZrcqnxgk6SxM4nEvOJYa8pmZrHqAjl0nBByHGgAqEuCfFaPPt+MBOViPUna
bCv2GplDPPTaENBNuAdG6deV6AdJl0eDiGDDBNHmQL8CPWGJY8aEUCpBcFavO28Igpaap7oKMgKp
jTmSDFF8QEkmZyXpIUBfnIMzvLC4koZ5ABJ8sQu0EX2BALlG8ZeSchthHYu7MLcikKuUAD2tCq2j
bnXROSBZ+WOeY+4MI35YUa+Qr62ClWQcxnOoXuS66F2AqMw8V/rztUWtJmxHbSNqCPEI6eyuKeoI
K1/e5kARpyMTgXXzw6i3eqohOMQwJ45Cf4NZRbE3XMmbzY5fN7R/w/VlXhvHp8JAn+yh2MxXjWid
avgG066UChv4dv9uYpPtoePHisB4Jsk0wJLnKvZ+pusRp5dXlruryiRIqVkho/DIAWdtBeFrrHSN
ut1dvPqVsNwjp6m62nMfDtymCE1CV6xvO3LcRf+hu/le+X88TIoVE1ENUFqFyufDYH72pSlVL1t3
AHa880RYdEsSC9z/iz9T7xipz5jRLNSjGN/8lf7FpdrvRv6g3Z0DBWrZb7xVZfNucCxel4SbowUg
EjP8B17g422sF3OVlV/W3BPcwTHry4LARZ+ZbuiAoPT65tMIUO6RRDamnjQmvNtWu/mvlogy3HS5
L0Sscw33b+V99bB4WFScX/0AYiAH+hZi55iO4eUZd29pV/f5I9kxtB8/yPuZoo5fyhJ3Yin7/HSv
/TQsUgYbFefrweG6v+eUqMf0rH6BvcIBiEcLCa3LO4DKvz6w6FndYcrms8dsEhvEJC9QWUvAiq0M
4NitssLnhhO4/T3/1Pp1mF/3yLSfjVq6QVcwSH9yA/vu3hUvoeMpPN2HcIbMrbRmp0O5SAIUBROF
nvX+A450GXTpMv480hPsTrzfBRscdpXLtpq4+i8lSPXQMDVlZQ4I2ErtGlc0AqgH+gii4wN5WFZx
ybPtCxHS355AfXd9Wzr8k1tT3I7BvoV2gv5NLRSFC8x2iygz7+c06xx9s/Uu98zFIxYoc0C3ZfJ9
3q9m/RaCxDwloYFCJpo+R4+nHvjvD5yjaMGiee8jV/0JKg3wu0b6kWfoCii2G2T45TVXgJQwzPxW
BUp4KINcvrJmKG1G6f9mqF+847pvZQ5Cd7h5k2zPBipGuYPNylXlZ2aI1YPqpdqn50qgSXtwrRwq
3jDuJFG8sFnBk5WBoyUXd3P9HxGyeuPIhcS1IlANp1qtQW7Y9jyZzU/xVON15onfHKMtdGkWB7fg
5ZQCEBDeHNekdlrtpfdW3BwLkLb8KRABUxNs1nKQX4bYNE5U+d4jj/82iP9wR7vBT7qyBMvYXZFR
g+ELNGZlwBAZNTuOav+bcUaNXS18xRKbFPnjb5u760pyNaZyWFempxqZm9/eU4c7LuH4bliBQA0o
JG+lRzuXav6LtxOE07gRf+KYcYIHX0M+chR5YKHBbmPQrLTsKONtCq7fO+C9JJr8BvoK6AQBMUxN
V46WOCmQMVP3vad5GhBBcH2uY1gDvlnqa2vRUhEnW/rw8pG5jYmApOhJPzmhOx9jDF51FNq2wbtz
S7IBt6f6ApM/nNjc7F0XTGeRCbqW71WGWh45owBpNgWJG87Ts9kdTriN+0oZ1rSWZM+M7pLxAbVy
dJWfqgCvPySa5d/RKEKd7Tm3qDUJdGZQPcG4enexuC8kBBzqK+kosi/aS+PEfIz5CWVoS5I9MNCt
rfRm1V9w/7+8I4Wo2gAgoAXHPwWRd35Nf8Lh4Pt6h2SaVvaAcvygj1zq5OJ+UwuGMNHWQudhRk8c
8xWAgppR96kM9mprXn7qyqhijPeKlyaC66A7k/cd1rbOkO7ILObRjALVNwuFcarZtFBXnCNfMxG9
+seBiql5lWm5rgbM8JPSJMdx6zl/aLJDY3k1S/88ZHMTVIv7+tAydOo0P0tGTC6sLEtxPrhu+7Ax
8AlYiC4/R/JTE3Ovn+q+/IABwXi1aTW1yB9nlc2JINcR2jGtjhQTDLdDDno+3yiSI37EFpF0NwP+
cEdoNB3K6y7ClqoDoK7sUtHlyGpSF0St/z6qI+v1MKzkWyTNBB9Q2dhfAerHNUTVW6I/oUIk3QD2
YZ/iWGxXU/SOm1Kud7d8cpHzrd3Voz7E5F+siajFh9D88OrJFA1k9gR0N1TX3KGGaAvUK4s1o5HX
hfxpQkQBplW6MKBiWLrQ2WKZHcHgmqwj/gGdcyKhBPcsbUzCXKn/3GATpJQAa3pAEXggU2DwkbDG
GAlWbSGKR/s39niyZSCr+ydQnJOwkNU5ELlVTFQMapaFqjzS2qddOGY6afPVHS70YmcLo5zUWNHw
02PWRnjN3QjiRpkmlySEwIbbP3pdWb4Anud7kdqiIJapKZgXfjMP0DXWmgCdxxAWJUDfhfS6O+Ef
ezq9QrOLNRqG2mG1HoFiZSfFXkLZPA4qYnfdKiYYl/nuY9s8nPyP1u4fCkjX/bI+mUoW1jtbcuF1
ID4BbhfaT737T7OMqLMvNrtN1HzGqFVrcEMLspLKmWmr4qI9sFULZqs5xmJbG1/VCABdinLOv2r/
Ratmz0JEVk8kGNchakCyVfMYlde5JvSF4dT59u2HxpRAopJpfNeG8Xom5x9jgklq75TMCNweAFyx
z8EgfmMul2/kPqg5UxPUtRkvQ1pj/UDQ4R9bkZ2De0E6+QcuUlZASTyEkqoeNV+OI0RMaitKVLQn
5Z6nCj9SsM/SfKfhZ1Fi8R0A5zs6mGi4lcuDmkNZWN2aQM13lUMRu+z3bFTEx/x66adKsnwmREko
zhoB4+NCZToKdD7E3geq9hcmW1IGZkVbKlu0RVP50+jPtqhsd3XTDmFzQwtkicFq97V1xJY6MKBD
A/3/RO3LS5jiaPzFjiKG3lI5KwlPwPmtEZoY0L1vERwqfYUwyOWGmEDv7qbcQ+1d+ONVywhDok3Z
UALKwtkrcFdY+xb286U594HVbvHHO3Os4oJCGtOdINKMKvDXzS5GoQtS9PzpjTuZBlulNr1dXaHA
+FZ8ujHHaJp4J5ckV/R8/9x56meKx8Re1f+dT0KaQYcc0czF/zV45ngT1Q6a8tgfOvm8O1nUAmjA
oap4odQfNIV3Q1Bdn1eVUv7lLQlIFX8wXj6bxcXF+PNxjnKCeof0YXanLwZJAs4zyOpKQdrjo5Id
OuHZ5VPPut5KH5cWJ7QnbU0nuoLzSbAfqliZsF6RAE0d67wMuL+kiq2CQcDwVX/7TETBpHKVL1ub
pPvw2wqoXOvwVi2w/vuHpogYekpJmzg6MsNBJVm5AdjwSB5ZO6daMlOlkuKLgfR3/9mzKQhqHh19
JzG440ZlyKeCOEPQiB117GBNMH86qwq3UebSJcqHnZDE1rxOsGHLhGoPH6HsCAl7ABRF+c9O424k
TMLFaF27rU6MQM+oLsjoQrnfG2Y1XDXMPC15OpCPB7tTILpmYwJtpjesU58QHsCnoLyWWZyxh3BB
zTPvNGfFYE6wof9uUL9JXihbc2bcA8gi+tELeYV09Y58IxD/tLlQQiAIVwPOTvT8ed2t2gbVZd4j
x4bqLYOW9GX1uPSamGTwr4XAvZMOmrvPICtWLUwLUTH+Kdlz2QNAYCiX6EjhS+hMKPxt4tq2Xjcz
2BK4Q46YgC/Rk5ADS0B0nSqp5twSwEV4O5uh98o9O166DunWqsdxLQoYPhTp6osBZuW6Hchh1IDI
chA4cf3sttP1sUZK/k0HPbhOvJitknuW6nBmNCSh7rx5DUAD1hfnPOy0APnN9kusDfgPDJe/sAeC
RjQYOyllE4ySEv2W9L54NnNunMFYAKtYiPvhG5nXwgXe0inIEE2PJ9s+CneLgX0ac21sCHtLO8i5
whySnQSXblO2RFfaOaEiWjQ354x2Vxlh70nSbeCZXxjGkRMP04bzn1Xq9u38GL0MUzmjQiNOCfGV
Zs/iOYugrwMDGTpJu1DMY0hC3Nw0Oc4Z2TIg6VhrkqTUryVVASniE988WULAUgp8jwN7h+i/mHCx
x9FtGX2dg6K3UzI4l2Azl32itFIFqY5bHAHe3wTdRW1c/GpMRxtn1P5RZMh6mQVUkoDXRYco66g1
jiQoapoHd4HF3J2rUB3y+Rp+ipTOyfSs6ZefCkjqfPCHpKcvHqaGH3As2e5mk+TjE0iR+sW1b/2M
mgMrk6V3JD8cuuSYl6nnk/1rbYcpW0l4hi8K6zTgFCqoJCZLyKgN+RRHi6RsZPx7ZHBH4BkC615M
xckPBDdVFc6ZRSDpLymto8otoS7bdCG29fymB1YfDdwLMrWRLZy8L1FqnZ6b22MZfZcJOEwIe2vE
vLaiOv6uV5J1z5Sul2M1WRKeUXxV+lM3xfzeOj1w56aX+biC7TBHcIqcoZmBpJwsNAMEm6kVIwdA
/RWuLnLNUJMj+k1jwDKaCxFxVYlYWIgg6kh4J1SjoDlvzVjlCzyzAqGtyAonYEupKvy8RqNP8vVd
aOp5cEgYe/bsRdWsp5GBmtYL22PByASgj0B8SaYOTWgMpaGlGPFyFvi9Ei+yw6Bz+ftVe4WGtbv6
lTuCdczMm3AvYHGBn/9AOvCUY0jyQ8J6WYM9H+d3zmg6+iAVxTGrg/mbH+9/eLWYjASb0CnRKSlO
VuVarjU75aVxAB85vlY2DtxpimenYTirWZgFJcjzbJvQOgbrL7DxtWcEJFlq0LYBWR+eMcSMbEo8
Kz7xinRwLKUKW/ruTI7uBaItsdrjfd+uU0si8ILSbQ1FPtxnI6FMcKcg2pksdcnuCusmJmEdZbO+
B3AOcnpqZvCZQXYHlEJEIf9mWHaKQARgG9f+NXpaZR0SnzYVLOgz8GRRxcrqKxafHuPIhByfCBL0
0elHUh0vnSVVrhJ8rDDVaQT7hENGn1gHK6Jz1YHLcPMtJuN7CUigbqsH6tTtcXqJlmTT7A8+mEG6
3i53hHJM69VvhMHA8mh1A/cjv8W/NUa6lggUBhr4IYpb3DlPpeTXcEi994+M/LfU6Aat8NBqTUdl
TM/BmtImT67McEdBBzhaUizceIBPePiHUN5t8cLyMv74h2kFqWeLgPASjae+Qifb65D5kASte0Q6
JZdZ/R0tidOhaErRfNsriMT3QpcEfLvufT7IhqOy/N7Z5IC2E2CS0vEzPi+ZLEWcC+n671wUTx8n
0Vv8rB8MtneXm33RJMhpx7Izg5vgZ+vnP5o8GQ2CiumUcgEK3E7tGQs/WrOCeL/C09glQQR26sjz
IIaEHe/AaNKmOWsJjxJK99vR0aTX3cHU/H9ehAis8VoDUoJ4mXwe9u1Cj30o+eCxSb2tapnaUkak
VBuYN8TYYveR3TSTQ6VP1hQkWkK4+gFiCYLoq6REKoyxscDO3owU3FQ1aHdynTbIoMzZ/4Zqki40
fuRp3DNVZBKG3/kTNdSg6CkL+OIO02xpAQ8v7GfVgK1WMGVyrpW9e+V/qGzw4eT+IHn1bvKHnY93
MbydUUqzhsUPcKVAt6QTwZ8SXl/g+tptmrk1i0sbiXFEMPKTkQq+vm1wZg6NoHyrDEVHQirkmew3
/tKcDWz8m1pKsZFxfNjLqCg3dXwaEaQ1kcV30qpQlmsQ9ZvN99pfpullIr+ROa6xuUUsMibOQNqc
DbwC7DMTYmrXWpuMmrNYGGIVoChqigyk8rIO0MoJTsdc/ZJSjnpsX2K4IfMRLOaiu7TQnG9kWekg
6Khtu3qCDRhw8mFJJDngf9zquKbz+hJXbVR1gG2xIuWnnp47iRLi0mKv89lF6ufg9ADd+7lWCWj5
AFc33VFqNevBzt5+NSRY9ffXdTwbTcflD4TCTvW0eiM4MwHcD1P8fU/V7GMAu7XEbHLH0b8VIvP0
frimjhPOtXt6JnEzapzll4cDMzvCxm0YUBlwKxgC5QTMwnv4M9Qt/NmX+dHnnzp5dujHfDUvn2M0
BTXdjtNgooftawhSlsBB5DUwCogA+CTtVgc+E9qdr6uaN7az9mlaJ6tn/Jqc51ChPhNZIlfv32rT
f3Ncs4c292JF+cajWbxlw03zmkyz0SsUB2X/Vwub746ames+K4hC9mg7I5KEy5TyHnX9ZJE5+cT4
hcyJGqAix5NnGFSeqx2vbIP668e6ety66mvFG8QHGkCOQcqbUNWgMzUfEA1uSPtUaVJLNS9AgXwQ
LALKetFSP6yYNKp8ydRePxmhdPQQjYrYX1izUlaOTtwW1BzLNxyAVawZ3cqWvQPpflJCYrDV4fNd
aYGSKGIUNknweRELOJbUiYiCbZo2b12zjDq4MY85RVpeWGArp0uLzMUYuyUW6KWiVTP2aauRERNz
avoUE7Wzx7F5o1soG72skWaLQdijHykwbGr++tBYC8oeiVZKR/JsctoCyTUQ3E8r4/eiVdFaDuxs
hqzZf/aIVN+PAGwrJHhZom4s37U0vg1Y1MdGAeHLuLUMk7lPHwE9GGr88rH0I6gaHHEWbDHL4iCx
s1ALg68sVkuxl0V0vnHCgpH2FfJOzNPPl7g/KEqX8gP3cZLBUEkJT7gRjsAgXhEEEkNlPRJ+9GVE
PniysEHxRM/LZ6CIiVCQpx8qFrUPDZpa4ahdW4mEGgX0zV959l4pQs+zYucPy3RtNlkVp1kcAZmy
yuMfUiSManf5tes/IqAiB7nFYjzl0DfDu1ALkGQ4dwYlk1b16+dAYwxj0uxYX8Mi9QWDRaWltL3a
v98CZA0hB16JX7wP9Qr/K4SFPx83VPES0da1W9X1Mo16+SCxGfC6UkayUk2BGRK3zrewuXqKJEJ5
COG+xXt1YI/YvquhGxqy8dMMWUTbmXUaP9QDBYA9h5NSGgHUWHXCJWKR4bbnlREe0j/lyrSkwLcw
oofsFoZnWap0atzRdnssF8a0WNkFvjbDxhEj7qFRkYsLQ+Tul0RYymwXbh/gMgZZ3/y1IDn+bpV6
GASinoqYjAawI7Rd/Q9Q1XggfYTlicH6HX8NEgnbTI+vM7Kqtcs0jLZ49KGZhbpmPmrHD1wwYyE4
itlU3nHQtmDRHFB074JI00j0wcxEGVbVZSZD6CFM3i379/vpxrXYpGkWYwVj9DT/8rUTFNGm6Eu6
+qWpHQvgquRHOlDssONGWT/CsKhn4TKYbzBVge/6gYGBOPqSYn8kM1eetNhH5QDyfgGOAakjzJf2
LqFHLJAsau70j5tAQmEwoL4B2ZqEAmq72kuFW8P265PRvvPD6qS/z1u//xbydrMtcTS2evBsKSmi
nSq5oOP/qKGTTfHbPWqcnJRDwWpxUFwaieSppLDvra1rCH8NLeuofcCQU6Mdv4an3lSaMjjj+eOR
Dw0Eonn2/S5HnWUFf5wstDlbauV0nM06Za1CLIE3zlqHii2YyDxL/t+QWWTgp2sWCK0OFdITzkok
jd9tdIL7L6bNQGAiV0qiZ55b1IZYwDme6vbqywye5/801Xx2p41SmbsBU8DK+cfrwY+R86g5BnVd
zSC8yBn5fJr/POyHslO2MpzoyTdnunbTnYOGBgrepa/r6fprKzc12Bv5Pq64+P++m+YGfAAbNlDX
ySZH9h1cYwKyDpCSZYg+upTyrT0BreOR/p/9OAopo2NkgUZZe9L1/zNeci3iQWU1VLD2suPJtXMS
cPO4e7Iddv1KpVP+Q0NKPzOfQ5J8f0DjoQSXIBmztiOFy8C7p4okL0n6V4sf9QlVbC6cV7EOYMsu
vsf07+R/5IwbcPKVSxD1N5pHVhPqMBfL7Yx+Oklv4+tt5TydLKA7LWcDxDtRBQr9SFURI3pckCIJ
9SVRgcUQJyZ4xXqa5sMJa130l8sofpLfiX39PmjYYh0P/fT0bZ/AWhk//xjT58j06Jc4sRuMFTM+
60jfj0zGiTjByQ3LQ5Dy6BrOzgZg9hOPQsI+M2u2R2Lx2L6hU0gcKww/hCRAz/N/3SXf6mmWD+L0
4r81n5NWZAer/RMsmIAz9KpN9FHt64cFIjlJ8h6QaXk/dIuLrFnVH7/y3R4ZlZZSdOGY4dCnb9/U
uSsmAzyinxSGuTL0CQHVqFnJETuMEj1Tha8Me7zc/e9b4kpP60gl+htTpQm5Z5oDX4T0DSQnzF4N
FD1s7ESVNpXpDZIFvA7IGWTsPTtVHVEjsW+KTuFxLtN640L379rDQ8h7IxgzqDB3Kvaw26YAq5cD
Blt2YQ6YQ/KPcuJLCK7dl6eRBZVGUDR7CRVEUTUJy5WAVdeLWyThsPo1IC0MMysdoBmi9GV2E3Lb
EPtfMzIwf+a+vEHgpsrrNdfwIKpPrgNuhY44xmCs2vzW0C8oMFklJTNKW4/1fFn6Lxoiozr6UKHy
bBnjIo9JuRZ7zj+Cv+QCiO0osxJcHZfjlkCD/tm5jg+JNm38yYKGxaY/8kl0kgrErb54MB3AzAH6
EnfoGGDLMB6sk8bM9p+xwUVMg0dx2Ah6IEMGlP3zaJBeHbDEdgV1y3Ftik6Zs5q1eVbO8jElTFr5
4ROrekcvAxVn5ZRKXQtvd5YVty46rQgA+yufQV4HM4AZdxSDotaKqr4Y4HqqhK+AEdjKEhgQ0a3Q
f7qfW9dn4G7m/w4ZZwYiW00qwsxX12xKzu7NQJzK/DfrgXME1UMEhrvF5MqpFRHLXb4YwU6bVLzP
bHGWYd8fDQ9TTjcrxMIYvHDFFoU314oPpCa/gNaGRiRfiZPdyQsjDIEB9ShrSPLj0/swvlGQGFH5
Bg3Q94ZV3YvCGr8XGkxCNntX/I+UnU3jFMPZIDNc8yMiT+xQl2fZy1kPB9UCDd7cVCUHCFTcWI5l
+/prdcHLNJe55p//XbA5dndcoDdKUQdlb6gPugJlrB41O0NalSkkcAQ4kiwY+FC4mZ/XUzaUHeL4
QNDHLHB2huf4W46PPCIDQbjHFLvsk2vB8hYlRdiblrnRQqrmMTQzhbJLCGgCsQCYnY+T/XjN5Erb
QuUB+j60giQ9keQ26LnSb2RCLxBiIQlWzlc3y92um6qvqYxPfWbJNiHB7SpN1T1BN6o+yWfWKH2c
exMa3AHJELIzXYriIr2f92X+RoJwL/uAwIByIakZQNiQMGh6y0rAzwCeyWqm847zZ+luxn4+NMo2
wKwCgvDe9enfFAAmnlt+OKxTFwXor/oVsydB1QV874IcFsvNhZuIn+76UzwRYUxG1FXNopMdO8HC
24q22BAoJB32q+yt2SuQJbKQuB5JUgYKybpVJOiM3CXTv67/Jz+TvtNaJVVQp89NNW9AsI0j2Mor
MQAEVVGLAUl7DwpW+37YVFFwosDwCgXWxold6NJMyzaYKLmu3G0ITKVaYqzDc6BejlOrM1hed++e
Jg5Fzb3hJEc+QSyZ/5/Y7JSXJq1Jq2DvS7BWtycuYym095Uh8ZGyn6TYhdih84KnTrLn+CXrIPy0
5jTLWczvGhR4gJ7dgkNLnAfg6JFKoEY+4Xd7+WtGzCKiyLUPgvLSgG1t0P01RM2nJiUOouxQA/SV
Jd4ULNV3tb8Na7N8LLawhd199yCtfhGb0q6phe7S+ichOWHKdmvwhcrpi3fgE/z7VgwQBwY3c+fM
LK2vO1ZVDKHmF5AnU0gLFI2U8X2KrJPbJ+nOH9WKNKctQl09TCgoZneff1JvTlsLOBZ6t8cefW7K
ccxBagWqDhhCMw8LgqmIJAgkKLBVO9g76wDxzjhwGHOV94qJ+CRM1It/+/YpPAkoVi475mZUvB6i
j4uUpkpAsUFSCZVNK1UWQSFiI/A8R8fl6VBqne6euzN5LqarNmeTmxMHMMbVqsTcrYzJUhHd57lG
h2PoEjBoFOcOfpohKuRibpb4BtL+aoBw4A19jwY0wIq+bgh36Q6x+fr06Ao8pXYkT9wcM1Va75OX
xwc6vA3ySATx9rEKUfEEB+hkfoTy2nm6GIX9C3VXo1g/um8CSbczlB6EHvKxQBQQooH6V/WjuiK/
QPXxQ/dKlZcKWmhaY3DEszgcr7LkEFEN/j6jp3HhDp4r8o83auo4NSg85mVwhMehza3SAdd1PAfq
bVe2Vk39thQi9qgz3I194/PD8J1GBh21sZAASvXLc5NMxfdwp+wk+C2qDoKW+FALcNEDtNguPWUg
w1D3kyKwCbrkij6oRxyLo5qIR+UEIicFc5RJO0df9FQsOn/cDWnkHauRnAeZnbfjQpKpge0T8yh4
IV/hdG7reog/t9bol5vjDH8FxbJWTqQGd6ENsE2opzaTJVOhB9Tc0XVWBXOGTKp0kiItVZHyDhU3
ql5azDGZThAXwnafSscwPPOVj1G06c6L4PrjvV7JHDvsylDVJEkOjl6an80v1AIlj9WOL5HYB+3t
hfSTnm02fC0iq2DtS8RcC7Cdpeyee6eeqNt/sY2jKFOTJUY9wHDV1yxSehepfAcbVUgq0FmgDlne
L4Do7lML3MfaddUjNvmlU1p71Q0bS+ONpI1ETvN9pzoXUTCSDJ3CWfQeOhjOx+W+OGE1NHLhBaof
sgz0aLc7nuSJDjcMD/5O3f7ufvzlSUAiXVEkBEzfdYU9jQL3pSp0uX8Dlho1OKazrivBfI3unBWz
C4fw/XXnuvJFcAEVERaHepn4ptAvhkDMPVJhbQFTFFLixV+olBnBwlPeti4/vrwv5mmb+60cEk9y
yGu1qqZp/xbHAz6Pjovei6r9sAuAgpTFAU2o33apMdtsTvAjYgqeqFg09vug7BeKYMXarbtQHM9K
PCwA7gCNuaigTXhqvvK6BBdNeh3p0r3cceSdjWNLGfcRffP+J1qRCsX3QiNiz+1IHjIBdk9byEEg
MM8/7imga4rx/Gm6ff7aHRKt0L/TQUoutlZlMapIbxd8v6ceDBk25hUO6m/3XhXSkHoiHHW47OgP
DPGNSUL98GQa7i8oC37wtJRIuEeIOOjYghy/PTJXc1bpVeOLrSb4lRsJLkULEsnZDJcrK+EVuGtU
tep3s5i8YW+QNOrCG8p8XRFT7YqUANui56a3uFZsnZ9raCmvXy2pUDCQyJC/OEVhwSbgLbfRFtht
vQUTA+fGVv3O1esUwxe0K2x9g+RuFGXdHjRk35cHzLO+rkg7wlRykp1GFitZ5zuIcM/Q3mQ7+eIC
b78jRueqwe3TEgv1SbXluqhx2stp2YNBo6fTqXrAMudMhYLbYF9t4kGpZPR9ZFsDJGtgqEZbA3dq
/alSpF09QiSGIjs7dD48XOTUbMMHFbr3dImnREI6ItnfYNMHqknj4valq1pHa30t00irN4fBXHCf
8xS/3kt85CL9PXBJqAshA21CBtGUMWX3xuY7+pJjyrIAui+I61ZN6cLnUEMSGPVkL7eXcAymn1nN
wxDj/btqrjq66LwUUue14nuhc1I3DWV0JLa5nmeztQ4a4axd54j+Jh6JW0mK2p2/Ya6zbdsyNKAR
dhvZMA+R5tJjI0tWnw3mBql8mnJ2kT2gHsphPZ1B/srda0HEEH6ZN9Y/wxoc+r+IgA0rT/EJGAmU
7YTpU9GxlH0wQoB5YXAvEKhA5SzmjMiNBOkMjy6u+G26MnUEgrYvZJnfmVPEXZC5w/zEb7D0vvxK
qOBqARDnypjSDgB9m8Yp4PU4jB+ky1KC+wJxmZCOEMF6hSxarRSVDnym89b0wDlbY82oyux5CMvS
xOkV5YzWwk6pci0zXVbwonxI9yp0B8tzd3wjVmblQCqQmciAQF9r2kZx4nO5HqpL2yN8sF2K6TT+
QlY0MUHK4Mp6eB334tx6MV5/C9DulYYNLk3SJT7cVrqg1f4Gbeop9kK8pGWlz861JaX5tJFWR3BG
F3yHvzl8KBrmzW6MetJYrohqp6ah60lWAPegjrw1y3a6/cR56eLEU1N8AoHkt+OyDDyAUu4nXeTk
hvZFPn6PldKed2rGJduO+IOGgEjSsL7RovV4UmlzG0ZvV5OEzzRplcMStw6/E9DG3FLxDJDFgObY
hon5YCzZLgWcwlfd1B2sF0AYq4XFHZik29n4I7oARnVtFwqMmoynz86mUuTG+gs7LlrDBAbBnnqr
QBNTOODanq6Ys0FI3Wfol3gPfr8GwE3BnVqaf2TNnztRWnZFwTKjpWEXWL/Cub1FvOOE2mSMgkZX
oQH5YreYl5CtHrPB0BiCwWvXuZ0l+5UUwmQETXP1yR/cMKzXl+Ou3OhC+9aLAfr8ZzjSXfiErb03
LVEeeOZUhuRUlfDk4XvHYF9Bs6Qv5cQf1tt0WXIkAAlP85GtRAYCj2ElfuJ9vCoEDVxfT8zFJgsp
uk4eqLMWYlxdaO3F4yf7LECkibeCrkvWuH8njJBjLKcNqVowqxuNsMcNWDOWoeilBUdCLa3tFLhX
He0YSpQcNUToU+RrO3doSLVp8Ypaba/dzsCaUL9fCIHA9mP8Jsx+jSqyCSUvf8n7Wqu9DVPzYgm7
1lrQr10KNda4cHEPnKDuAshe9Rk4Oct0ie74gOc6daMDa6xyj62xbgT4VvAofe5ciPlMmib8vG8c
akyFAPCS6w6yvSC6mzE9NvahLxcrbN3hAvzOTzzcwOjFUqOEVdv2WTmTW3ehqnKMWuE+eldgqLDm
I3KbdBsKUnBdhQ+sj6plD+eOIjpX3GKFN4uP54a/gYmDTfw3GTMl2B9aKwq9NYeuLKVpbr+GEDBQ
NR3SKhvICW3HOkT19/DmxZH6yU5wTItszIV5ATqD7WlJx5QcaCP7cMUDPfegPLmTvo8/b0kcSr1W
g+tPsC3eJML93USnW1oFilU8N2+zYIvHY9gORO/n/b5jXZxVg0P7kzutnmsHSB+ZK99f1nMpMEct
zkNVsew/F75nDMxgMVZWA1CbZ8Cil6TCkuYDedlny64+2Ryc91IxhEq6IyQ6CcJa25TUeUBNeC0R
rHhwWH9xHjs4zjBMVt/d5791fDDmc0MIL9l+23Xw3wQQEcdEINQgiKBKPOBv5mN9svpsAH9Jbpys
C7UQq2RKlqot2xtR60gwXjH19xAPN4jDZvaZGC2+1GSzFPtoE+xCjQQ4OE6AbFd/fESDu5EX25Am
W9GV7x6rRhU052oQ6W9Osz+D05EQx7RZI2v1b9ndoYP3XJ+TbknnvyZaU1t/uFiQbtvXo/Mp7N/M
QhGZ4QNW7z2aFLU+txKKfU+zQKrHaKSY4ob0iJUDCnLYPUJ2k1rAVyCzhQXgfTPY1uswGc1fpr4F
3E2cJ63YAa6fjKg7sj6Kv5+DXkc9l7FZkbug/I35YaVlvW7ZaeS2r4s1AFh0c4r4dibdDBAYLrYe
++04v8VgqSO39jhzR74d3OxrcEX4hks30MZ/eO0m5Yrmft4vTEljOh5uhliStFvqt/7ZPPsZa08c
SHCl088rguj4xL7m0ZlaOXDnurpLckQ+sjPMQntirYCajHd8Tva+EJJFLr2GmxWmXo5IjRuAQxnU
WiQX5WtX6SJXDWUWNATihy3EUl8A9xgHGVixEs6hqGEmYialCykIoUAxMB4AbtSrYD1x3jqoFVxI
O7VVnDSrhTsPmbRLvnDWYOW7hONyOogfzlmkd7u2i+TS76eKalsdHeEs6NgIuPRqEkYQNX/jXdve
dPaFHqKGezsxz6AvK06tjDZv6+w4i7HDMLAvL/MSKz0LbscsVpjwHXiOoKkLlNF6lTK+B2oqow3h
cz2+Xg9qO4PoHIVghjxLUJq3g0oPw4oSuY8jXbfrFYYgs3oKcrTBMzkFA9kpZZMqndc+Wi9kfHGY
PTN1+2UG6X6wFqJLyIsM9r8w9iFpmF6d0wx2WOwXPzs8CB4kQYhSw1WIo07mHP+Y/JlpUVNmjHOd
z7ynW2YbPGa2SkA0/Mq0vGbSaUCgIM1u2c/Begumvang/UpI4MAfVf+3nHgzawfFafwzOgrIF9te
io1pHMcRHi/t1gns91ilPEoZfQId/KSeLubblxoiozwfAj6JdXsSYPZjZJ8fqaOU0UidGpGDthcG
ShJQ6pof9/z1X7ZUttD5tUiZzvz29C1hP2ODH9vEGjsVk13CyCpRT0nu2Gu+zVU3RaVXGAKC36eB
po73tUfNnfFv/Gsuv+dZxfs5Sh3Ar3MxuRwkSHivZlu3rtnEjRIc6xTOKCaFij+6QMi8nfvw/Bbo
PmtRIC1z8MWZm2FtAuDJa/nvn9D70Z9i7Leic3rpDgppzKo2vnte7HOqv1XcAZDb5zZYYG162aNh
cF/CPBHoswUC7swTNwGR56CTxcW7iNaOHc9hml5QnOewaD4ku1ZwREnZ7USSx6yK6sFV4+zzuZ+U
1xZws4b+mPM8ALPujBHCXTTJ66uPEyVEo1F0nP5yKDhxEkD2P/FsyiIQJRp6c97R5L55NMzqX2dE
/9e5M9zG8M8TLBz53WZtZS1cUOyCw2FmPsj7ScK28rBH7KtG8FWxqN3lCJG2OxSWILQsLRmLxVtp
plniowH3cQJn563jDTPJjZpH+vXkYjPohjOvM5NufekBg0YG1173+VMZRmCe6meupPYTn5t/rBLr
+1cuOybIlWa9G5p8V0nt2eRcxWMwD0OMhi66br8ySOWiUikdYcgxq7dPJKVCYBL57ORbSzQe5I1W
0ywA/tQRSgFhfJBsObol2CNVvIadHEbZok//keXzvteZ7W02X/2U037I5tf7vdOkMNanJXbcOE22
ySj5zlTwi/H+aG4XCsD4WydOrAVZbehPf/J8V0/ZRnUzhlc0jjzBwTqv/mXYp5uyDJhe4gTiXLcd
peEzvZ56MVpFT1iUoch9arjSEphclPNdJWU4Q0lykkV4XDWuuexD79Us0Mx18VkfacP9rcMP5YwL
rIYlr3nsUIUYvZWv3rhybEDodPkwfaxwc00jecO3lLFlOYryeHokSEKcQsfMoBiw0154/i/B3AP/
I9Ez6u947xCu1ic1lcdekKhnTorLMZYXoJioxpluAEUrfnuYxr4C4ztma9ehGdVySyF7uiXLSFKX
4ck9QyOMt0gDIPnPpC+HWZfPOtgrfxEg5O6rOoD/miYv7Pp4wZIUIkc65SdqQJiC1H60WF+uu1wg
DttlsyLcxUWt6ELuQm9uWas1c5EciLqfutxYhP5lLrDOkK+Kqzq6myXv2LyHnbWbChUPYW9qpptc
8BsFjvkDiGxFMxcm9q2sffYTILCoYcUDm0yG6zIRgOVbdNM8VkZfgWfNlJfeRfqauI9jT4MQGVPx
/dQhKeq/myRT8y4mKS585xfthA1zZN28DabjLJab8hFMTDNBLQj1mYxqAw3eQdO84GDnZTAQifrk
iw6uhDSd6qs5NYRXSWNOOzU2uElFZs2l2hrzoaLf/xqJlg1vOoeeAshg5ROGxJEslqx8ukX5eb3h
zB7V5jCWRCb03G7/TtWFD0AlwB857jmIUxOIMnnh7KI+RTyVfbwGO1VlOYP21v+nmR0dkgVP9Y1r
EEcY0SA8CVsDjKe1/OXAzT82cMb66cFhhuytEe2mivIpZcAYGEgoC/XxC2xO+H2QLzsGRcVlpb05
7cp49TMYVAz0MRoODHX6X4mEIKOmXXg4KIbdIs3gkzGa0y7RbFfD1yLzJjLa3+vDhnW0Vm9hja7Y
OX5YH5LQrT2L5uIhS+HF12RWMa/U50iiFBtPPZpzplMjwde5dLuKZ5Avmg0ydGSIJERaygv2isQw
Up1pzbF6lSj+1fCt2IKjcwDoTyAMouTGerNyHL0Sb3NLPPCTYtPUUPA+FFa7bV4sJnIO5ipnKeDX
3NeRQCHTcCom4f3zvLwWacT2mTNZZi70w6aU53wDz/x4MQfynVPA3WIMNbwZSrT4T6dXnu0bQ6v2
wpC4mULn4XuURsSqQzMg/1oTpOE046GKcuQeAUA66D0dZI/9KzCYfCXkeljTdRWe58qRm6b/Onu/
UbJULeIwtIguXN46anVXpVDBELAxc6NhCzqXfJIf2zesu00Q8yBrESt/N1Ny9B+ezCVnU+vp1ERx
pU1RQ95smsjHeGUy0TvqlSDsezGmM3d7R9vLotbnpPCOFnxlu74a9v32/d3VuAazRfQrDS3ttdoN
YSRAWvyqtALwyybKUoWRglc1xf3rlkxOJA/xQLthuXo/lutNoRJ/rMR9xkXUIpNq0ThNdQnWuo9m
kLtIH1SriK6M1nI+bXSGRGVqxb1wMO6Vj8WJXy9g5a2CPXpKzuM3YaPOPZxAMRgcMzn1mrlOCXU2
dwev9D6WNoYCvYA+DRpH/MmuAd31MRuR6SK57To0xJB81Kg+jQuI0MO3zeshMkCTlj13wk7uCwBa
eCqvaCdpV6H44kZjK7bDl10wY7DUMQX2V2WN2DNv+kF++cmXQSopvyKY+QU7GeUXOLcUAtlaL2b0
+HHQSqPAbTLCYPCJJuGR/g420Eb//ed444UnBKFDH+8CkXK8aJaCEPr36oOqut0ExzUVE8NKF7hY
r0NKVmo0VFXGxToLDUs5jBOTU0We8boCReQi7R3CIgF8CuZeWGi97k+vdcmK6uDokNlnxg17cZLH
JS/XbaOaOkuGzT5ym2Xzw87gSNO8df2OfuCAtK1UP1ooL8ktIuFMLnVgDKDDv5ZQuJCP2NYyTl1z
SbgDEx9V3MhyAiLtLNMGiSszOBUi5jaduc/mpRBWokNgi8sgJzY6yIjX6E1q75hJpHU8IqM7NL/4
gusVAzQUmVTjGwBVd/MBbsOPB+4xeVgiQ+NDapdNz4Uu5Y0d/0G33/qA8WdWeVuuOCMxaaXIh6t7
V71HyebfRVxP3A20GMTYQEYthI5lB/Fg5dcqr/68PDrA79fRQr8Gh2G6hVA0CzFs4GdEYwyZ0luV
UEJxyRTbop8a4ukOKLIn1eEz3fjj2Dj9SboyJnZHAbRdOYRymsVgJQB22Ui3RKHYGr7I/4RKkljC
mJIm6WyEXvaRGKEwAlFXp05Bw4fKFe+BfCxtvVJZN4RcJemxMnUQO6BD35nkLPS0Bm5V0dhCtkfH
jpgc5ufAbtX0F6Ss/0GP8D7sraMPLFx76wk7TI3doWXjP7SAASd2elFTpGWU91zKRUFOp6HIbBVb
zmFbelOOTD2Szn11mN4ilwPVxPA2FuFhPZ4f9KXITZC/SuwYu7dyog4NSd2FkX4WWtCG9vnD8QIg
ceiLdm3hPYoZiWAV0gLUWpgO2Hjpbg3pe80oEXdTB3QRVADwdxM5XLQfj1vmfWl7BVROHjboMwuy
jtlF0tSMiyowsVXrg4HKzRQiS8+CvRBrNF9A4bIQ/VYvNtMa00EmL94JN9rvRm7iOJWkVJLAMzYv
njWU+UWdh8Ih0Pik+UC76cDNewW8BfQOZBdcmR6Jyc41/YBl51hWQdr4naVNTfpNql5meboRAxOU
6aBqysPgN40zsLEnUW/IhyjgIT9PY+PnqysKMhB3nW8hBj8cCc/RHjPeH55DVkwvHtMKnCOwPX5w
88wszoqK3UOTQLPRGn+LQ9fkmTZf/Rj7FbhRFylGd/AfP1MmqowgOIH62dWtG0evspv7n2qDXuiB
9f+5Ra0lE878NdqcdOZUL79qjsKAudWWs+62L59IwbgBDmBlspKcgC1TK9Pc2IOPJsTCja3+89IE
GIaS/3JgCEZ01nuWYeI93Bf7lCNn4Yfd8pWyHjPUkONIFw6UAXRNzj8gHTx5DgnsjTZthzA4QaB6
x/D9nkCYmU5HDxtctNFN1ATRe545UbY8O7zj6QS2ISwj+HQ8de3FdyMP2CkoNr3B8HO5efg7A7XO
pfG2FsdnMY7xC3An4Z1t0njmwVN0WyfSozyG3E1apJQWz+wgsNhT2MGcfSK19yiqft6SyiDcGuDP
kOC5K/OtjiKnUs3fALzCL3P0Q4S1xdXDpJ9PP0EP3ob9c59Zdj/6x7edwMWi3N1RTeuIB6lVpKnk
Tdomrivy9B78doxX8gqMS9h7w+l6GkBZXs7zJDi6xNzY5tnEI8vf98CT1GC3ozxTdqcEcXpZVVTm
9nqvTNLFCKge0TfBBWUAwyOuhAUGPzsAkwFFCmLXT+/YBNME4/cVTmGuNh8+sGE7pByqVzsFuc1X
SmBXcZL8XrHOWTSjbxOrlXBjXJ7bW7b81Fbkabk3PCDHawZJQPjw16WRCPvTqgwvzHpCHNM7AB0y
gvab7VhW7BvTKBEcrMGQe5p/96/4VL5Fg6OaIPCmmefSt91b8CPVOHD7UBZtKvmDZa1rJoQwNusz
RqqMt+f8BczasTnQ1wNWD3TALH4YzVike/lHkd5Wy5M3dctnjnzRUU2KLbQVchMWoJ0DkneLtgPz
6ppw8o5SkmtfG9yVyxfaZNSfSrJT11Ke0MQ/42+Ew6PMPiDyYdYasTUWXzjvN89gfu/HwPPnNdCc
3YwIAWgEVs0WKNDNH27xf6D/z29rT2AUdQxD01tUnnZTd+a7s7D88kv9q7A7roZuVgh2fr+v9Gq3
RsQSC9CUUyFkF5DwRdUs0rQzJtip0qXRq9TzUygGZsGOpaFHRdAf88DZsk8Z3dSqrYnKjGAiNN/E
5QRYHio606Nuyy6hEtv43jXXsN2rScYgV0E6hh0blbKZfezfTCdl+8I7LNWZjD+7P46ROoroz/Xc
braFYP0nh66gnvSjhRTvd9ZkqpXDQAp+deBMU/V2Jv9n7MNSotzfeXmHQUZHfnQt8MUHkjJ9fR5V
BkNq692CjPgcbZ2i2/mrBewInJA5hPHCsKZ6O/9t4++TmrwyAb0Qqf5DSXhosxthkXkxtJDt1hI/
Xn3PQB4KNezYjBBC4EivpFg1zLkgCGDrDj+/ZtIAOlly3NHD5ONOLoTNS7N/+SqMKKwnHawyiSiM
zl2fPsHZz5VUMzhGlkdsV4lHdOebRHAduhVY5JwcN/j8vqqF4ehpL7c6pWDIigl9U9tEn9/KrNFR
tbV/sHdcjbRqljpAjER2Oj7hvjGpDPKbWlo74WGMoG/WBm4YMqEy9cfcLnsjTkdaB9qaQZ/aVhLx
na2bltsDdIVbhTYCd5TLnmf0YydvBxKfyhvGHpW/bfSo9tbRhVCmIlXYr0Vt+EB6EaPg4jGN4fD+
s32bpm85R9jifXN/qq8Sd2dYpnZrucCofKE+KSSzOGTuR93PZbbfAMNnYKWGWWsOPe8tvgNzVHS4
irwL2dXbF0iygORFEKtOVJtyTClrGNwc772T3+pDSe38vJwTrLfDvxCTJjzpStA5woS4SMxOKpkn
dHQ68a35FOas5qJFqQ7oCDLtQJm2hWVN+9ogW/gETwAsz9L9b3GBsMnyfCUd9iZvNk/UtoDtRGce
ZYEDwZ4YoZ1hGFpQgf7bBN8yZQ5shV9qTLEeA0mGqbxT9ECFUO0zLLw2ZbHYdXQ/jrK2abcH59xj
owg47sFi3OTzzSUo8a52aunv+dR5wpIfF0OW4cWzpQkKZtqDadDtINNjDQjNjLqYpjv3QXQ/fu0H
OVv6Zsnz4PZHhv7Wut4kx6rJmsNYyygpW8TH2Tzc8mm+t7/g+iJJEKtwzMgruN6BAhIwFvxg1iw0
EJKFK9PHKGBPnMk54uI/FHeelFtodIQpD2AeMfpNti7gEHC6IuSMjhbj2xAcKCo3p0l0x1Ko2gH9
nZa14Up5GCC/cuRm6GCsTevzujwcvMpMBv3cyZVkI3iXVI/OTIvCJ33Kb9StT8Y20qu+x53ZvRPG
NUBsmqZ4it671iv4OlDSB34IOwAoPfmVHuXVfvKQ22KWXhX/hKH0R3fGVTaKRHaKZP5FGbzhfLpe
numAgqeOcZ1nC/0iENoyEGEgd3PnY+J2Dp0DUAgo9qnn9piBoeDH2l40aVukdbbS4MVBxHvAindX
luJRWEvEzmQe0yrmMsstsQefvIyozTIZpWeFXuh3+V62bIu8zlegWQTQxi+T93z8W/7jVsn2rPCN
skd/EYYO0LPWP0SlczDMYkyIuitH0JTYCE7+K/lw9Jm2sFsu61A6v7dGnjHhB/ApH8UUQvCbLChE
JZs5DAeVnoTq6tn8mQ+kNkP8Er0M7WapgurtwGJr5eGo7j289MwhJPa87RKnSSN4ax5QGy2RV8pn
FzDqlupKpCvDrrrwEPtsiweqRmY6oWa9ovWmDzjm56UNXsvNHFUis5Qh49XS5zp6tjoRkE2j6k6i
U5wERM7GZtdowFFPYflgI2r+Y331cy7W2120vb5sL0UXAQDJfj6SfB6lunlmSMxnLZXgYHh8E6nA
pvsivp7sDjo01HgHmnAc3Ef8Tohk0liousWBXrKaOySQCYFR0LQGK4YujRXiGvAuX8Zf2GdT6zmJ
i8YH4gc0NeqM/6LvXZGrPN06gILcjUPI2J6PNnCXmDSVnrsLNhatpVIoCtdmu8eAU6m+V79dQCt5
viZp4phXqpNUa/f3qWoWT1C1zdxyDabvhkFMYJT8dVFosoS1WEhg6R3d65UyMZOQOuRaIajKknRU
ds4LFfPbhrBvpNkjL9T33WdjFZYlHLVCDnBnFyUb7rsbVVeZnHhUvzhd6WGfDEYqBgti/Y909Pnl
tYAOSvloTRHpYMQul5XWrccDZcDh4Rl6XwMibPs0d0OiTy6TkynmycAZAo7s+sCEm+dPIrh6hWny
JUe5uBxsyd8pBQsOoGCLRSwwVXo/UqPm1MAx3HhOIaIMXg3ep6xkSqHCVqMKTdCEk2c6Y5LkU6z4
uDTFiQ7W+nuwBRP0nv020NAZU/Yei3plDSQF20YUeNSTzIkoaF/q/Pca46wA+twwD2Q2as7CKozz
Z4T1Ro35ZAdMFSbR6u8E+EWyge+USmB1jnJgLOkx2otlF/FB8gua42qgCRZIlL2hSLRqsSHP1hb8
xDJ4SO5r+CDgPyrrvlsVPQlewh9V+rrMpSaIj5AlfSZuJo7Nin0mZjjAR02yMuou9wVmmrm/l+sj
UkJfau0IEoWh/mejQusDa1imfWPmTAknM6FYTutPluMFCc4aRG9mCa7xKUM/N9cj4wlurlmm+h0r
S4crhPNK8i/ILff8EdK1dCQQhqqkzHFP1l5LGAHvbWjMNruSQyXRXpx3Tg3olnVhN7mJSIhPwIIz
kyTk2xbFn/fhDDsf3nhaTUcSAFjujQkUb/1azgR1WuR816cs1LaXc6cMBI0gQ/NP2i9m96KU0tIR
Zyx5vtWO9tSUbKrDZe2Hk/+qjInfBs/HHenx+eWzQvAthtJhFUYNNAiq3bSXgG5fvK4Mm7gtiZvW
6v4aG0guWH0johtxLvMGp/6ZGqgfVz2fuNAE76souLudh+ZtPZ5/oJRMKiH3GZDhAIdsMt9X68Vq
00b85OeSziWZHCqs0ii7xC7XVLCxndsZNW5vccUuh1/GW+2FCZeq1e4NInGTVFmepwj6Qowc5mmu
v9NxJFjMmxQn4/URzfbQmluQYWl2mOPzHaezw1JcpQju/qxo6ZnBfilPKMFbwU7/B107Zk+mPocH
cO2ngoUQck5EL38l0MRcEVpavWoaWkAzvHqyLZRdadx7seDIj6AsFFxikbU0CvBtpMaoyf4rgH+X
ZIufMKQka2O9snFXWU0i3PtKO9RVGuPTDefvsCLBj7/X2oLNdWDJfcFGaLjMR8vJOBXHL9DlH2RO
MzcdoUfH4AWfch57IMnIOJGTW+nAGrK70wEaDyWsbXLjeX37Cfya9ZqIL+DVbyw/qtFL3XYsODgW
7Pkdlq5i2Z1MJRNEHcCdM12S+kEdBJJD80UD6KZDmskf3QrsQx3ysuIQX1orqaq942nStrIkj2jK
JInJu1qYkICX/MlGS2CixcfNQ4jT46Ns6acmZmsM4AOmu8KGZk+4JCj5+TOJojwGyouxRFihtwWd
B/5GVGNoBIVw/biDhxfk4neUe37oCsM57y3tULvxo1A1KfGdcjXTPdGm3qRm+mTTv47ubAFFY3iq
7ogr5RB1bXmRRSog6e2U91djOxYlxJuHEJyFCMqxX/ofSnK/HCPu5A/yATy3kAl5mGoYPkjWnJiV
sPnUnbRKhKwUNSYGY8n3nGYJMnkccVjNGjm4M3stH0a4AAGl0aQMWyWVyGlWx5UmQINkYKwbnLnG
WmJih98SUE5mjxdHnLCcNX29o0IHuvNTc6CGZj+d69+RDJ2sLOHkrwI3e6fdY3vPGIPt3UvfOiMK
Ql8i2YxPj9Ou0J5D5EmJqJGtYd7ZV7hS68GlZrZfmSHkI+yJyj2HeRZXxpsCZ+FlfVnA8//6ZrxS
MjR0vnwUK2MymWJW0iM8coTLQlHDw9DSJTIJd874273/oExSEU9W0k+5yiP113SVh4k/kqCtH8Qd
H9r3ID7ShrBo571AGtoB184SagqVRZbyFDagrLE2hJPutQqDRVK2z8o3LV5KRUGirdWepvpkdmUh
BG74AorMaoOjQnh8F2N2hR3iDUJwi+BRL/3Orj7QvRWv3OOi4jxkzzAmd0O18ZNHwqbreYNphzQF
djjXnTGHS4WRKE6wSO1a1l/2cTnMsrJSlCyMy/tQJ4leUUORFQVfd8MBhzMufUCw5c60KApXg+He
gbvrg4qVcfVrMa/z5UObNXrsRiv5q039gVk9mFrTk0WW6S+6ztwjLD/OXZcPsvaJDuxO5oIW02kq
lmnx6wf+sOf8hFMqH8NLyDq91e1WR4Xb7ZB8CfmtuZj/LtW5q+rn4WYINnsgkuooijTrEeunw7gV
NlwKsjimomObfpBiNDhOkt1636tWgjx2ywgCo2llUZVDhByilfBkCRSuvVhm/tDEUPfIoNBYASqQ
acJNuAbp0TZR9fFjbDVtfrALY6EkAnF2+9CmgSjggRy+O7ksUofuY6NGrmedzvfygSd0ThPsaLEv
lAsvRfWwPEHA3a0680027DXJZZcHraHkzYpWofE1cAxSajMA1jvWsYe3384zAIcRcEujaxoTKKjo
fhfRjhXwGeEOYnlNb1I39jgEil2BQeblIUTig8ZNYSEc86PG9QoU12PwU354JmOb55QU/ZHZMsi4
ySYAExtci2v9fdjCKC9REvWsznIN0hX19Z9z4QLQl/VGQWHtNQLl7Ofq4VPDmVQGpu/ifDoA3V1w
e5zokvxUIZsv8Yf7QUBvwI+gBnFdxoNaGxJ9/Lkmo02Z/6htGvPNr8TQmXTbVjsCPdmz7LHxFkkq
8raGx+5uz9pvmKvhkD0pkG3psgAyjsAmCI5JI04SbaiO5LLqyBJ2mW/aHjjnbv4Qip9awIHqmAiT
/Ao+Urh7WBsD6bAsUIQlklMMERhcz4WcRgDWMSPwbru1ickDlHwCCuc+VP/uAGfwjEGI5WahyVwt
RPyE/Yx+XCawzQj6VUEwfmckm77y+B2ryN5nt6gu300pp+kw/fp0EnpxR4va++KIG+qMokponzzN
6MwHTyyUEI2RTN5N3Csj6EdGAwGcFqSZvk0rzjQgyU1FkrZDxEhwCYZk9Sup/NzAd7KiUBjHUsk+
K+sqOHwn/Y5BWUsr0Jcz8ime97BUkt3FBYkdUXkvNjSbJ0K0t5eyHfI+Avh/ExWBHX9LzM4CMAOK
EkBx8SbRzLfkHeYsfQoHBT/36TxRWN/jQfP9NoHZlcrkcibAMS4ajf3oSDj3ejCsofkPJsShccKH
2KgmhARk5gJwwrqbA4otkj0OXeJgnWrbgsWpxMdXi8y40IGfAf2i05shrjhix2HA95ttLWUla/Oy
ujnQ88OkDo9sM0mg2zXIw0KHFibvlf4K21IU+6j3TjBVme5qoT3pGVm57gqlp0I3bcjqym0Bz2kl
q+VEY98L7vc8R2Jw+aZ7arxvov7WhvtzKpP6G312P3sbDAw5HH08tTmFSSoqlVLk2/I/9hsAbhNn
l/bGqT/nwTmdzaaG7rmTmLfJkiBIaoecRGDth1EHemlg0DOgYxVaeWHDZp2G4njtCMdwbXDhiHQs
VoPNrX2Y7T7xr/FyPniyPaf8NdOd4kHp9Y3Vhwnvyyr3E1paMcS2eiJq53wAqmuUbD5JKxGqs58S
T35zxAOUXWlSqZpY2Wr3/HSX3muMy0g0jZE8m+ClvKy/F9spfnpZzNFUXeJfzKGUxC/M1fN9z5MR
j+oHujnFlssQ5o84ahzf1/GyJhEzwWmiC+Hf1AqF9yuky2DulLkhjNtru85fNG54NrnEwojdn+Zi
uRZk/Dr7yEXI7r1Sy/WulOcR5x9m/9raUFtcPSlcfa4SGyPNDunabmaqdNufzhjsy9fcszO4LxV5
b3UgWXxSJSo83E7XxtegeTd/tflg0Ytuim3MXtgd7CE+QQay9rUQcRbqZvuNjsySl74RcL2XEAhW
cOEXjHzD965RWr079zJ1EFl16hKFBBR+QQvMsTupIO5s/lH956UO2IQvfzprdkBmVxLvNYKt7G/9
qxrFA/ahpunxUFydQoA4UOiaWjHorKPysZ+5aCPpt4LYMCQbb5Z7A1Z+fkwtYBL8/j5vmnis4XpN
ZOIq1CoX5Pff2lDRwPaFefzm+/X1NTskMdGsVHfp7+newpUgA5S4+UjisnC5kSXSciIDKi9lHF+e
+Vb2d856vNLNWbGwnSQ+m223q9wFPeK836mZFF5JUaw201M6iw0chPXay3JbigOYOoFvGyFhE8IE
shM0TagXF1rlnMoQproYR0eM1ulxeWg+faivWMglEK1X6rQMHVpAWuKx0855wy8g2DeDPW/0lroH
HLBH1AD8YGJUokjXKciqbEWBRrwpfJTFrqwqfEg9cNyNQV0fLf8zYDeBS+8yRBiSGKcqz0NvoEZ4
nXWY6WHFl6527/SfEeeSeTkbA8YPU8n++nShY3g5qVv5xl/K3PZvQYqDPmOR8RLWp02xEHDfpW3q
fV/3FpvpE397A90dQVOJMrnmdHBxEPSINz/EryMUzHM9WHfrIjkJEvWZwa38M23eh4GvmHEQ8hFm
z7+DtNziwDmHtPL6k2N729KHODNu0P/zVPjz/gzmdOmNm8wcazzyjtNV9Tx53PXg8S5IEH3e448E
gwv/XS8fzKkQiof2SVjwzL4kBwhS3jDtADrlNrdhA6XoQpcTVS5TXqDTUVZ/9yKCKGYg6RqMxOhA
2bdVq/luXyw8rDgWOg0hl4JZA6+wrTWPxhG+acELo9ZOQdN36mOspUBdhV5vHgPay7DIbxWeap/s
lkg+Twfyi0PupH9WeLhzEtRlWkU6vxegXzDfybCc2GkNdv1ecjaj9zGnomBNzoudEaSfOL5+SPQP
Uf+rHOVWSGOuUDAOJNQtp4z6Zkn7PKIGf5E+veJQtlWizhg+NhqJt/7KkVVsgmfVJAp5AjyABX3P
+4bQR4OWGE/LaVwRwreashy5C7Tjj0N8ib0M3ZA5c8K4rTNI0MGRf7+lWlkYQa1l9Tz5xc3Q6Rpb
MfXV04158TQPCMr2SeV6u6nPQfIYHy19id1n3Keq76rzdL88NEFfawpMlhnoLdnIYmD4e/ifzere
cISDWx0CxxYTX64/Gg/qfA0pfDLVc3AKQCPk2Vwj2Z3cDUOUuZ3c6mkFR2U/oLTT/FQIeuF3LsIJ
GRp8BENLWuXwLuzAHGpmgpsMQgKMQ8REMN/nf6T6oCfgWJz/0Koi3mzH1umvENbyA3T6sHYuJq7B
ZPrxZcs43IN0j7VbfLJGUJ5z81lOOqUx+n+M5HsZRsQ+6xaHHoFyL5gPotV9xY8XThhWcZjHlP32
akIjYBseYiQ55HW6vGAY25BE/5+/58e/ePNszB+8CnfGvci86h9z0cxux47tyrEKoS9HRMomsfoo
J+ZzfETDfKyM0cEhF37TbBRHA8kxiVsKouSlFLRCSdweuNqNKnyktUdij+o/45I9F4DOmDmWHe1x
AF0h+V62uHbQcfYD5O0cgOWqTkjh2V5gGAACZHUUhDnwIumaxbLYlReM5jJwaQe7Dac2YpKBf+AN
R44Cu+OjK7rtk6QukHz8DUwNik2ucgtAprQVZpc5CBkJ6kZrnpjaJp74lgrHEWB6lfQ7hT/PN6gO
MtdRd30OHqS7anJbiw0q4OzxxFDnZhGEGllLivwOiK2pGzTsb4XK39EOcEqwOrZFG+X9UO65Mkkw
TimguluEMABpyr9zVQhcu5NiaaY4jAZ8rfBsV5RXx7oTEMx5RYSP9dJid2Ny/eNKH1UWS368d80P
4EuKAIHf0FZ+ofOsxYOMxpfaFivV9yKejeJXGf91zNUVkjESNfxAJj0WJXm7hfkoJxiS9MTHVfr0
ywFWlhNO5Xdd/U1GB9DV3eH0sFdXnQ8CHPaAkeM+C/YZ9hQeSyp8NUbt1lsezVcMJuCZOk7a0kQe
cvWn2BoaOoK4i9muqojbT2OWVt0vi7TrWGZk2RVagYf2lio+5Vgmhk0sdbPjZZhJXEvV49Wdmi72
rkurm7E1OwHvbXelS+rYROqdEz0YmpGn/OiVGRQT2xBFolvUoQsL1tZtTJtb1Nk8M46wbT+vlle5
5y+tePNPZkKzBAwS/WLh1NXkPr2JcJr4ho0SGI5SX8pOxQXea/AKdoj6DDRBczzp/HbvpfIOD0bP
LnLDOYi6rO5X1Aui7lVxDKHXlrtShFIFFVktPYEoVD9efqcyo7PWV+2rYjuf8OMxqeKOKQ+KeXSC
cSrrGZCO3RsTT0Cti6guS0xduAIEZjWKsU3AI66bkpSDq3OLmOY8Vew94cGpZbTGamSMZd3S/mD0
4Pdjwu/EOLrnjJQi8ATqFc32trXV+BaG3wd3XrL3PfpCv/HPjCyi9lEIt7ffjwkiLY5BRA9kayNR
cZYGqKlioNoZz2IWP8TtYfsXOY+4vHLNGxdfeWjU8IO1MabZ+5gpNrNUDy3R6mUNkmci8fMKFCXW
gSjqcZqp5MNzCGQ/LdI5PV6cPAe3zJGIzGrAPb5gKk1qeaEKFa4ooF8cYzZGcLitaz/6fBitr8Nv
NuejBR42Uch0HwJiIBFWuQk5bxZ0NkmIhA0tEA2GvZXhoyHUITlnz6UfHqRnxZDbYih4rlOHcvHw
lta/hCEFh36w0VbdLAphKaAwZEuY56ygdSE2ZHVQqbBuokZxqDFutAc/uKicyl5zAIfr2eSR4Qzr
M7kIRIPviRF2MAor8I1ywrWVDHpX3B9rVJb5DsDjQss77xtdprhxJCbsxuWRsuj0DDhg0802TBNI
/9GQTC/sjdihJ0dRLoobChkPxO8w5QlS9nRUTMWM0LoNc1O2Kicll00P4xlOw1YYAvMqIWFoPD7T
T4/W4PmL8brkeBHFlYBLyvz17SQW7/6jtaqZnZ2FwmFIt4nM99Bw3fisn0c3Fj78HrylGF8Y7o84
/jd2+hLnXypAu3F5Jlpq5nDy/uYF01azJwAJWIJc3grVUOVitlP+r+LxyomFA11LyeRweRfTAiCx
QIJDUPtFSSp2LY0OAU9dWjNMU1EYRiBkrksERGmVZswsC/fpt0Ei1d5kb6h7btVFB3FL2V6IfKKh
oB7Vrh+8FKf3jeZiwRH+djKFam+yAWHdeXXyRTiSB/vKKleGubjRhlBCYEbvsGG7eUGk63WWw3pk
4NOZUBJCDcz5bDInb+bcfsfRW4UE5B1waxteHsQRZDWFOt2goLru96tqmm/tEEMt6HnMuJL6WBGE
SFbMS5cBo5xpzfOInfnm34svyE7YAXKw9cBU+OhYalNYXn64C77Rv1+IHLEHgC3GNlWZbhPRGayT
xWA57EpfJx4fV6RZyUhDCdpwEy4T7rf9IIj90wm8lLaRGy4Yg4UHYcL/YKWDdhtuFc66NkseTyfb
1hghc5e540sGN7p6UXiHAfbTNmvflfRssbtBsSX35cWjdzm+cRVGDOJVNQw6efKNQJqfT7gR50dd
tHCjK61p1IJDE+LMM+tIvFGO9/GySUwiD3QxCtYIn2YEJTyHGF9Oaxy5TxqAG63ERSz2zGu5tKFI
SRNqlFPqEtEMepXV3KRi+pIFcsIectpTJmTza05HS0fxVxkLJ2YGEs531ty0B/in9MV/49unBJhd
q3liNquwmodQUDns98hsNGmKmtwTJgcp6OtDAO194Rzkeca0sKOE6rBtBiPSpetX1YWjtt9JdlCu
XZzYi0gonZf9wbmzBwZC9UctEPPv55D5HD7lul1rCe92HDqzLIZxmzd9BK51z8bC2yA75ml2Pm9y
SpCCvusiKvipSv4O7XDrUjvueeq1MH7aw1egaLxws0CT+nax9XVrM6RElYkMsXR5t8KuMwLMXLQQ
OU15I++CF291CLu44+zLI6OeXVNC7FMSM89HntE5r26feChmD640D+AfCIoawxPC/yIIGVgEswmR
DazMFz5FwlgnOkzaqTseEwVS4upNpbC1mUZKYM1XerP/X4RhlDuDkbaSfOetdyzOn2YSur6/sTXM
g6AMEfNU8q2tLNqzo/TdWxxwspim5dsrccYY+NNVho8EPWzaXV9XgpEsCpLNX2uMRGNgaQB2ccGc
62/7yBaxW4i7jlGpZNnPC5lkoYBi7HgFBsRmXcMidFncmkbmbVYXpM6pMfUSViOsBWraqdZUq1vD
FfBhAsW7JGsWbD2E8UExveYuEo58WmRXj5JIsmac+pUqMRDDQDLNvjIVfXJsbI6MgsUbDg1yML/E
jlN3QHESDb27QYXbNKn6fJgbgj5gu1CNIpYZ5GC+j8VPsvGCXU2rSsbiWvmM0amz/z3MsQHWnxkl
1S9cF6VgrqGYTRzg20zpJyJDGczBKQi00UMkks5m3H0Iz4IpbtbDjaIRHxMULLRgJs8eWqFU2Svr
RPLzQlWL06SDpjSUeFwhucMKUC2hQ4X1ANnXC3+lhzOcKdycF/CJgxa8SVpWvrYIwdnYlwdSRIWl
b27VmjVvc8J9JB6OBgbn2EWGUz30p85mEwkf/F2ie1WId7u/bkIAfzxh2FFCfu0hDEaTNb1/155J
IC8PjkBrtnMXjcCVwBpf9Jaf3Ij85tXKJY1NjRKkEy4z4Bc4XWTWJwCN7j2dmv/PrBOthcDPDnEc
me+loGyfDzqNvrXjS2DTD3h2XXiHBh6Q+vtPn0w8wuPcAiZjrrFYjqokbI8kXsNiaD8tHUYX108V
N0ZUvl+k41iynrXHOOJEVfghYisxReFatQO82k8A3shu3IoUpWxZ1f0pvmYx+ulsUwggj+h/zVnX
XfdfRWp2oIUI2r1CNTLPMS8viGUiLaQc3bggZD+DXD4kL9CXi1UOZZWpKbrvAnXS6+E0Xqv0qQDo
IAmQgvt/+6KE8sW7F0eFc2O/10mMbmkHFaFha9KbuWUjZfKkIE7kyM8tPBaayKaIQQqtzIFPUX5I
iuN6qsGMI6WM73gmsleFEuxXSmwt5vSInWJaEBf42xqto1w+AunZG/kHoS4+V1h6uXo0VT/sWTDg
lrrc5dxN4nC1tBjnzWa+zKhEZGTEIHsea34bBNShENPA3ldTWLUVsVt2TysmNK+we615ZuG0OUDd
5vFQ7/5x+OO6k3m2bTgM3gdXpWQC8mX6viy8y9SHbf1vnxtF4oJcOq7ZDnUAE8UB2Xb+qMeJ1k77
undOxpnCcEyIrix7aHERZ9PyVYBUmIoIxvnu9LqAr85+kbd7IVVGPkhqXdgXhjniqPdrBUM5IL09
MdYV2+m/Q4ev9aEjLbcAfyEzCDPG6fAZ3rw0pvaYzd8jL2F1x2wGSet9pdEsaFFIljwvpeEn4lCl
ODA2OYyDDzHupvv/d7Ahkw61fOEgB5ZLx9ud/WjqAdVk+f2nBP8IHJhK2mCvs0cMZ0J48zbfgieY
s2R9PSilpvLykOBrosbeR8fkyfIx72dQhpZ8fZFGYruF5iufOigkIZemnCzuSsBGv/tfVox7To1E
KTwPWYo1IUcHL0Iq8dQCpWVbjJBQGHNoGNNUl79186V38k7hD0nDqCnC6lkTc/FFSsbWSbN65JGS
yE4eTUDiwl6YEIAL1x4AMuIpSakTnYXKCCj1XQYMnHMk0lPAdUbl9mfj3VYq43QvYlEOH9IHebyj
wZxhttT2e543bIQqYvKlCaMYsJRa2vJTcU/lQyDpoD4mz1DUugxU+BvqD4mg5kWXcsihoGTfunzI
5nHdseYPpWK5MS4eUkS741TXAN9sRU7BDc3g/xN/w7LbczQb38UWmZWiNqDbn39qsRQKZZdc/WUu
rdCBBXty0WrHXkyWXuLSSFLSYhzmkvezEwdavP5R2rTmr0+/FYplLOzPsYa4vYO9/1EywRIVlsSt
6TXf4BDXgVo8IZrYUCEL332RzroIzKMu/NKs9DnsctadCnFiYQOpsrZK/1qXHqi/tyef59tAlz6Z
fFR0/4mDPGJ9TdFXwG2o6M5VHGIj9YQO5K2ae88KErGGiU44/hS+0uD63q2DuuWTeZ1LBCw5WlMI
8R9OfG71A0PAAu+KU5pXqm8uY+wxBxEJjXNzywJ5005dzIRS2u+mG8RhhE/ssbGGw52aBmGfJN4n
sshxm3zh0X7Dg/B6zRWgTK5E/Y8i2Ukk8KY+Cccn/ue+nlxQ+3E1CprshMI2HxGGlzwkOcL+eYwO
bBfY21ogm10pv2B9DY7JNjxUBCK5mMk+HC3T+7tIWFLbRy0Wc/LvSfAjzSKl1tkCafsQxoTx27qo
6K80Fw71hku3SsbkceCz5ia1z6mfsi5RqVGThlsgRwwf134wkKnSALnSEeftdgcpCYNihTW1SlmJ
CLcelcZonWE6TipIgSdg4JsisAGn3zgQ2NGiRdUnBpS7LVskRIywKL4DXSFVPpI6YixiEe4x3JSc
Dml0ivI0erjdZqpp+0EfUFxgbuAMpwewp53DwzKBVdx2XFA6YrAc9xOkKDZHeT2VAaq9rhpFE7RN
gDmpk/47LKSrhSlP8RgrrZpRi5ymQAIrMuS3Mxv2bcpDK/m7D2kDjK2EFi3dXyZekTzl7tyXj0YQ
xct3ybw2YQnY3bsTw+DQTHO8ECDx6J1N9sB1r+twuhdcPIbffzvjCs13tr0pg7B05mRS4/vFd6WI
Tr7TfYqrrvWv61v8qCZpYeBH81YWN6E4v1njRIYPRTxVQUkEgDXBdPvSBjk2J9mhZu8bTH+1ZDnO
JJZNdzDpzzCteToIREViffGQUpYcHCiIKqxhrxqy+g2oNLT1HuLrDpTO3sPPSC2JMjt/th4uFvNO
PT30w47QIUPShS5QiICOalIkkgtJ91LcHhvV647gWki/7Em1jQfczbShz7bbUxP1rgJbUY2t9LBg
l0plIOPDcLB+JQT1+Ul1WiXdccBsdfglAGduDpMJwxDsD3qelGCVWG7RJstGI1AJ7SD3hgEFwO8m
Tt6SFGLLXYUJfdWy57I+Wx08kaAiRDtNQjHLYzNgNHkUS8b3sTZxlo6PWRjis9mCD4es0dithmJn
emRk9lqZkiZzKZK7HVjKbxaHD4MT/c371ayh7y+uyUnmwj46TAy9fDJ3QSxLk2CtHZIj7QL2Lxzq
vOVJ2kt62yvblETdr17D6kVUhtl6Zh6RYRpYpwruH5Q9C6BYungANy+NjGH9GxbGCjzz7UJ5GS4P
qGHnKyY94h8MTUo6X58JCHMqAWuUTCeKf1N0+MQS86w+Lt9MVWcmsNTwKkYI3EgeKvDpVEaOCQN2
t9RiBvXItgr0eS4ItEWBtWfZuabZ2SN6XhOkL3G9iMAkDtnqR3jWDQb+xep0fDaD0PtSNhm0T9K+
vk5eKJpeHVk+ozu+kpGwLI6Jj/oQuIC43OMORvmMUcJsyXzEKcH3eg19riFyQdMJB4XLY5c+mQqx
iliBodwR5XWEcfLxNx71ZKKB6+RHdHh5KcibgPsW5ktE2OM57sJmy9GQw3IQhaAx6Rdo+Kg+fpOb
S8kI+H6RZcbcaMn8yMktvRsl8pYylmpEkroJnn2uyUx8FS9aCIhfnOAYjk8JBlnrll9nDVMO5z7q
YNhNA00P3+vOC7Mpvxo3SjufEvv/i8lzJHzP8PQXWxnTbhTn0F3LciOEnD/RFyCxupVeCaQHSiHu
Vx9Xe/l7bJ8CtwsArWbmNwJ7OjiCoOAAooTJ2exD0/PcuU+HWdRqVgDQKHjvYJ9+XhegglV+aTVP
1NwsQ/1Py5Vc7Qvtmr1djCbRe11HutjpbGtJbazJLAJcbLVPu0ajROvqMXhvR0iYK8AWTbkAYoCr
XajHvJBAUHLo8r/hUvqHNuzdeTXRYIj7O0Llw0ijAhv16IIOfO76M2ZMgfCyoQnkbtIbZe8qiNjY
t6QI5by0jKeRpHgb5m19f3P7+oFwxl7AURFlKU6Uqr5hYrLf9MvxwLE+5fNbs3Lq/PCCH3Q/+7RU
na+qrPU7788Ota9SmChOB5+PCAWIShrTx4CtdhsBGzQVq4Qf2M5Fg8JYFQluWgN+yDIljPXuda/v
o3jVVGm3pMMHA4LDrp+TnrgXsaCXWCR0oL8GeALJ7q07x4jUwfGlpuZ9khAMnFiAcNR4WSTG+yqh
COVt7jKDxajHFjoUXZP2TmIIx9qwS+4ID5gdM0pV+UnTSjtNOGvP1r7rjrmxhlxAXapuh95Fdhm9
4CJVJZ1VSPspwPL9A4oDhyRtr913pGnp08QvhCocpVIlHIPI4vMk/KtUVkfFxZb5LmPksV/tRWGg
qi1m1ts2ctu3p2F+xngW2mv4huAkH2j5CzHD9dBNea6lf6PlyWB3woUL7HRV8sbsroJFKWcK7PU6
tLty66cJHto9Z271L7E5+Hc+YRecRT5WqQhwE2GULXtnEuGzh0fXO0L2kRZqmODydwKpciFhHi7h
mjFFRnNimfi8DL7h71oE1E+39ZK4lMSjR+2qlnuxHbhZlQMIYwsBr8yyL7ZDCVPZvcAdRgE4cjSX
KM3z40p5jDSTTFmxxeZw5ygTbqS4+WZO3UHihZqO2o/Q5Y/euFO7IyGOud3deXX5HsLTlcH9T01f
C/IiwlxdSmAcYHudG6i7VdbLBgnpMwuCM4yP1ZKVLpJbMX+YQrlONXBft/tGPrgCssX5K+CeI4ne
OZYNtYKYOHW5bhnVPI5TpGwpgOSmevDhJz/pC2U3v+iB/GPsEdH05boHINJwOV6papFP6uwqfoq5
Zr6usEuXG52gdWQAavXlc092AzqQD+uNuRQx8yQRxEpE3DQjI6L/4qqC9HBbD/5EBoA2OLX7xxc7
sdsxFf+mrZSuijc1KbHXlu75Iw/Cska/Ebz5q1AxNzMwHq7txXhGZdF4zTt3rGOxU74qcAJRLb0y
QuINFJLKAR3LhZPkyuZh0tMdkHgVWo5ta+AOx2L94+79s2FLvT+GWfc10regPoqygwx+VFBzvftV
q/MeSp3TXJSXNkOBRJKlgPj0DBQhlG9NxmzTWA11+lgEsWlothQ/J6EhV79IBmzWCjhx+Yd+M842
W2L/Fkuh7LbaOY0jS4cBIWvExpktBOfpdxtt5prsdftVjZPuj4wOpfRaUXofaVAJibxBBSW83mEt
j4AgTSC/6XhKwX4ZLDNN/BU6DuWARBHnrgYVKDuHogNGP/LpzRIEGX88QpERLCc10IWNecD2jXuk
h5ql2XI3N2tdpdjbUFHwt5BI74D5vMSt2drcg4+Zo/hjXxzK6PgIF8FfBfMULE9EUqBtfnhKHTGL
rNzrZlX7nKKsm1e8PBeqTciVl+Z9cAhVHlwYxTjxX4eKVqHEiXuNZQqExgCyH9YC55Mzqx3oEhEO
20lQkAMvGAvskJmnosmeNHQunSiwbSitomKK2/lkbwnip2RLSJF2ojhpHKhsPcX4UDVfqO5SLGoG
654WTPuHG6YeK+lgHEWLu7G3B4bK2zYzOL4f5b609BK7mVNuhtZvdzk3zDGXLlmPyIAWGd+vPiAM
QfTJDIzoLuFv3iLBa2PMj/IF1cCWfIqf0GCLzzOz/mxQJCGsvJr5hnu/2QCEX2aub74bzd2EBLku
oqbIOwrlkxY4AwZ7E+3/xVZGEDTrpzBrRXJTJO84Fz+cu5wM8U64eYzH1/H6sJ9TvGt0akwYqQHc
PkLaQQPpa3FJSnma3WLMgGoZ8RaDPRApz87lWVMrtiTgUx2Lv/jWJo2xlH3FOxhVPZqjEm+xQz+7
2rMePT9cgcBpyYMXaVBsB5F1waqrUkaTr7CpST5saE5sKcB2yN1isgyAsqn9/jyyx83lzcsrBIcM
EBPpfDBioWc7NQf5IxuxrqKNLyqu3dgmjVHYNwpn/OFi4Nt3A131kvCbbvDZlkV+nX0ud1Yoksp8
rejLdeVGm08gVSwsQT8mzDAxo8H3l+suotI3R2zRp9iuLDORFHoAhmpyoYNWyE9cEjWWz41vk2H4
y0AKhJLpaMNQNIO0dyZbRAgDejadwNL3hMQexzL2gtEvIu6oTD3FX70Wr0SL21HEtXpl+mfgiTSi
WH1T3bCRSb0Ixws0S2o4mhNI5GmUS8dUXkhIU34Scb4rXcWa5f7lMg2ShXnHbtiWL77wJBjnIn67
YHZnlkm1B+3K8SKeUqfzpTxpzbwwDCWkOpTH2LM/IB3LB6eME302DXIidk3xLT0oadnq1pxpgNLc
mPtYMj3h1j04PiAP0KtrmFzRbwjD4EyDK1SW6aVksIeSUgJolsc+b18y4uvseAx9+ufJQ69o9O0j
MNI9/aWwebBICVFlR1lGHOaM4Ukj9oJn6t6Yx9fjBVed0bmEY9FPBOimp/tq/vyU6vyPwlSG+UDI
SIvyOGH2yBHHB5dccrrn2mCsudHglTP0DftDsYe6/HIYq0CfCoDKabmy+t556XgzhiLNHQaAhY0u
pGXLvYHH1RCd7SwkFlbEj2ht2l3/hVsfV/lmTY/W7zI7bCGzQ3Tc72wuP6G4h9xsjsxB+r5aGYqs
/JGucf9f6xHGWOsf/xkG0chZUInMGuD0xLHaN5RKlTrSEQqA+++p922UjdSTZsA2+oYhHKYMO0an
wfWLKN96/V1+ykfObu+GefezZ1Ee131slGGOWaWuQa38A7U8uaNvIm4tPK94j9Lgbf4OjPrEqt3O
zQieeo0ZZpDqsj55UuItyDfDsn5cQRsH+l4+SziOj1zxWMgFjJwoVRJsVgH/XJ7cRG4tiJPluElg
D00/TMZKEocMid0uwgPrTJOJWB4+zjKPvImCHVaPtlo8FJng1vv4FizvysHpc4oQm5cBxff/Ypdg
ukbj9BgC8hkH5J8T0k1DIFfOCcYC/lbOC/ZJe6r2ebbxD4Y2lNPZjaolOrW53KDyEfAe8osNTO10
mOwyvZIJymC5WxDRQpsvWOTJsLzhXsxJyN8soHymzheaKwngDX7qVfkUvk17rhCJGouJhum0Gt5t
8opLLMwleIX/sOz47bj1RKebF5VCXVNIh12n3pvSjivqsjoQxfBCLr+5ZVLr6JCdkq+b84NeyFrB
fl9JrK9PGRaUO9XLrhoseV6sgWuTWbcM4u+SusgYYahwdRFtcG84//BEHJDB0QLTYdW0DTJdr4cW
7nNZ9haRCpVZs43A5+mLN2uw6th+HWoVTc6/15sRzn/R4e/4jQZ/HqbvlgZh5iR7aDoGnopIOeBR
Nd0QORyXyHlQOswgTstPnAzseHRnFHnCEGO54Ope8w8b28+Ea/2ncZ0/MVgRf27GdoJidS82R/5d
u3ouaHxPOu3ZTtaDBaHQ2QR/bhMXf9Ve/zSWKOLrrOMjrCsryTMfszXgwaC1KH5JZPA0Qn2yZRfT
e8QB5LeSv/+NAEi/YFtcdO1Ko660866fd9WEzwNqD4Hy8hQXX6Gi3bTM3oYyTEHGf16DmanufPUg
UZAu1AHINmMCJHdloAJSHa15VjDmZ1M9RIIm4RczL9flCjwyz3PIYR8itvl4F43U/7yisHMLIRvV
QvLqRtozfioduXk0IxafFwjG29FMIkZ+Gv/hpz7MOGYe4NwupX4FTNyN8JCsgM8Jatz3RGhQU6kI
alrf55XC9ITCwCaqoDh68G8g5K8+NYI7FRFO4dWzBslEl9Gw2QBpJrthbuBpm4/FBC0RK8TDnZdS
RRXf+V6cCSwnMIq8lcQ5P5CGZ9M3msXqso4mDaWzpDJUtob4EQmbUucR1tg0mkMzwueXJ4JSQuId
FMAlZd4UuVTNi2FVvTVrIMxGFsjWpFio9Q9HKZy/qmJne2k64FH5e1ek0u/Qt6Wqxr9Z+40DLTt+
WpoB1rYKli84WekYGScPIGhkqIs0iWfVp01s1+AB7SEUwpTnQ3CCxDpwEJ41laNTHN9syLHJN4ly
OaGLcHtmiz5GZwAKcb7qCPMsl7dvklIWaZsxArwhhCmmX7X9Qz2ZdKKhz+auMz5aiL/21gXgC3XH
nqwbpwgEi5mVvNiTfnSHvQ1fJTSMInTRIDSEhQ9jVn6q15gNW9QOmwTm07c1QJISYNYWsDyCqhfU
RDqg4K775Kebkp9FniF2u2ebubN4Q9BhZY5QJX+hQl+mv3792Xq0PmYFIHLu24vj8ObnYtWd4kT1
5ecLVSJkKnDVhkDRLvAPblseTQXpaB950GAQeEmUCvVv1mVZJdNxk2jpN6Qhnx3O4HcYYKl9pSow
oFMbFtZED/f7/XDD+0u/rm8blHIoYAVseydY8437bneinx2JRefk/ONC6ef3T2AIXitaZGOSBP/o
aUpOAzkcHGTIRYci16RANY9TQGy8eh+oGiV/2A1ILey3LpX5iE2RunSwfaxhOCS4zXObZj86EViL
uDD8E1+fmRn1bupmzK29VDD009OrkMzWRZSfk6lP9iypQ1d7eAnECYZLJlKBhhs4u+OggdKLE3AY
AVXlJq+/zKlclObZOv69V54KQxLvrgrpL6mS2GiCxHYvSlqR0yXWpP8IIjjeR2ecj3YYlAkseGDf
Vii/ayuzJreKjLvGIs4fcs7YnfEuZeHR/jImeWk1KSTL3Kz8YHQ+kG2+g2nHqBO2Uv2Ha9IzGjS+
y8LlUwy5uN/kIrZC2hOgTdhmj2WWWpZUSmsF+KsID1cAj35cMp0Ns167hJheKWGtXByYJr9uhW0/
klcdHPqYpwQmKqNBDl2gTGCJsSxd1+Xaymnw47aM1V033rrzVC728pVhh9OVEmvxwYSVeNqF1SN1
qS3jnVcn9F5pNZKGXVYU6Oxgj0L8DyHqNFbYb2RG7p7jrQz1j7Ev51JHmpalPzPJzikCeBNugA3n
g1VLAk7+40mFpKY8P9lMOrVd1LA3GmawxYL7LCjlAaXFaeLqAGamaa77CwI+JQG+ww6a0DY+6+NP
W+6vYaenxXS3sUtP3ItuCoFEcuBUbgd4dtUAydLT30zVkWyeUJxpafCXKEUEw0zpe4hiaoYcBJS5
biTy1RtCdU+lqsij4f4d80pLu1cSC1fkUziAl8/VKUaKnQcmB46cbUjfrZJhf4e445QToV8lfAjm
HIS2o0xTFvSI7piiTgrqzYElPCA+dHrxcXEsD7LEDN317aZN2tgYUvWIXI3yApm4eZ2T8qhfhhDe
Jq9UuQO3vBi3w94jtj+DhvEH5664HQHCO8vAO66DQ+WpAoApMMfUNsx8TKD+CiyzsFXscEc+c+35
DmZOTDsHq8y2AmJgoMsh9+zRq3WbmbEptWjkl61A90DCKTkr4evl4YBKJZunVFqLMmFma0gqPCrD
4Etzngn9n/ycgNfLchlSiTURKhafoW2i4XpypxHCDCCT2Hhk0aa5FB7BWdiWM//elZqgZOEBWsVV
L2IUMmnZWoBTT3qZ/JDykAfKf5mgUE0JWhlNkJD35mcv5KPFdQdA2R+v1gXRjFVsZ83qe2iO4RgO
mxU6nI4nsxkHv0vhOV0KTOKQVHRHrhhIM2EC7d7DWkTfipfjJlYlLBXw6pJpIbIJCgwmh2jmPVDs
WWUwXnoJQHKz65Lcy6K5wnfiKcmHkIdA6AbQSotkbr14z0qyqjvMNYsvWntgv+vJq/VHesMkjLtT
fblCk8oL0mvKhWY7nAoQVteOxFPI/Luf5gC9nXa0MGl1uaKTyPvp+n95Bk1td0VJqwPEWZ/tVmgm
1BVjQfiTYgzQRdjDpI2PkffzhwkT2/RQEsVGdbDlwtXKDd1tu2OXGoVtEU+XFx25yXJavLPOhV48
glAxo4AsJxMIGeCsNJ2HHj+CHuT1MjzXD4HtLKSQQgJcw43B8uNHW2OGipV+Q7SJBHDV+Jqgd7Am
piPOyrfJSbgz239H0JtkSOfp19TfQwMpJPQ2w1XpZVi4jfPBgS92ncim3t8t0km2l7u3T952dsBd
J99Qd4JjmRarPAIGiJ7QF4YNj47EyqeBlTQoVQoChhst8py+Z6c6cCgjdIQHDh4bLQfnt623robz
04xtlcy9sQMYG6l00PoZe4VXkReCrZo4zHz2f7OLuBR/26ZO+zxi6dXb5Iv9Cx9CxAw64hgSsdid
7zs5K2IZGLexjJ4nnJ209q9FuvRQV2MIx4xR8tTbbHaTyajCs74HDHvp7wtSdrQaXJGbUsm8f85u
r05SPoWZcinmOyy7JmZeMZqIbTSx/bAFn7oFPNRT/y91if1ajB2tNw0bdYYwTcVaQKNSHgTKpUrU
iR101xyAVKndEI7qasMOq5t5X/IYu1y0vKtmj/70zezjTzGXOIh5Nw6b/XfNFVDVldT9RLzvnvKP
H7rbPnDTu6qRi3HH0XD2DboxSVZo92YlAZ/B12kqupZ1VhUkYzmHY1Sw+EZcWuD3tueDTD/ajfD8
mkMpegNSy3xcBf9NjXdJ3N4DPQlmVXtbow/WxgR1Ry9KUd0N8UZrV0dCzfGWTqta0o+72JydZMEh
5S57rWZGhIsVYdRXq0WWhPEdWHlpTsC11jmFHeLnC2AEqkIF1PrHebOMT9YoI2jS/pepFXhfs1Wp
nDGxCsFn/D9+1I6ZNzqoyjgOSgah6Khk4yK70U/4zJmcy8SZQc9ecWxEWEnOQR0LfiRcshdqHfkH
y/onKenG/t4tgmmk2uTFiwyoZa+3z/7DW0r2Gnr3jetPKT/w1s4ZVVbzasjKxskOVwtypRXesZy3
4vJ8GYUOU5ZoXTqfrU7jV8DfwdyiYdHjNF5aYa5ZMz8rrmWy+DxuoUyZzP4ZwqXQmCALEdTnzToc
r22PaGt8XvZMjsUyDT5Bzibjrrb8Tgr+DB3M6PMLQbs15jO9GdPTQxCR2An+11tC0CSMwHoPcTyC
YoiFcZm/8XED2xH2Qz6/5g5QcqU6DUkDv+rvptJEfQ4c+MCOaM04Kh+yXI6vkOTM8232fNo70j88
e0zfYmmgQyBLXDEKcUP3avtTWZYi09bcW7phIhioMN+y9JqLdfu7fMMoMOphaz4aQ0g7EWu9sFYY
BOQGTBVtB++RK2WJIA2HfY7TOInKYv+3clhpjuEUMUAL9qklQDUT1yh4oaBMyrOFSI4EtQfk/ITW
Kbjq1WQSDiC4f21Zt+cRF0BhVukq71NwzO3BfFIWialmdW9u4QrVV+P49xiEG9CVksv2wyHEsRnM
ylC1hYUTmr+AAO3Ov5i45JV0IV8UXthM5+2vTZzWmpTNESn2uLK9kzOB9uR9gTOGlx6APcTMIsyJ
sXuVlkYHcNYzhd1okF3L3z1/hQBeNzOKUNy4sExBWT5cIl1swoU2WFF+WtOIBzFM4mRebGlqeNI/
YHUsmpp3HqiSLmf7zxBmumInqmmWimEFSXI61mdBGvCLz6nGHw6k7g+FpQiQW4rvdi5ORVmqZ/xs
FzOYpyynUODOYQvQg4qvl2QYEYqmpIwHKAaNTONA+DYVXr1KPpnNGYb3kNLupZEOis53SVDe3uDe
u6JyOv6EGcNI1C2B+VRH0n7qjmBDVNAAgn2nddn9J5aDWM2SGEFgsUKH0J4iHUbq83yrUE1I2emX
owlVH0ntjTM9zjKGPpNo2GzCANoN60p03j85wZcZuJJmC9PnJO8TxbrNM+aSxgG+HdRrLimBLbfS
tFdoJNAImWrWSCmrcqVq38p2DYc4FiF9DE+MISv0gR4c/Y+mo8HmyjSfCfY2OIzCNvNt2M54VL6H
D9SV4f2AWtqkoZl6FMzLFZCG0dL2BW9odVyEWnJQ0Lyij23EdoBzMVWfPYCjD2lwnSUlLc8qAWHt
RB4UfnEQhv/kMR4mnDkZDniCOjsRm3O6VI/WVGWv1A74FjuZku3Li7nlkZAiT+qg/EWX1YG6iiFz
Vk6swNPRXnFr6AMBxA/iqvh8nCE2Zqf16e9F0EY0HFU8LELRZ1N/OCoHDb4tGMGL2+tGoGQFDbfs
MfMNua3z66XWyU/2FelsdPAAMVXWPG17DHAcrUwaCNNPR7u8o2Na4QBoPToJxGJxzSzC2v5JgCE5
LGlJ2oLqFU3J2gOf7Svv28dSAFnaeG7+nytVMuD0QnmUuUWqhs9szfbJRfttYH1YhKp9/zTTR3zH
6tshmbia5oRaAALbRC4hHvw7BsPiGLkYihB9CBiKIxrFXpmxaVoZX5m/iupp6BYYOu0Iy+9iHli7
nPyOPyNbcUP4nA4If1lDRQdcDaWNsscIvZeoAZVGANwsEQ0Chev/DJemYtCzofuzn+aEll66U/uw
Om4zHRLQF4PX91GxW6zng5ZXhzR9UKiJAs0DfIA4JeV/qT9CRCaBsSTMlfngkPJawGxp3C8VeL2I
xl4m/PgrZdKs0liSj6paI6nTPgDw+own4CY3dsdCc1JXiDCuEq+14oOKROSjfSdBGS+ae9jMXzaV
5ThJKFjOEmsRuoG+S3M0i3qKK1xOvt0ZQtCLSU8g/o2SI2EX6LA+6K3iDUlk8yxQSt8cbdlDG5BS
R4aMt3QE75HrbY3dpPPJxMFTMCk2jOLKaL6VwHLRkwRjX/zYBLhpV5KeVAl7Ce/OKPmoM5krWQzc
rDlnVm1Dv3fGYIZsIwgahwEbIXo9W/pm7UuijS1niSGR9mRCxgCDrfNakRnM/q33/pdaRlsZuxrb
jS0d1UMq7FSeKdoG4LoOx8cPtRdStU0EVnVy/YOI3XO6EGQ9CV+B2tP6+Fcjh29G6a6fqrh+4KZP
62/8QxdscLWp6Ffj6tqZGjIuLu0PPTo2ATTejp7ak1rxjPvvRilEViQ8Hqxg3oSprVqjbaXFP1gf
FmOAMDYeYv5/rL2ZAT9E+V2/QXtlsPcsgWM0ngcQ53WF32zcH4v2iAKA4RcUYtNEkHlt1GOL80m+
co4a1i7sQOMCYFeetwlxjgdOyAFwjrefPUAWw1DQZW1cnOiROeGxmIuBV2EEyBlkKlN6RrOvUJG7
VMWlA/KPIJX2Urrc8VS7Mh24qVixOleTm4QKI3ssBXiWQx5zfFElQsq4fchiyFpIlCHtn/XjorD3
d9eYOStWJt4UD2xxFIXJIcUU4Y2XOXFzp28p39O1k1CPtOFU6PA4jzqJL6zk2Elt/EFc6B6DP56J
XKi5UTLCEiamxWyhz0dHGN5nAG/j4Y3Oxl7iWAByuGuxFtVE9d/WluE8tjcECsd0g93MuUDWB8EP
8kqDxb3L+voqJsVcEgQrjDsgbhJfpf9heED3s6XWhZfVX1zLBfKj31dOXu56EKVni/H6Z2AyzxdC
80LPthwMZmGvozsR6o+PFPpUSHgOSE0EKVgW8OKzehP1raxNjlophmOLZipZiCh2LSau8kcPaQaa
Sr40FovZkh6+ALyhTT89f3MkffknrNBOXTev9civmJE4qNHG/aNWe8guPlsyZiHe1/xEWW/aInEk
UBI4vInZjXQvZ2KD+yWYNhnLE3jIdYwBOv6UZubdmwLgYBP9And2Pg8ya14CdnQZeUTEHL45MmFR
6jaUmS6Ab6ZiwRi3P5hZ5PvxP4a7IfeeLhZ05O1+rKIaNq06bVhnnNywlpVmbv2g0VIV89drqdT+
2LZ0CBqwpTmamtwehq0KYR8jRnHfF5HwYdODBAc3XQWPWqSiY3b2zPU+NkANI7FUn65xbjE7dA2y
WmC29G+ZCP4A3yMR/4FkC9waXQlPmDSDEHIB+vwL0/NXtsYLn/t5Yz+Q/tveLVbxNLEwtMX6fTFP
Dm4oh/lviFLf1SaiFFF7X1cj3PS0qfMkxVVQ8d7CmbZiEgiG8M/fnutc7D3HXS3IXCy3vUJzjlPI
dnqAe3WtjScrWI55hNpJkD30LyMSZsqrnP8LmZb85X5GyzhSmxBaMfcQnbUZcy9f29heVvGhREVt
yUVg8Ulk1h7oio7Rw2nQOoKq3tJcJb0YMx9RdTo2pOj2Db6O1qXHcYfDLY1pToMlVzLTfcdXa0kC
30M21TODYmtSsCJ6HNPp+9t6msBLPO1W729P9qTQDuH1yGIwMY4AzYAqV/u8DF7ES7lyZHUKsmbK
ChlGvaNo0870IecVNQXPxezKEfZKULtjClZUBestQvyxGtifx4O4jt9MhNp2a/V4bkFCdMvhKumK
xJmZM62ugGMBj+ICvAD5KlqKY7bLSp2inHprEWMVNbnOQll3vACSQS+C+3nJwhUINGdNc+LSoq1C
1Fx2Lw/+xeWOMn+N1m9nZDboxPRhTD22YPkFtUS0Pkfe7HdbzzWoA4/PogIO//nCwviMsDHjmam2
CYjvl7hGyaUdZbke3MlKJnManKQPUtz433vmlnYCzkDmvD5tJM4OMYXW5ixxBSsHe0SjO9VvNpSZ
YEYNR6k+Jf3cpm/GufN/Mg/oOJm/JPuVgN5R5I3laPkCXCRWOKytao5WOkmYFHYmN0iRxCOIcYtO
9s/Bi7Apgc8RnS46jEIwfYScOedAEWiRcPUAYKq64Hnzl7G8EBXmPKV6ydZCI9OWV4exc0vpaB7r
VLIRxUZRixspJif+ytjxorB5yVq5mJZSSgEnoDRwcnT3rP/LjT0wZigiBePRYXI8HZHfk32IWXti
6YYSSlLeYAOah8+gaBs+auaHWVH8rUAHcM8jGzlyQl8ViSrVjajJ1sLx573Ztr+y33+7Mcn3l0fk
6/BlFbEyAzqZWbp/1x7hD6ESkqyfdaDj9KPbyUc203LjjXU8LYlslshPGYnZRadzJQDwtSfDZPIf
vLVhnqXxMFSrZ2xGymCj5OOGlGkZCLeH+yXT5eK6MtgPkfBGBj/Y2ezz22k63QkFc71ylOId5SOw
3xR6VO5zA0l7MMH51JeVToKKqphZjS/rSL62vsUSBVR21eUnMeTbgeeYFPepaDBZdSwhYImLKWwO
adRdZV7nq7Qt2x2GdFkdjlerwq9sNRkTkgqS08WuC/HAX9nUYSqNdhVSHRBjjqbiwya0WOSHn6Al
AL3mkn55uWmA+oPHfnfTiJ2DtL5cpgftcxJzlvgRqayTkl35ORgeuVMxl18pgqtKsO9Af8gVwHGp
zfGiG4NIkd/HtRmIXq00BNpEpXqx0zAWCm2shi0dzCrCpbGKGC+JYSZCquMD4UmKpzgHn3W8cJBQ
LhmRqpWEcfuHfWFN8lCB/3ujwYhhQsbXUAjGjAMS1/ghb8QH9pkl7lhbIsOox78fRLW6glZ1S3gD
b9Cwdq7Uu8LnfiZXpoaGONfmKcdresJ2zmh6OEMzO7wHZ1WvXH7OD/a0qDHBJJdUT5NqJDybb6Zv
MEZ5PDSlHa3qfPsHjsJvB/+h53jjLiYXY1ftBjUeS4V9AuVDAopXmM8TO1/H+V/wz91N2XzTan7K
5G3zWkdtctDwY5l2WVKqkRGZpvyd2A98dsgR++Q8LPCahGfpy3oZZRQBA6zTWTFYDgX3+DG6ycwT
N+yxywWu/x4CO5qRauLEsWWcatVGV3acOy1FOXh4F6IBnO29FVve280Gm/WRG59XS6TTqIstZ1zv
IykVQNHUb1SwG3+cgGxDhdH6j6AUOS771gORYJvVmt79bczVFU51dIholDl7ac4Wis+3HRufDDal
t/6w0jiWSV9hf5g8TNt9tfLiTtrQeAPKbZ5Pz2o6RAIZAtDvJGWMjDRNOr+515HmtDzdOYeul0Ga
/cspHX7lmTfiam1HpT3JzPrHuhVkePsK90TzFg+EVKT+F3wHKFH51r8edtvbWTwPNtt7gtMhUOnO
78d/pNvw70JUwXhoYGdt3grJgsZ1f9bCtT0SiUGYjLZUJBd/gYmQoxbZPbFVYaEzaGvb7y/mP9Py
A76mVzbUdAEk5+MtpY0Xc4WLaoROaG4AvaFV989FIgrQjACXt4h8Da4fhZhTWjC4/5OB5JqOXgTV
+AaB+DxvIgYqyyzBQedc0rw20brljBzmYxZn+jZlM8TZden6QGWdwH2IOW+FQOc2hb3E9MHGXvgs
gedRaxoGeH34jNl7HBUuUL2QU4K8BFI9olOSo0c4lUXFWbzPBqCodJG9PQ5IOdVvdqnW9ipH9YOH
ocyIhsCf2Q6lcXQmX4qhbfU3C6xPv4vKm8v5Lf0JnsZrQENfasttin8Af2XLet7yTp+d4rQvC1RU
SctoMN9XRHdGTWTFIvbn6PUEFGss3Wn7raG3/xEP59uywGG+j/SOK0Bb3wLT6i/Z8zN4M+mfrfBl
lXDTF3P1yq3gWmkDGpMBmGb87DU/WvyZr/WjcdGqakZPQOJbIR4N0jv03FqkCGdukdt+HbR9SO/8
aOaFRbe4g+3mB8xOuknqHa2qagHJmlZJjswgN3O+NfZS7c4l3LwqKycWF9Y5bEFnhW5O136Pqqdw
Vm+bIcoFeZsVE99FRsWZz1M/sJIDY0iS8H2jxCUKvyFHJtgMz1sNC6WQL7ROJ2UIt9PnHt5YFY4E
gfXF/Tnaum3fAzkhVHwFm/mHdOni1oviuNky1VLRBJ20B4GUrVuW6oTPe2OjldE98v0bbILN2xCK
B/aLF/7FrDnQFnu+0BH3w0+NncKM1xxwmcqfhkuw/iYYVYLLqSWzuOstHA28UK+iJ/HrV/NUrAPL
zRX56ja5aE5BQktupd7KxUDvh3FQR09NS9dN4kHf9PV4fDw/siVVmYsgxDdGtHqla8iD+L55Ck7O
sgyo6ISkA+WDuWFVd4VwABVTJk1MSaa2c9/eCN4Q2yoXwgogpdxFZqbI3zFwcwHVl8AriROl0AY/
Y4rQSHqSFlG2Uve+0/8YD45YbL0Cod13lLszb3wY0Hl7H3KDM+jnsVmQHtwO6vBNRqGgaI9ULUUC
V4owI+a0VW+5CO+/+TQFX6AiJCIVTkoFHiknc39tvEXvOdGjfZyqwk0BI84s2/WB3VY0jkLzGmqK
yWCPvdfzPYokLudIXqSHo8TXDhKrxmMsD2by7SC1PBZDwQA4evgXd17z4UVSAzFYuLz0xErDTpk6
NJKfZLLGDMr3jWqvD/EH0Q3JP8QxzEOa3KJOBshv/J4dsq5fzLMnO8t6BTin0MW6U+6kKCT2t37z
lqoiftVuUc2bHj+hym/E1T+Z+YXQv8vpMFnMeLVj/K9hno5ImIf8koOqm0d+uoH2ZZpkobVl3DDi
I6HwxOxnR6MKbww7Md8tF1Kgo52kGhKxLghfN5F61hmcmpwB4nl9eKNe47mDAxL1thPTfjFwl1y6
vwOxHBqsOaeYSBRLmPvL4200ASTnP9D/5zSLmQzdOZabwcmYPJagWWEGT1It3s+lDo+JDOV8Tcre
CsULTGmOgLGtj0uk9i93TmqQAeLk+bePiG5EsyYFR2E80ApuBImodmvH5ktZGIl0DpviVXLZqtj8
ppG6IiL0Z2sI9snzqdBsdviLsUuBP3dFQ0qQDafyFi57War2JBtYw/+fP3sAWIQX2zXek42xuewi
bfKlAJQI7Q9hKCN7eiqJuOhV+QgjF8aobhn5xW0bybXrlLRoBWqUnvSj+FM3C8S6Xx3i/0cPNWo+
n+C7I2vd3HVpkvThUtJwCM8IvXBpCshyOHYEXxnG1QUVKwaztwwcjs9K7LmKOaO83VCqp3jYenF5
6G+R1RFfb6CetRagpWC6Pb5yTqq1sPlmRwOkiRe8I0sQor9ykBmDEEhpJ3M3PskNUh9C9EZM1Jlq
jRV5Yg/bsKcZHiPbJAR8GYf0SNq5s9QcNhLZORdn9myhphhVIEypMxGc2pGvgi8aqSgVcrlPehmZ
8VjcZQsR9B2PC6WleiQSYVF5yxZQTgoML9UMguGQ0dSXdFMBcktBeymKr7lmoXifKIfSKUUb9lDM
VlUNg0wwbqF5HWyeofOzAFV5BgXOafN6I79ffsj4ePqRJDkQrxPq4S2nR4A1oC+3K6T8K7dD81XS
+xhtfTpwixH3ki0jQ1K/AyJhGBy4f4dMzfrrShHCgfy93C6t7fDjzRnylQPWuUR4a/U7DFyLmozN
amVp1RBXXO3AJ/YfYRvoeC9TGibc2OZaQIGUWst7IOOCpTtmvIMyp6HbZpmCTDf2iNjPMUwwOARb
Zxva/sckcvrAxylhwnX0LHxVy8p19mkDeu04xw/BRfukvfLybyLcOg5N1xC2Zn2UDYdCyP159FEg
QkQXX+zuOwdVepUvPb3PjnauUT4H85X0nzVv4kTuquD2eF1IzCjzBhlhbCZXe33JV01GHY1wqDqm
CAf6K4ygzUQNfYAE9AvobckBjFyFAk3VWbleyFO5+4gBdYXnBBrrKHmW/ZPqT8keqL5sPwbCAvkR
WDFdhIHdTfd0dFJaEbeD0Lqs0GgpeYrRnwa2awsFGkD8l4FENf+eQzHVNNvKMUEixjnQP9BdMCti
8n/ornUvCp/5JT0+o4a44xOiHk/eR95Y+w95OFb98s+qY0JdSFdZ0A9DXBQ0yG7gcenL24xjO9CC
PqkGVuqQ9PsjNywrlNkjmqbhP09QTeONFj7OazCf+CcN3E5m+wiTV0/zOOd0zWQWDkfr9zTDf1B4
mwF7YWecR4cuEWbw1+CSeIKxH2A0zbKwgRWq+X4aaeO6PgBH+BJ2E+Wn3V2GtFZtHck0WD4dGzpi
BzEpxeCd8tFKY89gqCKuNAkzRN54NqjI7xwsKkwCLySOd0/npy/1HY8Cx6oGw0yEhzZulejQxzNk
6fqZTZqk8DtxaZcCFqQPOB2a5wGXZIDBuEKUA1Fb7xLXWW0hZhK0jbKQC/5Vas3NFZJWnIq9Yz8x
2DYDYo9O5w+rxPTVFKOdWWg4OvHBxklQF80lNENfuxX7oOinfUUFA7X5G/67+J+INtRouNIKuhjF
l78EMZclrXyBHCU2mnydbBj72BaxuhUS1S80Bz/CZNvpK9aMA2/5XHDBxsVGp1vmkffCVKPsT87V
W7A185gRVpzNI1C/HkwRWieTajVvTGz9zlCrLVOBTRE53kpRMAr/vaq1UdM3H5Idgay5eEtrqKIg
1sgGCJzNatDfagR8oDDVjKxPHyTuzry0wAMuCnJRbuTAAoHhIIEZp+zd9l7Zzrwxscu4H+Ju7cet
lODzZZXWN+Qlvi/l3C5pxekFsD6pVh5oNtLs6XUELwO9Nbu6hcwoHgChIG9SkTkPvHtTI4XrNBS1
cdy67afxPwhe4rSHQB22clcQeJM/jz5CVP4yfOjlmjsL8+kS93m/K2VQNLpm7AHSBLqAdKhGF0Y2
uP37Kx6zbYMKSUKGBU3TJKehUVUdCoR4MX5o1vQ/k2Ao0BLhASIxwkS0ehDRx+NslU7YAdF/TXXV
x/VynLaXKiVMpKbZwOz1KkNSXpTC/rqH5y8qsEH5/l3cGQ1wWbtIyr7lgSYWOCOKzDhqpFl7cuK2
geCxB5W02Fk2neuBnM4RjQ9lqcyrPBxeLnt1muAukZiL8fYIG1Gs0H0RGgnD/sd6OiUxsYk6Y8Y7
P4jhRccGTCzaTTP60OjYB4AOTwLTCtoxnXrlPbaqULMaEdqryDqxvrYVU8a5z0kwtiAwznVUp/BM
0//E/LaTaIXEvlciWyyuM/LLgkooqpPkRs0gSXH9fAhT+KuUNfcI31KVpA2WiEL26oxGTNARlf6g
FIBTPWUpxkPxExaGzssT7BvV/HJIVyLhfx1ukXUj4vi30SAZ/TC1UYwuZJEr+1cwZTX/n77Qjk3p
ugM0K9ClWHKCWI6Cvl7dSD0oHs8ycq5LCETNAgqx6tLmfji/UQhjQ+5A8pu4T/qpAIHzRVp2nYY1
/vpSAaoLtHMIDjc86vSGCm1CH3PFIs0CGzawAGjnz48KcD5YVX1Cv0fcd4aDeWiBbJUdZ6lTCymU
mDpEdvdqzzxnOB8rFB4coLzBne92ih9YZ6RZdsgg6sE3AP/k8Hto1Y2d1XhSqQU2Yr1iBWe2poUW
gS8GAkvY6Wii64/zJ66PkqiYGD78NhU0MezHv0Dlef0Fj+Gafn9ssUNlXr77KnjUqe8AHgJaArCP
tL1Z/SJxY6A7Bf64TS8b5GVmDQYhovcGRbpHPPNYHdbvY08rNG/a/gL1DdMfmP0n23wyKAeszPfF
C4PFdij8lsmNVm2DMKTrfligN0moRfAYysN/lFOMJ9UkVjn+x46rmUxgx7U0pHQu056GLXKjvdw7
7yMmMkzY3cL3WT4NulqTE9l5FgIfq2jUhqnX9TfyAXl6wftmpO4QxO7a29cU478ShHkQIYXSYiny
BlZy7VTY4pQSSf7V5xDwm1koWY+1BbF9X3y1d8Kq7+vfmg8QzXbdAMDE5JTnERkmgCyZhKaDCNvs
iDIZgV8UPg3e9SK7RBDFSwH0PtxqMT2nRq/B3VFX/Rnsje7O4zBvegrDo8llDljN9pmc4tJwFPfd
w50cZC2MGtdSHmx5Wq+sZUZ/o5GUVX3jhtfTHOgRo21m5XA1TZ4EEH4AGVsZmczJe8fDXuRfrxEF
MCzopjHR1YnT5WgUzIeyabfAFL6Jcx7duJSmgI/1K60APzqxL5s95Rco8KXASbrvMrJSN8NJ4Bvt
x6gzBdM7uvO93n89XCjQg1gx5kqF3H+X6OPcEaszLWSr1rh/U+Ju6Cng8e0cfYZkWAhoTsefSfWx
J/gkAGE5GxPugdE7Y0A1vd8qAuuOPhi+LdloIRewYb/KaRR0SfglXjNFQidp/xqeK/w1k4CjfU6o
Ux040R7gpJv1n3zOGupoxVovIesNPJb6fgDFyeK2Ob1Dx4gt2vqUcQom3SRgFcwcnd1gzo7C1CLW
5tH8Uei0nIBDvU8ejKhDfuK5Q1Tm45Tcve7McBlmx8n1oR1r1Ar+SgeiSUH4N7/L+SZDRnfLVJva
oik1M09u1KmPchi/UWn7m45d/OkEbJC5rRer8SoXlIEzftM5VnCqfyCrJCy3lpOZLvSAOIuZWAD/
P3sCHh6U0QV8pmRT4HpJT/KuzBwSV1ScJO9fPAj4/6lCVKnGH7QKdoUjr8/AWRP8jmTNmUBd3hrY
7E/0I0yAineFEecql93obFC7JgD845x42sn8/C/U65fql5B4zEBZUWr3yILTcwPLL8l8aXikqoJo
TKFzk6/QisQ45VfTujaxtMWNaC1/2SGbu9kSuNP1vzhDB3FyuTX2fG0qLUYHIrJbba8je6AWvwK1
W9s72a4qsWdFMripxIQjiwhD8oBfwR1hHSQWxE8tELgLWefcuYK+A5fQLvqz9C8SEzHZ+DQEo80o
LLq/1s1RnblLLIVLduvVqB1quWYXSWzLOtgT/Gcx1O4SkgMUUfaBZZYY7NclRJvBqdT/m2QWsorY
pxMucgrJJar36G3xV6GKUmOFolxPk7vSWU4ZqT6SgBvF2QC19mCUawdk6xCjHnqTGCOLuFKqcgYs
IUF6iP4F3SEI006VQDCX1VqNX9CM+SgZcKCEBCI3Zqz1x9VO1zdRPwDDn/htGB8TBeczmAewlJOU
H4SvVZT3GzXa/bdtsPv8Edrqh2XZz+7s/j6DP4oax+sxXi88cYMvoXKa5+oHudkuKv7pL2dQHMrn
dGCS3YO1Mlu0hP3oeoUxuQum0e9LXmejCayF9hwBjwHTaikUi3pN1B56oWxn1mGjKhUz+gyOHiqd
u0OB/ctTV8mvTb0Gb1H2YT4JXo6NIJybTkZXzHmeJkTI50nizngBF6aEF1icewg/Wjlb4AgsoRCj
Yh016Wy+prtuGvjeT3VDcNpHUvJzvTsZrxwKYdBrVr1fjaSMjUvs78lUBr6Mtu6K1GuW1aiw+ZsE
YSQ35Vs454SlmE9cYMH1W1LulSuDiglZG2/j2yJw6ksC5UTymW2RxRMj5sMQIcP42Zk01V42u3I1
enr9N7goYzL8Sn4m2kFP5VdRDcIscWyiqhdkPDwyaJlsJyJroz2KTKUcdI9ecbPauDQcTi1JqUQd
VriggkooRBelIMD14niO9bm9iMWko0slZ3GtDaDJJYhq2BbNSDXJJGp9sHghk3mbDgs251uS9k2C
DLX+mr5PyQHvtFET4c8m2PBW4TK8aYkG3eujuJbRM0wpIFYjfswg8ox2G51Y/2tCmppWDFFv1ElL
Hzgc/YmJnSmNf9gw7goZuMmtGiEiYcB9rZSqKCfXrQXjmoQB6WU0eSc21Q730OA1SSin2D9hvjvn
usIsMuDZYkdH8vNfw7aJBR69x92blr7rbCun0/hPhJJKdtRzfDENklhFZRRxIBSIWXjvxikfyZ4a
vfl3rrIVJiHSqBWRwSKhYe96CiP+LKwtCaI7fV5owf9Zigp70lHZZIXCO+x/QVosubqJJS9Dl7E+
T5p/JoSvnbJQ8P7K6/Ev2f/NKta3UXu1wrLHaRX2+Bj9/mecx0ufdfLhIAp+Chkl56rhqboPrrAw
Gtt9TmYX2k86xNCgeamjdxgVn+xFoSS6ylRljohtwu4TGFrhl8Pjzxmd4QVObTmgREMp7L4PZELL
g9CH3j8aStf235U4NQr2droVWqLLX0k5RvS+C3B3ZLT0orXSfb5LkoKsGv+/GFOt6hAJ3MIC5fIe
1qeq3i5nyUhyPV9eCsNaY/aBIpWHKil7i3nhvpHHgmCNVggndghPEraa4+jhUa7zWNdK+eeLytuQ
iMkn8LNXCtxT7G3S9HOlbjWa/seZRCz7Z4W6ioZ/G4RiLdbGG9DusNFxXcOVDjxxmxwqH+E901rv
/d40E9afY40PXF6eGNydCcCKlrh48+TY4+rft6fMA25Ze/5UnRtUSpjizMtncqPTQoeyjEvKC/vv
hLU1zkgGJwoqYHUO740muvYC20V2iP6uB0I1jRjN7zkzv8e4jlI1J/Um5WbSvx5BtQvCW7xd+rYb
pMMG7Uc+twhtBuHZT/4nCq2Ft5F7qSnGbMg7DoGQvG+dojyC1QZRUcJssZQ7MsaEFQaQG124tBbs
10DGeGxIPE+XCrw/MbflDPKAzrfoj4umn28YL9h+PxEG5Jok2o3c6bs657PUn8qUKlAG9GvUbs+N
UU9WBeRT0l32Hvb7ncw3RPmuN0/u+IG1JZmFFJ/Cusbluf4FmkQ/g8r9d24l7MO4hQbnA4ZaC6Nv
q192zRr0meFaOCj+DuU0o/rhUijRriqm3vY3xWRKC9LB05QtVJqKzRLkxqpXBDfym6RP+ZnJyuFY
GBtBt+VoI3C8W6TrgAnWE2PnMD0FeqpTuIYDyse+wDzoAk6xbFdks0PtPpT2F4tC8wfs/2yxJVcB
qSrrbSZIcQZ3oHDSAhlLtoB4mM7bR2Y9uV62Gq90u4bP12EWkGusgfUpJgB+a3CBoLzHzMY2+DBJ
y3pTRwod8ub6RrNzfOSkvMYh2YUXo9tcPbKbVG5kGELHMW70CA2oUwJsTNPxEYGcZZ10xFoVuqd4
lKtQilbgOK58cTTYK22MuJsncjAUt3I1AOWf6VmYmCExluo4OquTrlOwXgT6IFzsM05Jjihhi6iI
kOJ1YF4S7BwEmOtTbQQtn4AJia9YjjOUmihOMgpvya35YaWw/13g0T+b7nvbplosUbxCueeIfX9k
kejXqT90cuApT6TS9/XiB9wzDJeh8WO5b2bQ7SBAmvvG+NII8EfS9As+sCf5eoGiks3LAsTmLVPq
vVprFs9xFAZY0rGBdtdR4P9cprO35pDikFcKUSvhYNBMcWuX25+zOAoFCmZSSKmc8s1E5EUWRAfJ
FQcuvWHitIyLuoXhD7WpfjgcPdD1YoNINnC95t7ydJ3vxP7kax+dz0DhxoxgUVl0GpfJ9XDIB6n+
+0d5Yrhqs347cF02t2ZxBjSoiwHU1fErEl1hIxXXpHKMHY+zVtMYM2og1QdZZyfKkOIvDuTPQcFh
k2wYGgADfVecsxF1Mp/K/8TLUGzIUanwkvasry0Ehz4Gr91XkpajYxR9GJhBZhOCdp5x5jyO206a
7y3q0efmakEOLeKFtW+Y994KrVxHnPmEaddv0YgmGpKUyxorQh1RZ8WSJGRVKgqx/qUk3U7AISCp
05lHtUmewIBWyPwCbWTcbxq3C9Rm33BH2zE5u43aOVyTPxdz7fAB7PClhVW9pzrNws8wboQt79sd
wCRC7WWh1z8gfIx+AaceGseoOOzhphWRx2qRTV8A/R0uxJMjIUnMcOiFSV/1lE1cxHq3//q7DQvF
jAenpzydGs3W9w575X42LD5t1X3HRTiD9Gxq0a+Cv8yaILBezOKxUoniqEZEIVMpgqfHmnwAojP7
pXLAsDkQUXXYV5RZIhfClvbnMBVmkpLcL6BLbQL/LLkhBJ0IrXHJDwfotG6skP0Zvs2Kqnmsuk8Z
ASBj15CDb0da3s2swAI7Lnkn9VS8RRs7LuYEQW9qzvSPt9ZINMQMpu3VExcGuybFS+l+7XUOq+uu
4RDp5MZgn33iSuI7wcnRVFL431mIUgqzCY82J/j3wJXvY+VNPJwEg2NjDXabF1AJRQfAAUAZtafO
nv0+sdyuBR8gEaC4+zPV291J7pCqPWC9gvOPCTvzrPUUAe4eIQDwwm5d3GzESRMgDhUBPc9EMC3W
QDBubLBcGeSEcbDBIclZcMS0qIgceGNg0by1NTvI2DQO+bQayribNMuCCX8G0mVUrzaGimw/+xxf
QNXrnKIzU7VGff1nQIFOZW+wTRHoXOGRinHkkbbA7cqOiDX+yO7R5J/xuQutLDVSeFJP21A/LOMS
V8XFrTTpsJ5/AinmDHRJ1U9S7gXl/Um/EmXpxRfjWLyPbXh+RJ8nuMQZA/sGROevWbRIgeQmxYiJ
drXEwh9lnk4hMkJlZPCKl55GNbpynCB39FI3rG4d1DYrG/b6JxVPco8WJvFF0Y9v0fa//eDmkUSy
Uog2pAY15ICoDzXgRZ/DcdOXXkHyW29xv+V+t+iiL9lII5hiMRGWVGvi39cHAWpUHvaK5npPBv9J
Gne4250kLcdkvloXu5VeABloG8ANPzA9DPUw+Qv5bBfy85hTPfloUtiKJMW0TvLZXTjFP8mqB7lp
lUUQirNd3b79/8CsqYVBu5yOQPG051iAR9HaFubwgXHI2t7iU2CObeqPEvXNei0g+Chrz+eOi9Rg
+aS7DJDZfinVucdAHdZrGJZDMWFWt8oK2kJRrGHsf7iVa4HKmu/MSVuCi8k3M2FucZq/CLfz2cYd
7Xl5NEVZLsQsgQJ+nv+QnmfPFxociH9+F9QwNSPVsPBHIYAj8YETRIYNRs3mU36snrcvgKTdsIE7
qDsW7zhsxfY2PbGyoL31sEM2ss4MwpD0VcfRX1VNFmX62bV7SknmW5xFZSRm0N/m241M1daTGJnu
GrO3WSqICZWNjfyqho8T9RUFiighNKcV/oCxDkH8NNgPpJ0MgDF8+9JNHMr4nnEIVapaa9o376HX
yq9CYynX9JChXPINeawy1Pn0RzL7Al8nwFA2FarkjFjRJdyKuZWBFimlnzVMCDFZsot8OUnKodZT
CBGz7X+1fiiARTMpU53RIpAXT2rCq4m7yBUO3LS1fgFLss++sbVr9SakDQ7kNmEwZK0RYH6GkHzK
0bh2zuS/0TIyEzD0sJcNjq9vMT0s+IVSPUxlDyOGd2zjeEgsMl7Nrw5oK4oxDostm3Hmib99RV+h
/9LltVxbGcSmwlfrlM8d7Q3Tj40g6vvh/ixkR5UedkbULO8ISaK/aHY+BG/tgeerNZRR9qRdERvH
CcF1L6iHSyLNzYaFqoYHIKEJu+gxjvXHQtcDxLrQnXXHWdzjtg1mrC68eeZznZ9pAI10XDnrp7D7
kNtOekZn5EfWmJAFtQxNpbZvn8VgLiEj+SgNxTfm2QXUydkFPfL/F6MgIwJzOt6KimsPv5Tzrpru
5nRRUWgcq342NS9XdCcSASAHw0+neGZYB4Zj+rnyB/ZLJXW5C58kfFau0XyYuMiqleLPEU52F0JX
06TYQDuGH0c8Sd/pVSzzZ9RUHhe5PVCW98whQmHGfjiSWkPInWGDMD31Tua3vuPU98gF91XSjWeb
Jt5cFjUdIA4Zsz9mW01JorcFxtm84kp3AHDSZiq8E9ZQshQ4NlAXoVzt/atyKNOYzqWieXt5qRr2
zrFqnpqp9aXnRzRpt7oKxbywakAJcCdk/6yEkkiexxI8duhxr97yINb6ox2yCfOuGDcPrBG0Fg1C
RVOshLjIvbRpzTFCIR1SU+sAViSIrsOHGhlwtHjOLtkaN4/hUk63ZPz7dQGTWsbPRfESaD2zUCVV
4romjbMCZFEyTIOvvtnmjL53aHXZWM5lc11MriiSqdeqX65XgiDkuzMoUnf2/b252LRHwFY0HQwx
W/crYOuPwedfsVV4M7pro+iqcN8ZHV+2SF6ouWVukfoo+TOwbUvUdRQ9nrSabiKFxGDSF7O40T9Z
K4c7dhmyO+GScms3iWewpitY0IHVpce7pDRPYTkZc4qNdAWB7IxoeHV/FdABsW+kyUewRI9bnNPf
JFhJKc8KlNejk2fNmH31rrv2sLIBBJhq+u4ddB/8C5nf9jg9elkrlBx2tOyuDW4mVWfQe1lkFni6
Xyco5sAxi40uKnJDSCA7KXHd3ZFBZXqjV0hQs7r1cZ8bSXZsAXWZmJSB7O8hmKOIDCnNsWheJ5mM
JIPf+zvqyy8ldd12EZJ1igKmnqEZKKPcxNY8MxjbMEPZwvHmZWDfSQId4KYEXpugBLydg00Unx5k
t9WzhKZk5R7hZcdT8JQa51KIAV/N69LTYCaIOF8kgdesuIcynhTufgjJAsTau0D8Rn6yGjsLBfnm
viTqWzlbdSYzVBP4xgPNGB0mnX2+d4zMxOGeJMi+v/CDJPy8b9jvcXNa/1KbKyyOaqkZUV0WgBz3
rCo75Da2mTOH4XMabQoAagSiK2Z/OpL3gtA1BmmU5bnd2GZ13hFUmqTW8Upy9cqdrO67WxoZhSFS
vD/r4juU8BpMBdH2/rOT5gT0q2/DPOE+DRAbRvse5SMQF3MGE64SIJCYDZjfzCjNXZzhtYKIAeQQ
AsBhxGzaj3OlpTLHnrQ6kbSl+5wUjIkixw0U8//hcXfWZYpTmGMy7nAMdPGLtrKw52VLQ4FzdILT
iHxs3Ke+3DzgeottI6So2TV3Fzj3uIV8LD/OQjDxUfH04VBvkLLfBbC7R7Rgvbd9bPUKUKOZ3zcC
YKAWN95rRj/RiBfXfyZNxibLnGQbHkPw68mZj9L5CkIpgeDayyWi+d7THvAc6m+JT9JCUk+raTHt
5zoIW4QyDgS3SAFTZAbZWTC76NwdryZ8ffOw0MeMOWneXWBg1OsS7mSv+lSiTiYjOAPyFJa+iCJm
TwNdo28SapHUgDvDlZeqo4dsS6eGKk4FoD0T/k+Q3LkSqXgJhwQg9SYoY7ADgNOXdkUIA4WNVect
F23v2xWVhniXSFeDsmVZJb7zmXInN48jh9aERJGhMCHspkrwO5m/YeAk0mSCyLo7zGqZN2jdk/yn
/o9T7wt/ox4cThrvZSKPd8k9gvtmKYpoFjpKIdGnDQPnRbbxO0Hl4+aGBgTa1L/q/NXKG60nGgXH
Q2FKa3OZDnTLqT4CoipIYEH2K0WK63Zf22gysxr4JtOurGEoPTv/p6R0MacM0beH8EvyQ7FrHrhO
vgu1DXmb092Qot7efEKlQiIPArDXCEdFXSXMC96ibT2MEFK/QsHb7WJOuAU/3fzVigw/iKCR8Luy
6lhSDZOv9lqGr7re2HJZd03npge9wGU6rGq2tWnuLVCWbD6g4bVhJtjJtfnyNodCswOdpAM3U+U4
VPF618ASmm3m7wLgFMY29bawlXtpIx4+b5FNIUPaD96c+movfXFYPgLNif775l+2c2SQplta4P91
+WbzLQ/xSgfSxLRE+oEel3HZkP+9DhoWBw5osmpLk4VQI8YFH49xRqBKgyFWbsA9+uX6p8CWS7oQ
ZDDXjLn0XsuUrsck1hHhmLqctEb/I2s+CJ7KmE3ekuaztt2MfUMcDhfVSKzCW79lbAZSC+/TYZ6p
PeRIQO2/1lVzNfm9rtmqiRloYb3EHDMUbcg7owx+yRFvBn0RD40TKFhAY4tvNhQABQ2JmcAnr9L/
/69K9vvbn000KlNLqa48WTI9ZZ50Q3v2JsjW3LyCBzJoak13hL+GmuJ0jlXNoZJv/Ir2KiY4Z91i
4tSdZnWsTcJA+x6olNWkRIallPh9ap9FlpygOTl7msjkmdtNto2tCLrae5SmcIslucj/WiMkBZHn
s62EeFyduviQYnYhyO8jtiZQpneBGnRVRclYUP1S69DxTHvDsNlMKyY773FTFgOMjlQbB+SPQ1DD
a7/OiH91toMY60nN0RV64KKKxLtko/lSs+tSUytrw80HiO5jWhrLJ8GH3H4PuefjX+5OCkGMZv9H
ficYpA5DhOjldwyTXymteItDHMthzZDw29quvRL4rfC8Zhs38OK5vmIrGkZbd1SfnmfKWESb66u0
iKyBIksh7+BI7pr8BVsR20SM/TlCvBqIBcdMyYHfCn+nkXf4qdrrS+nR23SspPwdiPAfm4lx2xxq
Dyy0Aw4dJT8iEKDW7uSTjdOTarkVJxpni1sgzP5AO6HG+2Urcs/4VnWRVfNhfctc3KiMldUyGRQC
wGlw7MgBIibcvW2yAmWcTzI//O1+Wi9uoLfLrGapEbhc21GO8D8zPVYfPGjsE4YJzLT96V4bvFbQ
nBXxbaS4ha4KvHgnNEiMJ8EcjlhkmjeRT3p5oilba9zz4HQ7MhZhgeJR1oNuJ/pKCILhsJI5JyL8
UGGNhsNEpKAsKp4uAXMcbaUKfqwp3eTu9OLqNR4dAvCrWvc1xS31zTnAv+PoJEX7d1/ZGIgNmfIG
QoxTV+68Z3mmtx4Nsm+HqCyeFCcumy0RmpptFsfnfiG04b0WwII9PNtJNPUA+N5BVC+s2sh9JGsz
DxDOsYFPzjtmDgcpXWa+ctWSdhRABoN9oBZmNevLHgf4RYAAE44F0YaHyFrNfCpxlgMjBLOOxrNP
to6CBOUT9hrp8U9/MiG4aByxo3lhlG1Ss/zPFLsbIcH2MuNnBHKwLw13QH37b/YQ8vTeqBcGNXtj
8igRXy535b7KwuLzik8dG0rsj2ATEp1y+f3Y58IcnhJgNd1/BSQ99ISDlRnwDJVw6XCbeB1Exkxh
5kKwgNnbsQ5n7OzZB3wFlfh7If7njdxyvrFDQ9FnRqnS7MLMJ5ApElJmGerxgstZjIaSDQ2fE2Uh
keFDfIQGL7/K/VD89oz4qwryswl8lz2aCLOQpR6pFdesRQohLlJZo7vv/Y7eyXmDzh5zhVEXVM/+
p3hK1sATx2IdCYtWQCn6aIeVH51a226mG3M7BiZt7sEyLXn0sHMeAwvhJXfq1Yr4LAts9HgtbOmy
GW+V8wEcJzH9yqJyA6gsFaCd+SwtnwPRL9vB+Hccgt/R41NRj3YkmCHzhpwzRNQLAHrA+PCwnujf
GGw9GQPbDQjZMq3je6OVAj39tEOXuqtV/YEVEPCdVJ9QQCt9c3KxmHzEPnXSNL9rRgvlHt5YA0KZ
xdWAPuBXRCMAAdNrTm/TVj0O1rWW1T1V4/m9p0ysMEOkVJkd8V6XjBaCGcyCJ3jW7txwUuTXQR4G
DCuZ8oim0pDv3umjX030rg+pCbcYVaj4IUo/nAFomv65+ff6VDpkoHuDDzJTscpHUrzxa1gXMXUY
LqMoDR3G0WOhg/586rpRMGZenF+C1+RQYFkcDxX2L6qlMLhu3mpMdP3irAawhctFd+9jk4YileX9
PZM5THCZPRArd8AUU/baGsBTQsQugolGRpeAaFVstNGLGIK7AeoX/PPbqhkoWIQJobgcVR2fVsMr
iKBCEaWBgnKmWViea9XSLA1iRw4qWSqpKknx4JB+7Ogfnog/wtL7JqMQfWpW0uYM6ben2XTbFj6T
fgjGA2mHUjpRcZjOasC7QKtdFDSJROB29vVeFP6rYCfCQ9SWbygqfSHm2reGfL/Cqn7LLiGOaw9X
WPwGhr797LHef0YuWDgR8uuaXRBsZmnwkkqDoVzsvbyDrcxNVTZRa1BBxfLldrhP2kYESoCl1WYj
wfdDayyERbFuXYZjk1ZqYqU+kqsUFmL3uiekp7/gm19iirO8GiRVsc/CijOkvvzzOKEeUrKkTcMh
VzDDYQo7D7O2EKdoDFq7SspVzgQlTYe1HTvOjERCRQcb2BdwFM90CMkUc2s1oF46ETMuEB7Ghoyv
LkIXK9/EDNR37PRLfjpu8QAD2WZVTtUILlJEKLwiDm6VrMW04hLxJJ1Q2y3se53FYliQorIvgpJ6
qlnJWJE9pYgpXLGba8TC7Qvzc//2UlnYsklJB2nw9d1P5HzWUsSihtqJ0bK0G+HGvypSbIbqYcqy
SmCJWW6sFlnxV/X1E1Wq7HAu9Ue+Kvx3i4hA/X0LwOVBp7JeYN5mqUa41qCwwcIOFdARO+2l19D0
dw+vo0/nUvqmm5SDWEizj2316hsb3Kgp0C4PHfQ6WYO1n2quUuEunV8pEGBnSmjxdMRHz2lKgFI4
YeFX9PjJxfX08jQmxcV1ipEB12MZHZ21h2qUv8icU1/Hm16A2rjxC5g53liq4opbEooF9d/8keYW
sbWPzTyYCmDTW4Fh8odLCK7WgOigu9om2gB/kd9/OmZQevJ9YHSNR9I/ejwuukdUnOWK5DwejIXE
LfmM/vyQLnEW575SJMXMfXUHU06g1ZMRnjYuh7JdGjIlNrGLkxz5aEIhK0+iXvJ28tiRxH5GYg9b
uZvx8Vb846jgwva1At/XbrRY5S73tljIZTFOEip0NkW/3EMscFWR1yYpC3yYOMOh7l1dJe5iuzb9
UIGhBbaez29B/a/r1hh5Hz2Muv2ja3GMD2XH0Fy9jfkzMsB+CSmvYBC9LAzR/QtFGaX/mFUI0yB/
XBtZoS4csZ187xg2S/SFexcEuxU6DZ76fcRLdVfU7/Y1vMxKI1grw81TMlwDqxs/YcdbDgeJHuBx
0OOlTR6ZHHfRCMAbA3vsQBstZrRZBlLt6f17lHIHcsfT6wMdUicwOxlfguUV1duxHZbc8oewY7+M
2/JAb4vOn6cLyVqx4F4T4UmbjfzNY8yXQqYkEyzb7fS8EoJFMI+H9ffWkwIUPXNyx6VDEcGFVEwf
msmwbZ9Pl6hVBHQTCBbwfExBM0SKQM4EBTyAJBP8pa33siJbk7PGWYWo+F8NIhdf7KPcCg6fMQ3l
uP650XeNy3oUQ+J6s7IFjVjEEighOl5MGMmRuJ/CVNfNoT50e96TmwMriCXwr6ZVUuDHiiz4abto
CdbrZq4JBqUSunhNmXdxUMnzKesHuGVD4fHV+2cYa8y7Ja4kRZRiP4pbI2waDe9ywHFnMtXn0Crs
vETWs2+wpnWGfzRlkha7JK9cJYvAjbIf2e1Eo1DFBsSr8o0A0nFx+KSdDXWyMhxIzJlokwUw+4KU
/hta25xY1TQ1KLQiM+cINFzo3iw5o5YqDSVeMAktiHoLJhb+cJ6QIXrPCW259r9XCPw2yQEVCRT6
PC22SfVFeDLYArOSVJdttfzfFLx7riyFjSv1dAd4IGxUvfgv50734A5Tl04SGor9v/r8a4eTNphz
oIaVXZPrRr1BuYfiNfOWPOTVYOlyrIr623PviBddY/q9rCyl5q5KQo40rdxKOFZUSRdA+LfT+CFH
1VjbPSSIfy1dnQSUaaD4BYFQnu7SrOLyyAhhz4t3jOjpBd1vmsbwGwXG65zTk7ITR5ZD3cNOhKQR
BCeBbdxFYlF2i2knM3ZQFnlNv8F+I95EU1xL6Ys718rhU+ifRszdJselxa8XKsX93VSm3T9yqa3+
CzOYCaWxCA68DL2tK/2V1vbhULoem+Xw/o179D7kmcviMr8D82T1mdLMTo4Mm69muOyfBxYZ5FPu
lX366E/ZL3+1v2E5rQbpOqntjb7CN2TeSo0Uq/Z8nBjUsikt/Wh17a3OzMWLykvWWcpeZ3pR7C9U
LGhnTCBFlrmUIr0iXiS6VdCQGUnTZL/To4X0Pl5TJAyoQmaL/Rw2oBhVjtxqWY+UKt7xBTsIi6kJ
QfkwFvlHu4yes2uyxJzy2CO+D1zswofZmRNE45ZMXZL5gMK2MHz40RRWeSuw54/LHJIMr5qRrgMD
EeMBod87ObVcTn+1UcCKtSEz7nLYlMFv5cNJCE2z+jsg43XETjHb6xazeW8O1ufyIG3m6kjEmA4u
UCJU7S4/7PKsTfXTOYm+lhDOfKM41U1IxFJmf5iQHYQniXoWGxzjvwPtwq7ieSErLxasC55yE8Mn
vV6WxSHvfgjWVJaZPUYYkqeAAJ+geF6UyhBFDZJRBPMZV++Dlq1A4SIRX6b9uoxJ6MKGtsaN1AS/
4FK9ld5mGSHFngUdPmoqvOrNeBbI2BF1hUsNyKtlQj3LEHoptFktwR0iZnRCdcVLiyj3qoc1zR7J
D9W8TCm3+rKA5/VkcgYE705a6DfE9CouZQv4andX4rydpmon8UFm+Trn4fYxcFpf8sDsJIbVkiSL
CGbU5Rw5MdNgTomLcCc8cE8xoMdtF1WPWCejC61+HoJja3KLg/SbsbIekkydOQcg7Si2vqizOCof
KUjQhJaUmFUJdYAvwG/MvS8jui0ionPRZUpsltpsuZcBQ9/9MyD5XCJWqlhnse7WxIP18Vo91Uyx
myD+cFCudfC62ts5ogd29vjD5Vq+TnK0cE2wrNsNm+w+jjE+MVlxYJhz9PmsI0PmIuEuTmaLqTzo
TU9dfPfjUkn/oNm74g99NRDSvyofojO8hRXP717mDL+5SY38b4ZdZJ1dUt1/SXrmdb4odrNonXYd
keoiU89HobHowhnd+akqlkpPxodYmzFEF8ekavgf72UUpAtLMIiCY1jsgtu1oFE4v6jllRGR7X/K
Atl8qNAzPsQ8IuCbMxjRnjomts8npB52aKjnflG3UiYkuHxdA6T7YXoN6V1r4p85V1/RLACPGVA5
mkzlNonBpsbjWJzy7vEo6SHKg1PN9snfPm8peMGJCihZnLS+cSs6V6ACbeY7GltCG9o043jWaoNS
STJ/8WKAKvONqCmqyUuMT7qM00mYRHaUBzdEu7heb8EPH5wThSGWr+en8b6T0LFbBzhVXNYD6tLW
FPN9lXPI4juzZjt/vikURgO/YmaZNOiSAmuwnR897LssOHH5WJCHVyBW6XoJlJ2hGgcwrwf2Msiw
kL42yHC1pNYATG624JkfrWE2wiKZC6bErvfbTIL8eU43VDqy1ItY1w854KXkMSqP9aPK1KFtCmV/
gNXaB3wEZMF2EGMSaavWHhBbN8VIS9teTiIBUgGgfFg6OTUeHE4Xi9VVLOV4SSABDpMlT+aOYnz9
03xVOCOxKTNv2/zJ+gFDiQZxWSqyqzA7ZTE2iIunkVa3adeyZD47+KKKLE7mkcUX3qfNkVC6E2Ja
ngIAGR7Ie5AGlZ8W5DP5nU9a16LRlmpTmfW2XvimjmaBdPD88D8Onv5c/HRU5/JthqEFIxzou2t0
gxbZhNqe9heKwN0fWZLawiI8xC//pImL6JlHVgOkp4tsOQT4dLFos38TGgMS144NfurFhWwwhcWG
Idk9KLXsuqfVxR0FxiOTZWQGxzqbWFl5t8OaQq6afUygJTDbT0wFt2IuA47TtRigepY2mOk2qurY
bxq5decfb6wOsXUGqnQ7WjFwIJ2TtmX+Vet3rD9vUjdjwlTvwWRzaIMAFVfUaT7oJpI+3l8r+IQB
iWF/ACtadvE7/c8uXiu6IxwMImdw1bSWhDojrB+E3rP6TAnJuE4zr5q6EnnMAImPTl0Y5ath+e0m
v4u9G3fTHWxjjgcSHn2im9TR/++MSSwKopyRfjvuSaoenE10DKh55U8KjhM/YouQOa6yz2WwGkNB
mX8g+l8odHF2NsOXbUspwp5Ad5aZzN4P48WKTxMf83baFKfBC1LsNjyNqfnnPLStNZS4Vib/M39Q
oL/cKRrGH9Fr7uGKdLzXO2WkQGffE+KNerOF2Xh3vjV0m86Ac5ZfMvfU5uKF1TMo4Ljnoh5sVbiW
cmi4AIn9VhnHoIB3od3yOhWWH6dZEd8qbpaD351WJdch4swZ26p3H0k8HG43OPclSpY/G3wnuTkW
cUKOjxUHCQ15yf3NR0MQiGF61hi4tQxk06NU+f3jvzdmNqa2CfiuxU2OQBDIHiGB4ntsfnXyM4HY
kaEbNy9IRR0oejeQxIp95jCzM/tzNlJAqjtv6LSR0ml168NKVjPj/6J3trIGNzl78PdoaqjA+HlE
8lf4KH6Yw3G0PC2hvaGqfRV/BCYkxAkpS49vKym9yVXPikLJA1PvBh9ToR5HLErxUIBz3UVzbGTg
78VOJAoSZajKDOBVMoz8FeOXI2XmKhfspqTKVWg2Z5RH9jF2jW+6ziksg7exwzxEyOST2qWfjogp
0orWRuKj5c9akzxAjyUzsLmtVe9K+3vLgbbq4x5VQZnO/tQM9+aj72K2Sd8mCTr+eKTr/sztMRR5
ieuIdQUWsEgR9LDenPLGMqVz+EhXw6lW3TJjHzG7a9Mu8fAUtROuMlQXIQSt3fk7R8eFxCFycNZV
qkvgA93n9WTVG2Dcqp8xP1jbbd/Seninbz4dxqlz2xp7FhaEhZrTukuIhD6nQpRqH1pAOlWNZHLr
AifdH2RCe/YHrdr1elDpDumMh/bAv/K4fbE/sGoqzXVJgHWzeb5TjSJReLca7iFwfm9mgGaCtpJG
tI6qe//CKGnw+iCCNq7l4mnyJ++k15XutajsYK1p56JZNlS1HQ87qIT94GwoKvMOs/uTfOD7gKep
JGGVWV9deO1x7nXsjfrlabYj3z6gLy+TXT0p0bSuugu1JrJgJQ0EvQbA7MPZK91/4H6I/0QBlAQ2
lv4XW9QmHrKCbw4nNG0OJBLZGFvAqzFuYOwY69uo1lnF5gnCQVjns4Za5ns/JvvHWCyT2Kk3pz2W
GPSgyPkuQE5g5Lf58HLlU+UcP3dCR+pAhoB71v1J6aV/MF3v0emqd3Pn2sv30mjpZ24ItJRepZxM
dgLkjVfErCM3bE0188aAe+ZDNZGWfLXcCjCv+ewuBJi9yNOiMJI57IpUb2FIG5uvb4lAcgHXXdMn
sNUQHqmtOoNbj1HqUdKVO7MkMnEpMFrEUCJXjWnqpc9GSCTPojUORiQeWp1C77XwsLLhqd2rp0MK
vf/zD5pRRrD/IjdkGOJkAyjSsn4AK4dbxAnMVKkRy0Kcur4zZr3cn7jNvK4pneu9Xm8+k0DwjqpT
j6VbsDHJ5GE4csgclnhxHcX+fSKTAncsCHFkhZf4uq5Jkm1ggEBGC6DE2Bx6HLjsAyVSL2tvpb61
L4YLCC4mPYhvuzxu1tapLLQdLans4BSJT3PjllaeeTsCdX+llTHElqcosjsdOtcojjCvvHL0Rctc
aNJCVvSl7oQuhX4YN+Wqo0bNgLz89vZRW3PCDfHx+JvOTjFxN/ZPtN/PL1dU/PXFiHYw5lYUcOIA
CEhF0ihOdIdQ6GLdL+5wwCoQZ1WerQtKMWB6Y+3m1ZpaikX1417Z6SdkyCEbgUDJ+AbmcjJqz4Q7
S3iHGVqst6Pw5m0mvVFW6LGnaDQnRNHOHndqcktlr3d9y66LTQNtgLXa0XD+dBIEmmnz9AQFoYxE
ccE84SK8Fbfb1AGa1GsGTEjbCMhGjZHq6DXmJM7yeJSUeJT6TNcJsH70RW3admGNV+01AJY3lCn0
bF0s4mXPJyzjdA5Sn4u0ydvZh5MSy4P/oJ6oSlzZjw8hsUUPZpoXwH+xJ3bC/Vkm5japsL092So9
zdFhRW2675SgY9TTvQw/FcTcsRotdZmev2iaIrZRdmlzLF5VIPNiMnC1uHOwEUESY28F6rWeZvmw
Sm9Q/17WHMdjdUSyhRD+xKWmQHLSjoGYjmgqvP5bel+ipjdNbIiu87vMprYkZ8pE3G/s4mZieJP8
nuaq6QuQYLs2fSsp/LFKOykz3FmB8SZssK2r8J7Qo1W/XLvXiKvBjV117u94dVHFnckJFdKGk7yL
6Cmmek4PYoOEW86S8V+VV4CcU9/zfwKeg3TuffQ3GQCpHjWOmmccOfv7rGuhYK8qs7M444nzF/UW
Cmy27BZWUuFm2KBSxVVBDJ6JlUCYW4Sfjo7MsQD2sxHS+kgxnVatpxN3PN+mklz4uQRIoYwir1Kg
r41jLVpT7Inc7YM7+AfKF5Hs8WwY72UMnZdp921BTZ/0Ic+JPBUIW2B3/23owuIhSaGsOJDGtEVt
H6W/Kj0ywfrLkRqtrDQypWdE5TpYaVf+Yp5l6wuW1NTzy+w8IoDQwYud0uOphPtgz0HURWsN8i8H
Tuv07PCmkfYxqLUfsn3cxI6/d1dr87CQ3E2vS5Hc8vu59mFDy/YjAMoSVZ9plvZtddC0q0Pn6Ebl
tAX5TI8Wj2MldQlgzm/oQ99ceJO6+upam+sa6YLVPqpR6ve/h5N2YpU8zJsbCF0y0RiE1u783fZJ
wbLuaLnfWKpGlBwMKCQBRg9PVK5OvvZYL5alw/quJYWqHABOzs5BqDROCU1HLglvCi8ZzXjPQv/1
9XHFiywVJL/ab4S2ZegDZ+keyjA+eXk/hZOVRiXV0CjraTqVXYRzcRXCAtUJJkDkqVhAANkeuxje
+9pdnVCFQJZOrZyxNwv3Y0nnCxTirH5p4YmGtlWxpqdwd+3vL0ZD1+soucxS1dTmwJJXApeXw9XO
LJSfvy6Io4BLHVKHgKa/V4ZwZ47ig+Eukxg9nPUH3iMpuy6xlQ4M/5l7p46D3TgDP3DLVUW5Pnfu
7UfbjS9GOSYjhoXJfw0aDLlDATEE6wjaVB7+xewCZGD9t4ly4f/wK5wg8tA/cF5CZxqZYwED6UEx
1yMiQW//SMzi3byxPBUhLWjOF3ZXbN7KO4dLYymbgjFR4+TkTyPPqdzVKfgJIFrq2H7xxLV6cerO
Zizcx9oZooU/mQC4FXB+IItBCL40GAUNvpqP2QYDJAHJLMcvp1r179cpEtLXSn3qKgzfGW9EUXhL
6Q5d4s7YUI0unGlVCiYSPr0XOw13qo+PYmRDy941rV365vt1QtX2wP0urgbH3zDNvExNMVFcSAQd
uZHl849rpW1V+0UF3MiJRzqy+cG1N4Sce4pxiA9GSlkf/yL2ZhgONgFPVPKDhYqMl9Z/wVahPABv
P1RMTzsqyePclRHYZaab4opXkhTMkdKJBC7IVCYJ+/pH7PLL/54uxZObvvQVQCx3OgJpfFA0/DU5
ag5yW1gDflTh9ooMIvCt+Wa39r+JAS/k611jH8K/UXFCGqg9SuGAm0lAXFM6AAQ2dM/3y+52kuEE
wNwZtbaG3qlsthJLIt5pKa0ZobQWDFW2zgBbue7cjs71vAB8QBXkU50RDQ5V+26ApdOv9Lh1xGds
zces9KUp/mpuaWRdRN+7cBCNNR4YaDShX3QDwRZFybc066RadJMFwTGtWBA6grW4xNgJYQm1h5xF
Hsf4j2FWOZRYZ0ADItgV5y8o85SLu7z6v7KBYeEST/Hnf1ezGpYwFS5lN3ic9mjVpRCpnrC8h4SA
LsobXoimMrJr8L3NUqDoEAewBiLUfWtnm8KgmJonw+d1E2mRqfNuDAY0ElhYJ1m6YxDPHAu7xp94
mCR7xTg4dtK65AG9ENL+o3CP64br2351GqQgTFGFZNdDnP/VTkIPsHikrjK5s6/EyD82UtpKO5ZD
nRyZzZTZ6f4usGAWLcv3mNroD4HAsMdtsswNAskpZjKOeh+GrWQlIyVgne5hMcdbEEZfDUCGOQZY
75zO3Y8Ts+vCLBGi0bcks4iQiZ1gC/OnIyHaGkGiuHTp269gZ5Tw7ftT3OXS7//PPjdeH3ebKEOa
aH2dIonEkVwjA2raH45rNjb0fc1x7NStVIDD2C/0g5a44cXwWPKPZBUmOn0igPGccoY3nEgBzkJy
C1iOOdOyYNOvlYDFu/cgeI+yJqoUxCL8wHzJEAXscVkMNN0lbB9jgne/7KF0sy1RiHGrIFYhteVU
Y8h/bvEbPhWuMMqHcaMlkdtwLOTUjT+si43hVYCCnk1dWDTHCiBijcRQsKUrE+aWjDJA7XYiLZj3
LqSHR9wbaHFCeLEUUDpwIw1ain9OR5KKDSwYQoCzXbEywpoHmcvzuV1SeGkpyQUUAt8q5NAMQxjz
ucbl1l4vj1W4bPb0giFrYgThvLMSVXv79FE322j8kfMHEfZotwAehwjtgdjU+aPUdBZ28YgGrbWJ
RH0xB67GXsX5iTR1KUtAR8UziwpCTQt2Hwt28iESwLjYR18n2PiQWvvznt2QyLH3NgIfmmxYNVFD
gkwL7i1RX8rwoySFwb7/whmaoGzj7+2/uic84QH8Pj62zIQWNMv1nrFpJacaalQz5tGgU9ZxWIK8
TzlYUp1H8RYnKllZLPGoCx97p71lQ7khQAJZRisN9BulYPoNuOpgIVFpnJfeFfYGpTQp1839Vp4Y
I3wIiuKz8PyakQAurQru9q0LH8EJNJhL9pakzo5beZi0R9QoT2lq8yblyHmVGdFV7dpOOIcB+jb1
81Hjt70vWFWPM6ekXI+Snu8xegaUgGH+Xwz7zAhDsr0nPFS4EmtIve1k0Y/GZ++R1i+XRNnlY4Ad
i6DoZL5EgGu1ZZo3lb1d+26IrMcW+HXK1juGbwHmCcxjrAVJh3ITUJuHe4q4Gpn5OYZ2J6DZkG4v
LFwkAyI0sKNkJUAGwr83gGwdGvrO4ieRFDv44Fq6uuVZDkZgFXFfJsRcbNr+UTnqDFNDH26adfJw
Jhu8oYSoE02MW6i6C7tvRZ73GZzo7E7/Sr+FQO23rVlTK3B7MS5BDPiVv9NTM0xTvHBHHOocdCXd
pxRnO3FtPbxTBBtCZAJ3Ho/32Mo+tvrDpGXI8QPp6jrSzpx4XtO20crXiPKEF/lO6F01BZaQCCIB
HS1D7L3NHfmLory7R5gBK+vl2IGbtkeabD5IBUZMp7Nad1o/gMNNLiXocDBx3y1OE3JJGOcS/fTT
izjmRgnKbOBe/0iu3fyvWqET/P6/7YXtVOs9JrxejP27NA/Db0hKJcNbCrU91XmIZgSPmwAhAGnS
3Wn8tu94zhUX5HgfKZL/T7jBkvNf0/t6nHytV+RTVoH4Nq9graeb5qKAFi50Kj/WCHbOeDYZucPq
Mm2xDedAVW7NN3+x5pFBco8kpsP+yY4gEV1axEz8818MVAMWH1G+kaMd/bdJn8YMzKu3A3eOvInY
Jqc/GWii7yxh7TMfY56SiVPrsoYbbGr3bcnyP8gLWpH2sDio8jk33G4NJumQ0B6Vu7HEBEtagPOV
DR/g4assl5gUiCp3RFSOtLD+Jm4gQLYMvcGGUAqCXY0jT2dnGxKVTyDFh6HAsi1KjCz3FMNdBY0Y
V541WklykkFurL62glu3qrWhEz4Oixc3DmQerLi35jHlORZXwGSQihsQRons+hwL/hQHqiHwiV3o
ia+aSn6VePZMPlML8g1T3ZvoecuIPJ/PULEGadDsyb1zffLb0kxO+90q2i0ZRmfBkGqovolnwWQE
j5LC4QIVTV4I+/Bb98yXucl60thdNiw1bBvPOGCopX7OztQNN03W0pNDHyR+s88Ju1YJyxvtRkgo
lvTFH7BcgFT8GkR8qvgala3d+Diu3TLbevOioTzUfDGVM2sCZRgbmiR8Whmdw7S1H6/9p9J/IizL
/VBljrdVdWi/hPLeE861akHTfZZkQhtGTYmRWwmaXw5KxzCs1AlL776C40ZqMpgdY5AyOnvsyv8g
bYGEV98AVhi4+9A+sUvgexpSduLIvPMEcWrrRKgA2YkG2sEYV3ZyKZOW3MuP44p1L+4p5ZB25YuN
/M5dtFD1N31Xv+Henqa9fej2RhhVW1GWE3PDh7CUAkvFGqUZDWVKUVC7UiPa5QchibuJARUZ/q/q
2jz4Ov3lA72fRbzhJVsX0DxQvFtfwbPAJeuVyIMFoa8KMImnYRzYvljL2GKv6kpNECfP0BSpVMWS
UYUGzmzmSaEEW0d0pHr4MceRbVcF0MeaaWYiJSU5v9rH5uFlNzJXwmHzePQeCBguGKVq8roMwu1G
M2VQYl2PjJZSBrdsI1Vsbjni0jQBUahiTzyDJd0cPtXGPB7GVl1C6OidWbmXro0xRj3LjOfnpaTN
6fMLHA2WSmCFqHIY4Js8hTcYeXwReic5SZ0mvw+Dl5koqFzvxF/xS+xWlaor7ddIktRFVrH4PZh3
8x9CWKgloMEXv5MeHipubjNX5rDtnYqpjcp9GEwe1cI6pqBBQFi518htt6XjCgLRCQyvw5w23Rx2
xV5R1v/d9Bgg7JUV4GLasY+7m0x0SZdQoX7LSCzXmnBYnaVxXcgSAVIjXJgiKpYnkwcuSSSDYWhI
b3AwaSPS8E2VE+l1zzhaETFXXMS2kCnHxnffduRD2OaWwOy6mgFFhDMLrGr0N1Ijjgpczxega/z6
B8ih8EEU+V1SRfmmXzVgbfw2PuC+VgwnVyAqUpUjm7WjU3mvgbTw7qTmbVdMbDTONQs8YHzPrUzf
ryQ8gvoPa5xQOqMUxBvpR4UStRMgeGeX0Ep/71WOBJ2saC/1hZaAgyQ4tnxXGgXT1YSDerhH3htu
FTtaDh9AoN8QM9wJl6yj4JElpP5H1rNuTdLfYvPXvuGRbWsJ0ofDIYMwGwp1NngR0oDhohARnPtO
uMX59O7SXoWDyR0kJI1UmvNfuktF/FUDMrvtWicnxGyvTTT4eMfHDqLPChUyFJDLgSjhRXQM3eQ4
DOrIjuilI22AeN1RfepOLKK+BKilMof4lBTVwWjqCvElNdhyMQBzWlMVBAYIr8X/1Eyh5gLkifbf
x0AaTzOB1m3fwKnZaA7Cf86izEDNK6vYcVrcQUsg+Pg/sqWQJ0TLPswkctCSWdbogQ1yMdG7xW7z
lapSVQpCdDW/etrv4cFsxPN/ebamR0Imz05eHU8K7JLPKxfDiUbjLPVg0+cV3aowTA4JoakVfNIr
nyypyPJ/mrkUh/5ICaypYY2sjnOqmFYYEcmAasLKAAkuGFPrCTA37wyE7pdMBUF0DxGb4uJKtSxI
KuL25sFCdI7tDkHgvrGGHcdDtw1dN2BZD96UgOhkbXWnmcR4z17tUGZWm52eMrJXQLgeNv8GQb+O
f+zroOjLW3dSClMLbW4HNwJGu+N0HUCNeTh5I61Klpoo46JQN5R/zGlEgsxMzh3aJ77F7CsKNzRZ
mJLOdHU7415cgsI52WAdeTBpWxnuozO6jLs5ffwgAsjP5f5IPFGTLeqQIMM/RDNxPWARrftBnFEG
02Zk8NhOTKLsmtLVUJPFsauoIomT7QnSGO+bjanW77U9z7iXkuTdhweYDXWCV3M8almzAG45DMQy
KaNOwDbE5NrBqYR7x4fjKHpgBgFlFgS1KlQMPKrrw7buD5NZCuS/X1DQujBm47RlM/4YYOu+eafV
sz2US9Ih5I53oSgqNS8GdIfzUkNTWnry1IZe7d0ESKrIQt3HpSQjLlBg4D3wdIOnWsa9fS81pBmE
RPoH+IllXG2ey7psTjwrHz9SzA46+gSu9WEz5QdIlDM9WQ1ysfWkEOGKKUHQhB7ZqkyN+nPX93VY
+rGCJiEB6eyrN7ORhvpRsB37wQnFfbGN9DReja3vTAwrzK/4Jjmc6nbFnAdT193Vxq202XZ/HB0L
i+LSYM+G8YXe3jVT1NOmzxytkc47u9nMObHSh/dugGPHt2G1ddD594Veoe6EKWWLCT0rzRdGfahk
tCQIWPeBEDw3wMdZGxqfZFx9qHREq6QtAxWRX8Xgt+c24JeYY8wrHAaF802FAeBb3Yayn5ZxQ++A
yXxVZ7bHrUMyJCOQWGXxaeLHITPMhYD+ropFIsjiDllFdMHt0fClwVhrEvlm5b7JJkgjjNE5W3ad
AnMZT4jIOUI1mKmw+RJLbfb7m7jeXEMJYwMZmUj2nFUHsx031x4VViR1ssW8Om+x4WIvWNqCmGuW
SMzR5YcEWUNarbZbn5Z9zeYkSVmP3nxY/J6m5Tgs8DPr28+2YDksc9OMnqH8/+YYBb6GIVkfRmAJ
lBJ0UFNOdKwbgfOtw0z2Wd5LdH6mQrRskFfdPehjUsK7USdP361ptk99i2dH05cDINHwFtXONg37
8u+8BwKIxEq9wzTV8J1Z2N+alrWDZC66R5TuDWqsmqTHpasg0HQ7aIEIbFYsCwesBkSQewDHbh4C
xrwt4N0oto4fKYxvoiLyUfqx22phCQUK0/w3unpcHjYX7mvNFBXE5zrF04o647dUJokHFasWO8cr
xKKDyqRdKv3MOsNF+f9m32LwTktgMC8/44kIG0QYo8PmdwnWXkSbxknpLvtA0NJvOIVE4Bs5bRPF
6Wsk9hW0KezpsoDuYsQa9HwYQLX3b6Y+nfQKzCqs/HHLQe9/H6WWlw/Z02PNBsldTYc6Zol3DrqT
Qwlgb53D093j2F/chJN980eZ4DGAUKYdIu+a1DOoSwYq7SCzcFnofS24wS1g0vGozbAk74esksjh
TaScP8F+0HthYeSQgTVLu2+W0woZvcaTXB7FdBp49wY1l1GVnceyP5EfwxSfwkZ/Cd/mmrZ5uaa0
IJHxdDJjCAD0Iil3W+PaTa6ucWD3lUUjsTCAeuDpwX7RIPfHWFkqi8cgW0PRV6iuu+tm8Iz1rch2
ec9Lrx6SVTcO1lzIrbag37SYsbOCNiLapkn0n/GMuKSGrEmf9f3MC4p3EfbvUwCW8FQ2KR9Ig0FF
ktkG8TakR1tnpznYoBDKjBh0waCLxi1V7QVc9qTlEq3JkjWFD5Wioylejbw2wvMPR+2AWf52ZrbW
Lo9YqhXJ/YcfqZhMFwa6yEf3Y3i9tyikdw3KrMUyNP5vlxGtsBpC1dlvSS+whw7el8h2kNHg8zf7
gGs7x5MxT1+qVVjjcbM9FtgIP7aUAQPWQPkaKUPk7kDY6Xu5M6i6SBis8rNviDVvwLfsmwDum3yv
+mpNCkn0hERbXv6oJmRbJ/mtfxchSmoFjO3RM/LVA4uVqd0p6haD0ZQGc8kNUtUL3IPrmoY64h1E
XxYMTz8gQQuOYRj6qQOVUMZVIkcHmxashDZFfTdndXVRupqJ3E+0rEVcY6E4LjS98D0Ie5uG2ELb
iPrQr2y9s2LU2/HAnwExI0wxWXl0+OKVIwQMyJ3MUtBzawsjyMwY9YLhdpMzyUgX1RSqk5f9t28C
pYjxXXWPOChOnge7nGE9V5fobyOS91/O6xgcNXhDwTyohQ8XJJBBcaX+WVObRfAzUTqzCA/JR0nm
KZfghyQuQFiNgkGKE3f5DO/NammYWMyt8wf1Jyvy38JES+We7HlHSoWQqyA0Fsrqsj1AB3NTM61R
0Eb5UvnU3AQiGqhnsIwknhJ1RpX3Xdnik3b+nj1vYV76TJaFJGNor0Q7LOTAa82+4zyI6QHe9gZI
iaO/ho8+/LwUeKc2vGZZTjtdi/T8h18p8XqSJvWA6I2UKfgTTKk3WKYKZuLs2D4Xv4a5KNiod2Vr
90wr1j05NzGZJlxoIampSzsKVdpbB+b1LzvW4BJTCqH8cmFYTphjqN7bj9poEaBL2Dup52G8R/iR
mgBNNeIN8QI8zzHcXjxGKpSIXrTZycetCD4cVhTVxdc2zl8RhtYuozagTaE9BHhO8oQFJamdWIK5
7oUIqTFrom+r0u3KrWlxjEVEM1rYkUgWdD66aD6O5rBzdYk0RISjGz+T51o1klxO1tUnonttVPtb
JqyzW2gj/dwwv0cLgsFkwmIqZ9FuS1EVSKxqXxzOLPM+eXzWcJ6AAYXROC2ka3ZAtKa8waKTb258
ulHmRSx/4dA/OF6rNRk56aiRPMk1rAsPTDKWx1lJItnwi6IB/MvJGSh4B6pO9pfjUjYE467PGHmj
tzWqPlRNYFHP1meOTOLEvfXmMbKoUaYLbiaaY0wnjZVcKUEm7OElgCzCInYutJO8yvvEnSs92U6r
nrQfE7gRnXepL93HwiHvkn5ZTP/zVV/+IbOUJEtQsItDO5kfsP6yokdL5BCCSp5ADaGb0sIsgZa3
NSLlAF6SuOCl9MbqPvLrbDrWQ8ggMlqHTDxSFloiaVgfKwG8+t5QW8KK80all1jnmLF6SWmQg6QF
BxgvWDhcTlmkbbU/8tJyf/5wk2rQrZB7hP531xFsv7huVWeY/1eRHIISN0mprIYjZZFtXCOv0HuH
LZ2ikE7OD6brmnnNml/rLlDqV1POuVCk9osZxsvycGSF8hBMFRrd3QCrPa5lamE1CjKe4YQ88FhU
G/FoTNEp6pqO+THWBhfvqZrTnefFN/vBgRi+4AQbNR6CA2QBNkobnMlWvuE9LX+lsKoO7fzlRFIN
aVa60JWPyeM9qy4t6pNpMOavnPS3YqOlWEL8SlopDtHIVqo6157Z2C/jR9mEZQt29mS2g+DEXy9v
iV+zNXchjrGePvm1rcoK9n0K3L46VppV17cgwFlK+C1d0yLlPANI3sDV3Y2fEjHU8hb9BoOaefkG
arJlMZNUk5uBJqB2qHzDmEPfpmz1uOUWRyXf5l+azHlNH4HI1GRWEzEXtPLIfNeG0/Gvb6LjHKpY
oGmY3B4tUEGlwP8rMvZeA5AFXVQ4aQ5iQkxURMb44yFTyuxK+JTQ3qWcm8Y2TxWdtpZlCWX+/Gcl
1/cFujgNQY7TwXgtjrLzHg6XMh6bVDh9cQy9BCy6JueA39pzM1qKO/ZZXVeqoeg1W2h49cxV6L9D
djtX1JD6F6WQKMOj3hi+fzbHhARxXUwirKFQP8u6w7SfXbhXgKJhgJv/CYuzKKgry28xJ4qzq3Py
FlEQUt0D9zdcUfc5GHxVjoRHjM+E6YCLq8K2+ATccWkKNL447Lo+ttF9gnCVZoGmmYWOgQgKGP1V
jfmUYzHlyo+xLKj9o2TVQrrpmx7VJKJR0td8UWx3gBl9Z20StmBL75FM9i2cCCUfRocgrxSPpGCf
UM9u3Fwhf0nT/i5lo1g/KuNsQLY/cSKAHTV2tGYIuKeKw5PVoEJyAyzx5MtAd03WoLMR5800rvrE
rX7dO8gnjNwGKoj4YVlq0LzyNWCdYxnc9OmRmwi+XvM2XSefPJrJlNrdNBmuZ8YbVpd2n3tP8kmz
mAOwYKs97cRjBfo6RRhIyEJ8kUU2gkINWZccXWUyreJ70hcWSmR+mUcCbv2PqtfmGmEG11txv33u
tvHmZOSj4VCN6ymugvdZXBprZtexCE0rGNDaWl54p0p6+cxpHTzMJTsWJwDY3vptJtQTnr34IlRz
9gNYyipvDg8EXq78DyAl6nCdTyMmAx9T6qHiwCXv0xUn8UmcNO6P6CvRlWGhMpXJd5ql5IZ0HH0E
0tYqJtRsQYmy0X3pYW86rsRZrxID+q8dcli0h8oRaEs458WqOngYWHSBrcEdC1hCzROMW3tdIjIa
xg7jPErho2T3FnmtBINwipTNWZxdO/ItJqj8SdMGHU61y6qbi+UY7/vvnuhQLBAVD54ZmGVO97bH
u+tY07dIDCvR2aEfsCsqHUQt9oVGWUGZxknhYdufwHGt3p7ODsHIxodONX38/RdKc0PcpI/Yntal
QMumzMpTozdi/4JaGcjUemCIihCf65GCpFoGztHAtcizRUi1HCk1/xwzJ2skIpR/3Kh3UAIWQ9Ms
IkqyLdvcoRPc78oCOYodXQrSCq8sE8tJ+CuvSLuDLqhVcLF+F2NrMlsiKHVJrgKkZyd4V55FSDBg
T71f2VLnj+Olh0IX9oEUPU5LQ3rXyPD7KMyvdDpMXNLnwEvgfN3fotOyckX5Vw6UE3IZ7wWfUtZN
xLJQcnCj4dDyLVd0vsEmFJGQzKLz28AGJNCAq30M8yJdesO3G0/7WHSfgPframCwWEMVT+RFFj7D
Ze7ZtTqb+WIlFsUkly+p69M5YfjZIdy57Wn4jZIK+N9h3Kp9WduXZDIvL712ofPsQ8T4F0xTuHAx
q5qx4jv1YkidUmkPUNqlxDMS82RP8KEvPSy5ZSbIbJOYSNqaJ5sObOLhf3DmoiFKg254HLrS4CGa
D6m06MKbtEoC/zo0SZyjMEu0t7k2Mm1kcmXyfyrZ42luXm15z0lT7HgXmT1D11LfU0DGLuZ4wFVA
pLEJwrlznx0ujo7u12BK0sZ6NtjZTPAkpKgWjEjh7EsTL4eEs4ESOJIeAkEd/+2iDux4iXAt0hia
Wywml2ZDI55raoKiqb8iXZdkqg374XItNv4GGt69FtGmcaKQutvNa3pO8f0r9wrwmck4a6nFs3Ft
GDjYwjg71vdtt35DNPFx62EF9iL/W5uT26BFNX+l2IpIDGG+hhTOx8VIFzl4K+bEVqvqJV0h126N
+r0bbIzAO5C22Ve0/ME08mauGYXZ/08tL0VUmbQlKKpcS8aG15tqTBSHSFcFUHiCFHqyJyQS3hZa
dKZaLXRQpQSmivydJ7DN6k2dmf99XFgmpfrVQs7CS+jrob+eME9bG223cTCv+bWjIv+Ol7jl5b4P
R2rXsd73+IMv4+DbSEYu269TGNFC1tIL1KSffK+OFlWBHugbHSvXveU9O2EYu4//jhP85JjOBwMS
K5Gip9meHzX0Z3vfQ4I07lKWQn3yfaxphUeURYSFIPwg0ovN17OL5F6vY0iBoJE0YlRwRhyVwG+N
z5QdZvaOo4AUVJlpi9XbxaHAgPsMRREzo8mE9xm79NFeAzqERLpdi2P21vqeTly2UNJlXg1q91O7
x16H29szMCRvN8ATnhy+0srV5XDo1bN/rMxZTfQ+fLJn+4EErIEpmsK5gC9YYRCN2gmkpcVzHFI/
jOxYjNsW+U2hdUbjg2w8H2Dlh4TnJYhxbiDjmKWllcH1eQ8ODI73VW6o0O/M/41qGs/2axFaOgGq
KQw6VR1vEEQaYIjx1JpsbIc8boOqaqq5fxM+S/xAxpJKq2JZ19xKAiR/rNK2N1z8rleGeplvnjrJ
tLnxWsVsCuqE9prQ0xO5uT+4ZcfbvE+d9AM6TMNx/yogQgWiD+KppctEkr5xWoX8c+FqFxwu8s2r
CHKR9pzUFpDrDnlDycyHHw73TmgL/XVT56jUaMNJYmne+aXb6875zXnhiTmamrALK1RuaBy5phGt
S7Z0frsZaeSbLu/0O2kWMP7ASSbBvYZZnTxGA8lttqxRqP14yV+Gj2HGuFQyhH8erNCyWjxQ7TaF
yGbH5iI+zwYScYJUjpnyXgrt1dW10s2vX49M3Y0Lnd+k0/NG+8KtRfbGGqpjfvztG/og0rUY3iCm
NRXfuyhJqzLxANs2Nku6ZA5fr9NQhqIAivCPzWDVk7zBG7C6Ti2frJv86DQNVwfg/vS7xEDx/KdD
aipciZS6+/cOwlCxfbgMoLFlenAV2k/uogb9JB+f75k7UBreY/p9xz8awmO/jfHkek5S8dpd24K/
sxOqMHTpP91JnECD7p3Ct4wwUDdcBuRxHjaD4sl4kOxJu5Hh/4Y3g/vU8961u//pI1WWBr9KQz0E
wgHIUXDoCqIQXqcKttLbeQkOkMHY+pULlSXpTojsOXt+epw5QxNVV+Oab38mRDkvWyZMLSOuCDbK
SMxTYWQ86SWk1PhEjvMSuuryIFwaY2PgOP5EhfyKpK821PMt0iWA1v0HZVAWsF5RlNwj7I8KdCap
EglPoA3LwddgFSZkU9+SFIxX11y4wUXLk1uOlu9UEjndKuKY8aZzdQU5LQn4jMIiD4nkgh53MgpS
Jhxvu3UMqfPB6VgtaYlFP2+wz0de710CnVIOpUbinaaoihsr+Vm/Py8M9oyaqEu6N1m2aDIRZtBS
1q0Z9ALSZ3YpQURHT7rqIBmwRnm3Ec68WyaNu1fvjn3qCNFnG4uSjzqwQ7M9WfE5r2rf2e2F3twz
SbDFPUBaF4b2Pt7eCk9YPKOd8cESSxGren0Ri7KW5vwTc6rNaidyGe6NQbHSFyz/zSLodw5JK3r0
kkFXwghnJFkcvvkIEoe5eTBL8rSC+Dz481j4Hqc9uIr3+U8VQ2Ck8p5fHiLP91B0Ah6ZZx/EZXjC
Qwe3sITM/GQ+H+sRrdSZUKPUVVJgcCLzECbjBL3/7C/R5WadMI3B1cdD3NQGjsPG9hLRL2ewpbEJ
lyXuTEWptHGZLIbI9Gj0VRE9VjcbExZz3pVyQ7aSIh4dfbsW7L7CSH3zBe+FUC45eHw8p2jHPBPc
HCzg8NpmSZICfO1TYxp4OGcsAu5D5hol1QMFEYbIWKkEjnxCm7Xo/gidOLafiS2JWMV97ikZoROC
hHFbw5W3S+clb+FP2hd+jaMY0to0owYrt0vuokXxgfKPM4n5tA+00FQra3YYNoNAettbPiLt2vME
YyoWueAlP6dd4JB2OgabapMh18euv95muLRX1PRJfHKPs4WHQ2zXQJtsj3ens1SqOgD516zh2/w9
W+nqC+I6Mwa8nb20PpWLawqyH50LQNDhlk0da0bd0v8U+utbbUlRTzKvAlBAXas/H5OffQMTgjUn
mj+CWMhsacBiPebi7IzRAT2r5QCIeAlqhq+xleHTPSJubEX4K5+pD4egHKcaIte/F1FKppiFVkKD
I1cq2rFCsjrc/csFng4MyAAYDrVUgV2aKbrESYovV3BLA8QWP6PeGLTWrMkny7B/cfaNk1y1LkKg
o+sFSLB79eYpjfo+2oAACFafvlQ2vfL9Uratd2z9pJPBYWeW08A2d58o6SoVh62WCY9tstFeW9o9
ftwTywJvXIhyBQ+FrLsnkeKA2y6NnpF9zLxMlxrf8EQ4DfzrZflsh7po61SPqovbb2P1+Y326QXR
EX/xKa+qL5wgMxxSDNtW+WimD1XsDPxd9FbCD72Snv41GfRHnVbH9WaVvBFp/82K3LQ9Va+J0GKY
gWm9kvH3CdYPj6eYpECdPilClQWk/VsgTpv56glTiMQQJA92gaYZfQiA94XG32KbQIaKcYvUuXTk
p5I/Zdd8Nt8iFvfqw6Wo4ADjZvJKx7eDIN3g16bb4DzoVueUEatAyDKluMmzch0gWWFooYo56En5
WbC8WhMRcr6n2PjoThIMf7z+dasPA3O5N3SHY/+/1OM20SRtONndg9Dtd8rCB4wtPP0NBifGmLOU
erRPllILsoeCJPoKv7ELW7UP+oYjpWX6En7GKmLasu2Dy3xQ+WR2E25U7NpSnKkficqYoj1R5EAI
3OQI/DMialICO8ZsAZodogm/rsnHouQ/olUg3LnvqLxT1UVDIiZxtS7koTCV2+E/J8uyqV8FLvnP
BbsTO146wBxIsuS3jBQXxN6WT2PHgGTIGV04SrsJPJ4tL6tpyzAFpEm0mmMAACxhsomTplRTl0FQ
5ViFHN3NK1imfoTFnVEix5OkRF6FIbOSsUOFEPhrQGBbrqx4whNRHcjLmFBDB5apCBHImu6vBmAg
86JZxR5MOWac5bGGbTx2hBu1m3kP/P9CtbvD7Pz53aPKnthIGmPr+zDtW/FmhJT8yEDBX15y08LD
Ij65NwWM7VgQrFgyYnyBi7htdn3X6nzIwTotL+aZpNVl6+mFmNhcHPpsvDgWjG5ex6RtkZlUbVRB
FMzBMydDAi8kWMHvokew9uHz3sUN5UH5rBjZZubnu3apodLYo2Jc8x9SnCnusvnx6ox8/Nzo8YIZ
SCOwMHyY8ZxUOTT2YycnxqeE6dpCv6FR/rNWw0+RGXsp2n+ldtF70hUiK2aPfGxQ58SVhrrnhjCq
6rfd7oWC1ZOsa6oU2Kl3Hbz9K+IsXDIOviOTqlXqm6wIymiQI+ottE8zx7sTC/6SgXR2Dv9oUY78
MhhelF9W4wZut1ZQO3bUam9t+rOBCSIwTmwWIGfwyLXRahMvCehHTd6RksQWFCVGDnAi/Y65ozh9
I9PgRU80ZtigLbKp+2OpIhkGQLML1fOg1skPuYoCvrLs+dp2PgH8XSeVwaOb04IB5bveJZ4AnHYP
mT0D4jhjfaYrx/TfwjcgVUFyDhiO3CjzT/oQajtPpqlKaGFdnLz21ofQnwUVQNb19vDKHZTCeJ0x
0Q4OR0EZoFPkmZriwof5W7vKZs6DSs0VYgPxXFhzMtfPO0q7R1u/gJSmkhE1eZpLENmvCImYqL0f
0pUrpbiLeO1zkzPdQStChWxbPXzq8PEtDOXbY5KH+JpzHHPIe3jTyk0W+67dTRbi3NuLwAvvu5GR
6Sg3yPlED5X+5VVqfyJCdtQSQE/Dq5glFqvOd0THIAdWQsg5EQN/ap5c9u4aqSYs3pfskk6i1vsM
mTcl4o97sa5RC7Q4LEYVn5KwjD8Cmu9cEiq3R2h7gt6QphPc5u4U8kn2Hr8rCRaV7Jrfm9+f2+Vr
TiwKECRXZ/Zz8NTJfV4jwvaltsGo2YjCxgWQJIcNtDkn7k4aodP2H9un8XQbL9sPTIXYKKAmAfGf
zzUComQ35U0msnJhzZXgLwccLY3Mrg8hsfYA77jrkI2LknQD1LdruQ765EsYOtTN/btgXxn4r2hn
kLh5VPs7lm5uOREfcHLDBiZ3T2hbLqh99urF/74Ikrm6rGjN1Hg/gTF/lCD82mMTbWFhVfAZ49hW
sL1Egz23lzsfC0Bq5kRfa4vA0h6Tv7F0Qk8HRcO4Sb28sZ8OIh+tooTjKFfAmJI3Ar0xAa/NanAd
4YGGFYq1cTT1WVyuyx/cbkzxzVVj7589RVzPqjfvAXZ+US6fbGEUAeqZZFA3lf2kAyIAkvJskTjh
bNuxZC9amWsAigrmAJvarPc8Mi0UZp/t6CmS2+qPtBy95SE6nC2RsMNnRoZFlhtOz2Rn6T/e+QA9
jvBV4U8cuBz5OOq8tKExWlJTa1KhcOb9bhSvrB3s4Dmp/A4x4NgBuCBHdCn1ISdm4PBQZGH2lRI8
DSTsD46ipZ3MZBjxKWn1fpFEykvCsSVn6k4/yU33SWRVt+eo4GpZYbqTfchaO7Wva6f+2uU1N1kq
MhCXuwTOa6tiYhdtTlnwfGjVzw8U+wvFU7bXfXuiwE9XQti8rOItyWEA2NHePQQnCTrnc18+NOhO
XWHhW9S56nMes3ZJj/uv3UH1VKJMa5ds8ZTunz8o48//K3DSq15fg9Hw5w7sut3LP17IgdBL+fed
p3BJQVsfR1YZRbSC6cyLd6k1GBVCmCSbMZa2EhCF2uhf+NVM+2uKnPJXK6AIujSF1E3MXcuiT0eF
QDwpV5uy6UOJ8Og4bDYtjUJ9JnpDbEAlo/kurzb++j5nr+xjpU68rF7orI8G9ypXKd1rUZLHToFt
LUv8L21YdXwbuHOV+e9czvBiMzS4XC1WFIvEjH6+x0yJacd+yRNk26FVEUVtlqBpHWEE4UIDTiWp
7Qb8vJzKfSrK5uGdZ5pMlJeBmcbXeNHZD7Acezj1RGiYdDdjXZkWCJW0qn6bZPBE7UVqrFF8q34C
rhAGlJCV1jy5aSZtgYFnq1FOZmsxdZ5zkAp/k0fNWnqT5tD8kLSO4Oj6U3mBx4h1fdQYAV4cxzpm
VlMLMiZI6kDF32k3sszWn2gO0ccIbkFBDULdMQPPUi7zCsOX6c9Qs9WqyVN2NvXSu8YImbeW1yAq
JQTkcCBaNJ+a5Mmls1WfGZ+qWh0xVpI2EByLwS7MG6aLs1s/VIyc7n5vPEiQqLx3XtGfkLDYNNM0
+4xT3BZwDKuH7RnL846NewMB8b+ZEo6CvtModKrbSJrWxZaP8AJtxvvxGv1zjh0z7AExE9937Dax
PISNtgh5GxTLGcuOfC/ChuJ7d5+vACRqi2BTNRa/u9mg3zdhcUVobjFSkmcFCPjOu5FU3DhGldwE
cJBtqx0Ktrk3n0sijdifSNJFdYYDYjpJcWRDslAM3vB4qn99hBQQl7ChZ9quu+IJKox5PHXDWm2p
3ScD1OHl82aNa9m4qSQggOV5fqvAXtZYUhlJvaTNnW5tp5TGQdHrLr4g9v3fLXlGvSbxFrysZbjO
tlaPxg6n2Koy1kNzKc8b7hHjEklS9RuECNA1/q7wab0rApY9UIdI09VQYKe9LJoF0wz2RLKiewAf
wCKaCbA5xfmJsmxnU/XmEMp9kdLZWsJqKa2G52YDHGbufQM4C4NSQ2OoaK5IJxtOV9q2+LORBBAN
zmdWN6KgLHwJT8PmWbaH6Q+aG9gdpL+PvbvMax9uDx0rQj6AbrXnHmMN90zb9FjdDFq4JCR9A/km
BApHzNXubrHTT2gQLtOuNp4zkyeJQKRvqvfuBmyGJmkZ2fGe9CLasMCittx8ZiQXNOjPsTRBUb2O
dOasvMfpiEj0oN+J7yfAx0/fjovAX8JspjQDcwXD5TSgRKMuCziHEmpBIXCf4CDb08KOHy2EKB/s
nASY0p7PFTeEx9Shlv2IBHrY8O/GDsB+Sk2/m+DytpLRjP7VZ1oAZFU8flSdPMsuWkCPubq3qaKu
W/Gs3GYCAov+PTNpJKmMxY/87i73UthnwUwNPLYp8YvO8lO5uJnXv68GNn4s5Z3Iq5qnZ67qBVCt
7ilt61gYRAal3g5KGVu8Dho4vUTxtcau7wVmHHSuSiaMP+bZc5cA483OlasORoTevyDzOqBzcAzJ
wtbMv58YFRwDVDWEU3Jpm5f0unNOUMdDSfeNk+0h9MUZE9obUvQ+CCbakD7b1h4UKrRwunXb2fxp
fcl2NaZIX7m054GFKvrv2zy6HVNczZ8I7lU3m+/ra6M0fYNwit9WBHRBKjmvSQZ4eCVtEZ29EPC9
hYLYQULqpuE7OxSsm1CqRyA7tSdJdN+ROWMFhEkQjQ1myav12hPj3Xuq5+6jt6t1S0l0JAcTrfLc
+7U83ZdPPpm+iyeWeZBOCLTFPyo6qN3p/3yk+m3HDAFf+qUB4iSDnhpNsXfPcBjOZXuCbtbicdW/
65hT+B7JC2qp3iTkapLSa9RTqo91wBAWaCUd9kXUaEJrVT/oi7YM8oC/02jUZoo6vwo0BtCu4JUc
ePPm9ybJlSqu28B5t2s1OfxezlmKo+cB/G+31FSPq2o0MELHEBQ41+h5VOyo24yagXWsu0//audY
QmIR8ztNCeESUlVLwFuI3JAaab9Y666LCwNTgZj3w7pkS0JiBgxSh/6drM1ZXPjoN5SBPLLgNHiG
JV7zI7uyd2UeKO2gUvul6fGMaZeiSzrnp4jlInYcyx24Xl0aaSrTDQ9+ZJHiz567X71wTDEboDH2
60Kbh2oBhGCSuV1GpaHW6Optxdeq9JpJKowLzBRAW1gMmJngEixHr9oxWQacT0iEXIsNuxl3avGV
g4kNFhQZxsY83K6V4WpI3wA30Xt1e0uyeQ6LLlyo29lNeVMUiqtJz/LmZHYeeDmE1RUMfkQVLnZM
EPe0/vEFNuAx01L9tRQA/0/m9hLtNmEaq5N+Fb9X1io4u/Brq7DJQYuF1Cfvlewqd5deWc9NkEqi
4rJ00tzJsnsiNSE1h5l8A2zzEi4yGX706UraiW/ZCyt6PizSjQ58N/NAJiGuBSnOehrPPzDU7pp8
qbOTltn82D2qNe/helvbISTUrok90/QzdRLrf2Lkoa+cHfcbtO3TS5I3JJmln2illv1XVprFC93x
h8V+9Pvu+z8t8krZs8qiHIQew97obVxLHJ/9vt/O/390fkzWDsXm4AgM+Vo4i2WYzQUzEadGWWzQ
QFfp8WgHhOYNx5rsfj/HosR2tbifxSxUcl6LywC1ApvO2WCBYJMrQ9HMKF7r8V3or+1M6j3Yh8S4
6sd/b/SmLAYQBiiTPsioqyPlq8r69MwqkSMrBnRvRhndxhZAaqGvAEGi6I060rmXOV4G0JHGlsRP
fMypQnlWktH9tH3KfzaEMfIz2eXU1G7Uf2tnhPkzz1RoenpFF1QR4pFJYU29kVUrp284yxOUamVI
Si/zW0M5jDkc5nccNDePZ3WJXJDrxM53aLMY5fUsv8xLI52xKKFXi5aS5rZiz7CK8pAkPRPldZeC
4jYuoMooYMJ+FfW+HK8IMSzzGJeSVZJWrqzRZskXzdQaq72OcfR2401pRrcvUbSFg3B7vtYOut+b
fOsxnTYPQl9Csn5HA1zuFLZWbEC+YY14ObXEytPq4C56HxGGuhctUOhvrtNSVTalWYrkWkin+TDv
3tWxlLktSWVY83tINTYqOA638O8DrWhl21gJ54AhiOHjX+SsE+cw8JGbZ+BZwVtkAa7rjfB8KaTV
NbGPFFKqr/gY4gr/ysjhdkyxc+37JIstPi57vL5MqGyQigeFZut8yeue3Cn6n9h8erqsrVkZeAOB
feuFRjtUTul3KMnlkzHVhvGf0RjdXOc3yYdyjY9eRpCrFhU4fUWP6zk8meWrm17nTBkcgjR6P6Xj
mV8aaypCBGkUnaM5KcUr/yfFTERg9+5wVh31aSpW3z6vCI2vgVqnlZ5NQqLdsvjT3kMSBlBg9HOr
L0rTnAu3FbNDkpL5bkkyLhe4pSSVVBMVlVtJFFei2zZDFZk3q1cjfYAVngZJP9YspPoIDM+tAek8
QPenU9F+2X0m6msx6z7brFCdd+dcaIxsYRiblf0TfX7dsz66BPpKHzVJ+6JKR8C6cMKdb2k2Kscm
KupTo+dXYS33hlStxeCw+X0JLLIWPYMsmtWbjEpLzOz1uOkQ6AsCCUgaOtDvBzRGr15IBrTYNJLR
IOVEHuWzjzSW1FgaTbjYZ3x+NSWTMRoBr0UccpLT5qQ5xE97xq+MG8XmJFxHtemA7pisHUvRIzz5
TfptY0OjUIJbyK/jPP3ZNlooZOruTFkeqH/JLdmZuilKpFr7Vdas72zAd3F4UJKpkFy2A3vTEI42
W2uuyhwwluH/16X1BOoUCNxCbE3dCrnpaY4GN0tqhcns0NdCH3VkqznN0YCFygV7ibIPkQtKOeBv
tGnf8PUp+TdKEPII+8rW87e/il1/TUwZyQYZ+d8HlNOdCLtiqi0bCMr/KFIjngw7VjaB22lmFypL
PC5Ae9ZSkq+QSxiu1/gRYciUyGetDxqFU75tOuB8U7s3J17SSCPj/zudqz25wKsVFec7Hxcl7O36
HbneiPF2aqiOqtIUVV6KzIm0zu5L4ka4J9Ffv8dLVlW2NKMLgqRW8KKPBOujwWjMDMxCtcKK94an
fwRceuHn24NbmzCGfaOBwOlPQqow5HlDEYkVoduCY6zwmcs0iLW7K6OVJsvXjemW4OWy7YrHwQFM
/s3HPJH4Y4iQKhIZKk5AmbdocYxyNpuGHZa8f6C2tbgm+lXwAfQLo2QHYLzQvpaqVgemUDRW48Dp
eyHxoznSCB8/U/1TLde3rz/3nZChkqzvxX5H1LYcp/mqzA8qOzdMZZ4bHdVErqAiP6XzEK6C2hLp
rweFSjbhhC/Q/IVSyHFnLeeAZclNi4q/p/8zvaaoQukpULvoKm9UOANqGQNwwLo6XIAF8wgx3ibg
n8322Z5YX5SJL0c86c3R3EaebYio8VGpQnCMsJqg8zdyYGEmkUKRqS8aPgf8Otl3O9Fzd1Y7MLgi
lS3oiLXEK/qFWfpad5ppjUho+sfZMDDXOz4BAXQ07LoKA8eM2PP56k68k5NP5DFvH8yL8C5ai72o
hHdmlvhvUnxTvXlDqdT0zPpEz2zR612ZQ5StWgQ8Vo8ioRO5nQEwiX2Kuhr07Q17rt0fYZdCNxXI
DmEvt7tH5JHSoMy2KF7N26Ty2hwGaI8FTzM9tDl5kwAIR9zB2peUv+/Ecr5ya24WygRpbIzkOQxL
gW41XjzphqXHFBjNQEMUd2Rf3tEsjMSGtNHchNR47cyKe+8413aVYi8bJs9mtcfUpay0zQnxSccT
t3NDgJo4z561/2E03vB5r6TpBHKQunzIzyADL+gJ7oHLy7IN3FXsVJ8jyW/TrhPMKr0g03RPr8U6
LC1ZPtGff9i23BB+rFfi0ECkfrJO9xf1DQbqeiW0osWvhpqe7NJKjhLPuQnCmYRL62c7sEVzNsxi
18+EypzeBRVe96W7dzbYjWSjj6vWFPtvAiGgLoB7wqmC/1VOx/Ab3Zvm9MRJcK0JFPADZ3phAAIA
/6AFt16P7PdmF8yfS6FYJOp0pZMtZK8nTbBZYNgnO8iFkgDunO4IiEqIDloGxueOJHpc+rYI7+90
nY0Bd0wrsxVz7SSnG7FuGaEe4zTUbnX47DIGzgl8Z47mzuOIPfjWA6OHy2FbtQZrJK7pThG1byyj
dzBPNYS3rKAcSE5o32QCn693PT1zSEW8aud5TaAPJZGCoL8pf2acNthbkvZFL79PZu25Aho/EFCE
7m1l65/nL2XOY3NFHP0oKROMYtuHvzLw8ZaNXVbPF9y1kGVzjXxENfNDaJ/+eFzyKsfJ67aU2/TB
rddrZ6F7xjNTQOlkyoylsKyG04Vf8Z7Jot/mChTs2U8X2/CD/KoObuNITd1hNBLDzST1HrmsagCa
UK0RFUtf73IzWeDFK6xElaAmiTFjSSIKRvNJEc4mmKZDsYeQNcrcu6dOe6c/7VX84q5KvbTx6yB+
nWRsbSvTWQ91VN0oPY1VtFk9QF+Lpnf9dPeUOARCV8FhSMgU6T/cGvwC3afr3Eh0fxHPn1ezaW8P
Hy5x/Udpmi+18C0ZD3vxUWn0QNruG51rA3Jb6FoXR0TXP9N29O46E2HGLLAlZOEmy2gpc6E5BgO8
AhUUe+ryTZAImQkzmhFqO0HCurVLmUgrRIOOsLrWNMoLiY9cn5CcrEGz9RFhWyaXnnskLlJYH9er
xuB0qG+3iqDk2SkA1AsQfb+q5VuhAQRM6CYAyYM7V2D2FEqzr7hcVD6YQSPvjUl6TyvBRfHqTBTz
k103q8LB8u8ufub2Bcn0DtvG4Y2n2sQAJFkb9FfAJ+NX0KDYTUwN9miQNGK6O1Zue19IppMRPbdL
rs6BVR6BmSlbNtqgsssZhDIrHKBiNY/VRauVH6gN51U5gy+21zlVb0MOMWiKKJ+Fl4hZTdJ7cQnI
dP/xc+c/b5jOcYSF9j0Na9u9mjSdijnm4gPf5CRZgJl24pCvqxjbQfHoFHXdDdbVkKnZY0OvOyjv
NoI5r4mxqgudOaWknujeX1a8/zEuwls2FP0pK5tMhJ7r+bxvEq61ktMWcRV4gjpYjFGcC+xL5I+n
J9itShf1EwTXduNR7Hci5OdUq5uprRXuQpxJn/vMe6MTO8PvzINow/Mw6QtgLrA+SecdD5csvTHZ
2qM1Tn/IBiV8o99yWOlES6Ij0mjxet5v99jsx6gfraBBxMnEE8gC9Dr9mRMo8B+bivTCoFotIEED
cW8n9WwLvNpkJr+nDaEjjTmjCk57soMmh4Lj46pzI2ITEukX4Uwo19KZR/xo1Ju8WAkFaTorMlbb
nVW7JpzulJjaSQNqrGwfi8q2LKOH+l2s9ooysTjCM2xJEFB+4dyozc2ebUVIgnGHwrgTRl/MYE7D
Skm0MB6veXu6RtuPJsXMg4f0qznuxdcO3OO8RZALThb+mYySdST7iY7Dz65hsMGGi8TNs7vaXm7k
vmmo9zZNOsrLZpdTDgJBUEubjMzq8VsO9cB/EN3Th5yO43cQK4DeDvhJAnWdmPTIT1XIU8os/00G
j8Akc/IFTEVzTpAqc1U9i68YNqF6YN84LAezxb0gHIKJPFEqK/5BFKuKwH73g7yHy6Nrjh8/4uei
82xkaQxvV+e9zFBKYn8LYzbX0fKsH037ktHqelEKENe9AchDL6+IYu/Xg/X5zIhB96LRNwL5j7ZL
ag0VHEnIOSGRn4Kw1L1GwlwvMIWjtLlbJ5eFhvu+oIf/5wwX4WCzEgub80KQdeI8fhgisrJOqRYn
8qDNNdhzm6BsCI9y4ysZf83OUGl7icMfUqJGtCYtUwZQJudbzN6ndHan8l6SC3V19g02HFiB3HDp
RVn2hMqftDKxwiJr+/e2xZnXGIcBTTjX93fS+5xjcP/w8Xvs2Jh0p3NBuX00CTXGHrmb/mR+51lk
01TAcp1F2AFHqUXlQ8xVrDt+GAT/z5vyvPjt5BhDhRt+4GjvrGCryBV7m+L6YLbPSi4wILIq/x7K
fclAjyXAb+QKO82kyL5DNG2SxVoGrPT0scd4bmRyH5ZmnP7vsNUfBm4EvNNAY4uamRlzUqvK5AfN
AEQv9GxSK5B5+rEO/hJwOyzFu/HHDAAiXc8h6jTJ/IJvAMttqcEagJE0ZKLGlnDnnHy6gtdRBda2
llHPbgeG+/s6xT38JsvFaxWKPcxKjQM/iBYtFvwUR3477nGCOqhA5Meb3XTdmfFgtFi78CHrmSxq
Y/VB9cvscgz+CelxH8JJCruFx4N3C2YdCKDvYIZsS+Fw1j3JJOrmAUxu62CvoRGmN+NQY1FbJh7f
PY2NXF3HZvUIS/22ZvBma23KVw8JZFYud1N4WFTBq+0tCOyvIOZDNg/yX0PyiFN+MHX0zKXpgOH+
wO4jh4kaU7ug5nEFI0znOEXWZ5lj9F1y5YpGh9cT44dieQWOnjjko/vF+5pubkpDkSgf3LXrPpRv
vtAJZ48inQ0a+cjSGzhfaDM1sdY4Ms3bnVsJoLS2PzJ4xKCH+4YtVrsmH/QQgDWixwntKT3vJQDL
JKroXBnzHuRoB3MxOmJ91JmKDiUMtD2Vzp5OYvft9TilnUemnZH0q6v+uSdZbRVxq/REh6n8VmR3
dmcWYuFksL8fIhCEhxy5vCxCe42BFePr5IqR2Q9dgHNTQVQErGOUH5D2s/wqWS4woMN0ER0ysMGX
OwO5NwEnjpWfzGUXufeX8ogkd0AxXZ5iaJY9w68gBjTr1h8n+crIVttxIo65N+eswiXqwjl25zfE
2JHF1LxaPq4YgFbWRivjPggwkHYkDeMXBJhAH0VEBPRfuPr8FwtT0oahwQ8F/dgnws1xT0lRHchs
4RpI6MKN+2EFCUiGGOfMVfBj5edKWjF2oSqlEIokg5G1sTf0nCT9516NShfiNkQH+51u5CSWVqvQ
OeopRjpFgQ/efGwDjt4swQwDkQNHh6FUl4+rBogsmFPDYYXgI7pkbSZuDJY5jZpeqY47lp9TdiZU
L3OpyZqZwdTm+w6oCCV4l22fj/rIlB04iXnTxHnDyVeGceeeIjLd7iFhrvi06ivCRSfPmRiWkVg/
a57LV6+RA1JR9/9v2PVEFwFoNTpKv0Qy0yxT+F16y2TdXyvCMsIouTTvN0mrGIMg0UJgErYDGyPY
tfrcwKMZYNh/SCWQUs42yyCElrzLHi5i82EZpv9iV4LYGqAT+Xed3o9+IDxPpMWj14QmOoH1MPQ2
vKw5M0EmpU44hM//pOdRAiEHelqgSLmnx9Rh6cwjkSTh6xaeWrLU/i2oO2X/z7DBuA+kEP1QbvL1
mpQv4uTI7v5XrHSumgBxJls7r0Ij70sx9z/+Mrob4u+x41LUmGuigKAXrZY4pB9ZyV1ZSY9KSfn0
qboAKIyNTtzQ8yP8q1f2XwgUTO6lWIvV6ilRAAmNQOniBv619RZ2iAiMnTC9cHyMGwbkgFd2W4ap
0gje1FiE4mQq4ni9kvVhajywdTbmKYKDp2tly8JIBubIW8m4jp9si+FBvf6BqD08GLSk3mGV0Zfo
IENATHqLIWCB4LV5xqlhHKesmSd8wbGITf+RDkxDqAMBq3uFDBfSDBtVRzWJTbaHvfbIDhbMY+JJ
+5Z7whinywidpdm4IxhSUvSsNnQIs56ncDEsGJ7im9BfUaXQ0mEFEIpwWMlAb/qtLDa+5EOMyfYA
ly3nrsS0mv7nAba96+Ur1J/F1xpezdAzTlIiDFAn+Y7wuFhqSlaVBrs8dIi4rzB5I562xbXNtGXl
+aHWNjUK2P3AA1njU50tGZIBouNM6sJPRFyFDPZqXmssHS5fhvA6gBsTG6l1cXidURoa9s46x71a
VgOiY0UF80HkqegMHWXfAqIg4SadBRbkNObM6J6BWuw7j+F/WOOV1AQ7JZ4FNRo/6tlAup4PPEeo
YycECRblJe2CZUMZimrFa08IvmNEi9RzqvpYdoOpaSGsbD0+11S0ZLcnlG9/IJ7H+NtYatKfiZyf
YINrs5UtkXsWWTKJ0AJdbaOIIJk85d+qIz7OZyuIwm84DG+g7rzdpyYijCX3RszDfFL0CVGXF5VS
0YRgp8LUzMO8Es3Kv7qdsA9CtceDSPtwhzz4Lz5fpo74ZWpzVnWtBLkzgsciYRM8R7ZHbTFlv279
KPDUBIr/on7a9PcJYTYRdpxBdW+x5bN8Or8n4nqbGqSdS8C74hui8MyCGPOR02oFzVSU7ukrt977
9dH+RKn/DeCfPUKqtaJkhL7snT3lxjhOpnLdL0z+fbWrAgb8iPOHkaEdTzp2/ugZDG1yh6V2ExSm
tsQoyUEXx+hskH/3fU/+ksHuRjFjZZZr6rJjr9szfOyHyOOz2m8oFlHY/XtTa+8ocu/PObvZMEUj
h0tALYnP8KH4gUal5JVjIm5wQMDh/i6BpV/kRfFB01rLp2CsYdwGiMJiATkq2bwyd/XX3xYmdKhf
MHxXRnttIBtmJqGjMRgdKpM8+jHSpXwtUx1glfH1wJw+4TLZKZTQyDQkwTbAIZF9/KDuHslQXoYB
n3veWHuln/5yGX2bRJVtNYzKJt6it/9y8NGEGpGxGr495XTLHRZ14mPGKJq/kqFGGvkWagMUqHgc
8wTu7RSqutnQe7+PWaZq0iIcrZZnNjd21Eiv3819Mcmmx9hgKpI9gk4Vfr5deYuYvkxxXSziIUal
Kxq18BLGari1gHE+NPur6+5+PwEH1Ucx2b1E2H6UOgHSJE5ysV+daQoi3QVN3YlvNEfsbeqiSE3a
yFy4okeNFKdeJxr60D5xOHGnLvVcZudLBnaOJBXclETbH3we5MHxptwO5tvyeZJpByd7nwvDhoXb
olr9krfoql/ahsZNrO6IGBOZ8YWm7Cz7/JJyjbpxKklT1M0isPUGFHczVujE0ENUUT+dYKbMWdb/
oqHjDPT9U84enN85JRet09C7DXBZ5P6QDHoCNlcHBPm2LxtpchzVI7lttVeVkxA3y5i08DPbHmKF
ROO3Yf/izIC3mPKARk7xtCRYaKqqOH9m9Y/5dHqmCyHg8UZ5fZSnyjy3KUm8KBD8qhqxmYxjR0jm
UGq+JTu5LCcyZYH9fS+0tyz83vL2w3osoR+cEHA2Oqm7a+6RWnzRDWEv+FtbZxvS8x669DJ3sZJC
2loJlluWu7s4axKGtktFiWkRiralYeUWGgrVrnrK44CpAJclZN+h1sqEop+cNP3OnCIAlsrUAW90
dDjJjysGBEefFxFGRcAo0snS3kFfHUpo4UxEBc2WpXREC5yfqk8pr1XFDSxB+7H5xcLB7PuB3ghw
VMtEm/drDUeANcMEDet+6UvdQzMnz6Aby9pv7Kz0EJfPJNy8p5Bdj93X5bMsu4W7stkvvNZf8b+U
axRZOQfCRRVo1iaCOpOZLOrakKeXd0s7mC9ZuqeZjjEZ+YeckrQ7+MTESe0Yu1+ffOqWgqymG8ko
C9DAPUdUvSNnfM8d5nMtX+FpDkRORGForaGBgyBIepUsaCMtsoUoSwIfnH+aP1QDzAIjZ7kaA6mi
hxprp0hrbS7ZcBbEhAWrNaErLM/RAzRFhIMkah4n/LtCk00Cu4h9elybTcC9YgvfLQFdmhNOfwc+
RU3Vgrr6sd0WxR9/Ng2/H88/RAIKpKpZ/mejbKD1dsNzMqI45CMN00P+KIefk6jVwUrAijpqeZAs
eBzV1TbNCQVsD53DW2qjHEt5/5dora4aqR+fXv9oaqdKmN3ChKwS9upwsAuQXE7b2ScyNVOp0Plv
HOPGVcBLVGz/a+6VUhduDKS4LUDH5zb19Dg63PNH3OqMe2eJ/glbtLitWTYS+PT54Pt+ThlP56Pv
Itqif2nsPN4vY4BtYRbWQMhVfSmhNkKLXycR29xqcrUH9Npg6VQkEEBXgzh95cn7SK6Im7aq4ghL
Sppi+zpZQNM4fuCw+RMPV6X4EJjXvyuK1uw20eN96ggYc2Fs7vqdVdfqQL9zidMwbJGQ+kurE80J
62HQaGhZiWzlsrU4MQHyCxqYApczWUdqCifroo9I8CQ1tCM5xwK1sCUUqE0pW31xXNTl27GnwGoE
lwlf/I3bJGPGka8jzh6w4qzgj72f0B7XoEXwCHtS0EV5ptoX0pbaAxhfwbptgLOFn2jV8vpJrG2w
/cBmQAHFk7x1Q3h+jfb7xKbJj6An/+AGzLgwnCD8MDkKGL+nLIKoWRlbMh9TsJIdFjqJMdg6d/E/
UEpv0lhz7ak9Q4yrMWwMVfzMyPeFS82rE0m2TD3e9WYEzRmauJePVisWwxA+6eCeOSNTjomoVTac
vwkbEYFtyaXLIApz2soOEdCTJ8aspkvGEa0u5XSizUCbypiJJM7M/Z7L7xhAg9Lw3uPsIiklFeUB
H6SDLmCZLQenrkp27hcCUBFMKyWzzppW/4UXkYcCxWx+7Nx5VMz8ruKJUBk6D1YOar0wkOOQqRqa
7gGjBH2Nlk/J5TL2hmBsn6ZNWPw02VTtWsOad1f45gXj57gXyqTHxnXli21dizmg9rrnNNUy+okW
J09+EFY0SJ2n0+k6HfIQbxdgWIhsjspCDrwM0OkeUKlyxIsDRe8MSt4W5BtcfTPKcuPsnV7hCYmw
VpSQiGKKEFhF3L0VErGAklGq89qQUpVUswF7IedJ5qFLc9vZsyJ1MFSW/x7WWI+S4apmkUHgRdwC
kwSlooN6wrK2WNNZ1L+iIxpezic1Z7TQ9btNkQ/7JY71aOGyJZb4b5HUKjXWL3a0gbMKbNfz4BBI
p66EcIbxpIvZTOyKtQTsYXDUeMBd+pPxehM6v9SUI0IfV89mTrlSTE1uzDSAoseIenIReTDgtPMt
yTk9tEYqAVvPI+EQixgb5o+DiUgtuz3IMV+MhD3/lzpCyN+7GKnQN8nc2VWobAE9Y/3H9xSx9DP6
mSZDtQMSjnInAwJk7bz5qpT0n6plwTB1pFsvrdHTWm11mTi6CU2KSzQs1aB5raOcLYP2Y/l8NHFo
MYMAAI31StydkKroBh+Yhggpx3IFC1+SH8qI+R7sQIl1u6Pyj1CYih65C3i85WDqhyWvIixCGMgd
cmTgIFkKxv2MFYLyrnsLnS/nMBvtC+aNuVyy2z9L/zunneOm8Q/xuNQPtMZxqzV33oo3EFtx1FNG
clWuBMkVknL6btlmANKTHCC+HdXRpVlTaf5Gz42XLJP9xJAgWf+84APQEhs0npaHDE1p7PeUJAHx
M9/3IZsDkE6z67hqbj5kECWmex5rMoZz2auCc9o5U96diHHp4N2rHKw2HExebNNkoMb6yZW/rPtu
i09PyLOW8+CJd+0Dozaa/PFHWUCakGts+/HyjrkxDIaZyS992i/OFTfC05lkqIogDxC3crBd6A8R
AT5sKp6wp/XS07x51mc7V6yv/oO9/CIndghwmlSOuMMkOI3OIcel6aP86kaMliwNF79CJE7cOkt9
mURg6iO11sDv2EoEu4DW2g5imr7zBj5nZTH5fbw1zUfjgEan/+SkCfbPxJ9NntTSzKO5ZfWd1QG4
M9TEid/C6XfJ0++FIkgd5Vrny+X4Pzw471XtKrLu5eLTXW41xkqvt1RKZsK/gzYAksFU2Bu8wMnY
auLvuHA4Pi6Px4zEl53fjOYNgGdEeQkUe+BT719YMRDWEahzOLDYTsx4UiaC5jpjuh9D303jupVt
N7M0gwYMlb9eFxSXotdJeK+U9aqd3+j5v2Hz03EgrqMGZ55D64krbz7w8FC+3SVe81ovVWJRckTZ
3Qd0IgzckoWmLn7L3RJwhDAFz2yI0Rb64gVi4E9RRWI/KjoDftlQCaUL+Ll3rEAsRANPFlN2Gby4
R+ZoQ9wEpRCJItstRR6KUAl0cPKrrXEcq2IWk/dQ2Raf5b2OuEMPTDqrGGLTWc2yIB45R5OBrD/g
DBFpjra/zCxHkqtyJReUSQORGWnPkeBSD60pVzFtHJUvDCR3Q6jRkv0cQzYZN1domiP7554uzQiY
yCLDBmBqamY4naVS0fqXZICdI1S+jwCNALG9zxEsai78rjUZnetMJprxuVmHT7Sh+KH+S6G+T/R4
9hePPd5enW3xXTeC+YBDiL0ExcyaTvhwFploItrGikiM6CNknII5v4Mqy4UBXHCD+TP14SMsLGTI
bdunKj5+L49w/+zLcDfdQrU8TsQMVeX7rcoFpRIhVdwLfhjctUbAjYb7XYekv94TzwZq9QDTVpd6
uWiPZopFsCLTWYi7BAcnfjOLlfusauw/JLmIBiEU7KXXlnB2+NNysBoALr/eWv2AmgQ4M+eMsg/W
wr4Gn0Nyb+JeG3MnOSoZ/vaCtMp67UC3YvoguIVqCnLbbwoeRXoAWcasNlnRC3MgM5iyneWDoxcU
+wJ4DF7j5prokQmnhlayVjO2ksUxtG/6LVX1ycTMYyMb/13EKLpB0LovC+BMCsTBpfXv4KzQCtNg
pR+BMgJc9f+2YD4/vj4fcHit0ON22eanQaVDLziiLCtv7FpfQAYPEvmZ9RlW2MfMtRvTNIeuKv5V
qgFojWYdzAMeUXOATr755C97Go5YbmbdDrlgzF8yyHucsFLAeDK2mmUs78Od6nl4kW0bWBiXc+Bb
BJypcTDI4ekm2Cb9UAHugO3fHEVeCWAJQjFX4tkOJmKqw4UoKzFLlAcVrhofY8t24ruGEy5ngm4b
9P89UsQTg8geGNCYY3g0JwOkpblltKFS7YMZiY+MMiwXLcyteHLyB5e2Pn3OASqjsGsJ+Yh2Ydor
aA3iNMIM799l64HvMWhwgqpvuHMw+uUK6g0Gwd8M2HWa4a6RDXfhjXAMtMvh11wPhJkOcT+pKw07
NOA+MP2t5GRq9cgb9zU3nbwtAJDRLmvo1t1jLGc98+wC4rGzZda3apOIovl508P4V79PZDW08WH9
T8oWNehDMXsonhYbr85m9dJyXKKHK/zPFCjtMhCIEDEabvBx/XP9PDsXuUxcgFMHBCRnWrGVmdBR
UPvPTpMkLcTr+qm5PUNtSlj1J64fTWMWJf/zbDcZq6aEja7eVw46RP8grwzywIlxESQWlU2ko70V
zqvgkmQa3PlkhgelKQSzCRjuPJX144BGGxuLlv8R0Rg78BpNdfVA6S3HaowEOUY4PQqorPkgmPFm
8uNZPwheUkwt9XakoI0N9ccmOluZ45l8m9pb7i7rv9Mj4Ip2uqk8Tzohy3F+mrFez32xk8yCfsEl
M2zMk20BM2qqb9CZo4rOtZlkcbGcJfZySD0jgO55DQ5bAmEqMtwiS2XmE1CZDMzHToRb6UyDXCAL
v2SR7m7iG+86+/7ZVXx+xoq+nswyIvB0CjOviLkyBUCQF4jRlN1VRc/LQzVGr5e7PUdPN0MDeWNj
cpJJVz5CMoPlbRYiYCfXKzno9wq3LkTliAMrQCN5gTuNhFyDwE6lA2zzY0Gctn/bnSfbKhnW0Khi
w2ZrN0RTZiNU3QHESytdh99xeKyeXBPAEZIgL7w0c5UyguK1cF9hVfhCFofHyK7ntJcBPa+Yn0qS
ld/ZkBXk3APJTm2OFXBka4i4swzKG73M8P2NKwcaUbOAp6Dwn466ObRcGp2S9a+4Tn3ll7d7caIR
VCdtXAHa4JeCvZBhhlN8PfG9pXMvelG9ld8Hs2iRcn+GE/P2b+X+BQviK6ck46JaXXmZ1djsrBfk
26Dq3zQ3x6yrIfu9WkdRl+pncRcqFwHb90ZsampAixzBuzPQDkTpWVyuIhJ17DyfaBQh3oVF1WBh
cTso0blKgBFW/VbiK7wgzOfaSVGMwIK+7Agmwf3cELZD/zuKBgyO8yt+vzO7dmBdZq+REx080AVE
UVb1nDWCwqXO2q8ddh0sqNwpRGp2r+3oBsAuyVP7YwLKBZycZAmZMlFhxBkVuwry5gyzrNoXBSKE
3HrR6ve6bSqiF5hbzW6XthRVnCI3Xbm+63VxqunfwaaI0MatGOvdgGUGAYjVYik53u7U/EfDgJHj
QRD1BILufKEbyvV99NlxFzpN3JdQn2qHqm1k3JG3YeRAmuwelJyLB2a7Xy1uPFdBVt1QtLJfsXfw
pd3fHoOvqKgGfytqy338DHRBMw9yBxAXNfxINfc1BOC0M+L0hh4+ocF/2O+AQ8AgBTOo2fxaf7Si
mpJ+biEujjEQ/hh0HsrkUZiaPCuB1Qb2Cyx4d3FCEI7AUgg1r5lvNqN0vmp4dxMIic1XmkYgbp4C
p3SOJ03S5+V2rs+epwndoYM6IAtL3fXRSaorvNKq2pdtJ3/6ifxq+GRM0aYxeZ76I4N6l1troBkg
txGL5UMfFwK6AL/1fVhGDfMGjKF4cHlQN0ixSpfbylHUJg7W67oRCbAv8TX+TOKDUSuC9Vfgdq9m
/Zd1lgyd4DOYP73bAwwTrxlPesEXgeWgOppDfq5Kgc3iVdtH4rYXn/uxHMjZXvh/d4RzhQY9BoOZ
pIYXrOOqKXIsZf4YxcVQC9mggpnsOLW6A+eiN0GzgEUniCUnGwQVD8W/nbhibzoVcgwFftAKMwhW
FsnhwQete2ZWKzgIP6A+BWYzh+Frgtm0qeSBDrRJdCMEO8jqbQw8osDhdZNBdces340gPWHMbIg5
qJZXr2vELWBOCLic3V+r8TvcpJilZ/k0+38r7HDywTNMw8jU4hvl6WjJgb317pgQIt/rfB/ZnNoG
GsIJDfGrTE/WjFb0sciI8C7VM1zKHHbgqruCbS3swJ4/skUBMv6iNiLl5MjkdYHiJTk5sZ2phER9
OAOzDCOeWOUl+xocNrhiZKVme3KP9y0RVqqEdlK4n774Y5AlfyCw4Bfaodyduuq9ABV0VDZB3jv/
O5Hecr4oixnwHARmyW5CiMHvK+AR4DmHEsExsXs8EMvgN697yfNtCBfRjdlI71Jzaz1S3vJHKU+N
TLdvLnKDFQUKK/RmX+wSEQeIr/5CzIetCoKAo1pHf/LXgwuZNuRGJSIRHG78opXS36+C9mFLzfpF
Te6c5XI6B2cac9QdyzdFMF376DX3JWMcP2vbXtV8yN5eiHNx80bwKInMoODp8Omckz7ng0Y5nRs9
/ES9qPxBkMnGR+XmvkpBI5JhbxPoR4ufDHfFrttL9Fvd6NPBJvrCOdVYpMniafik9r0UIoA6k+JZ
l+bWLNBkVEtq6j4kvT7vp5Ofa3ZgY0VFAr4iyctc+BB3GuzXC83TpSYBUY9K3r8KDYweZm0P9ZRp
OrfFF6/H2H6aljd/f5Cs4sYO2WSuNdWK7uMeBxXZIDzoCd5byhwOYHno9Si4dJyyvNZnNF93iRy+
ZJaAeoQsSEZqAV0yHvVqqQw+0hbem0tWtG9j3e2p0poXrFVMHvH4xB0xqwhLc73BJ7uflv/zxoo2
Qx6zFpoeF6rV8NsZlrnR5u5wPfrIPk3OGahR5eW/qF/b9K6vycTLVQPhm4J/InONcHN8/T8xiO62
X3Por7YfxwmC7X7znOmhtEe0CcbiBT0MaYTK4YsPTvCiZZBjSzj+hlgYrN8NzAEqWWOZFusAcIPJ
1UXaIMLbhDRkwBhw+Vtbq/aPDjPhwb5jgq4pOA57sxqhzijiKSSDNoj2ZCGo96uO9uoAq3HkjpY+
F+hK/eJpfTFL241HVbdTws/vFoR3icBeob3yoQQXcOiDwaaIOz324LQGK6BT0x9EQ7duxGp+ja5i
/SQhhhCmrrKy1sCxklBnbKUOr/stP+lGLw2GmTX+LgqwTPeDaE9ZHbC6K2dY9Nw7DHu04S/pBEsQ
UDfzYJsrcfftFrp99/v9YDmsS+5p3mN4FlgqTQ4TwFmGSwzYF/aAri1Dza/4cZOt99PFz0FqZbbl
4GtAJWWau7/304FXr1frXpUBk8yGA7Do+QMwoBTg1fnVn+NNnvdkwarTcNuQA8nVKdVefLvv2guX
91/1BhSbq/lOUjtxiKc6PZCFfYSm6tFBI2Xwcrie7lsXV9NOWlG6zkFU41dnjE8MbGfKUY0kbWyh
AVMGASp8O7aQnJXVR5LWyjStmlkSdOXv6BWBMlNj0Q+KsNs/J/SwRJ1oP5zQ+8/gEuZW/SjXcU21
/nqdqMaY+tMkxdR3UJccZkxBPekc8x++lSewDjvbR7nE+neHt77sRyv5YaQt1vQZH3FxA09o2Eaw
48cYhIoTh80nt7VlOYga2yFEhgwNwY2LgG8ZZUkmbGb/hIuqFclRy4d/9lj0anLCgTqbFtSmqsxO
IfJ74/nIs0u/J6RAhRPUFFZxsPPJdNT7+DdTZnv4gJ0jc2cOKO4eNj930R1pfTytDZs7P0YJK6fp
uzlwFfyR6q+H1DAHUtJ+tLX4nfY7W2srxHyk52JDzvdxXO4biE5+q5LDZIp9/q3wfZqheFobMtav
gnf84rXJ9y3l7B2Nbhn0Tjvxg3HTKFj9HYbQnzBzkd3qwCre1C9VJZOVUUX86tp19lwThsdI6HoO
oOFTRiRwwQuEzBu7lQ5kpmwrhFHmJotki556r+2LjnYybHPHjLBNfwGnDEgMfwqHwOCx6IPEJF23
O/qsCbQIDvliJNN+hZRze3VcgZHWJYTQq3ThlMvgUPu4oqekGLR7Kf/11DGifCy5ENR9hqSIFKRr
C46Zez2H7h8HmQv+iSHZwKbeSbw4krjjI+It3pzCJb/bCUym3ijtw8HuQvLuYLpUhQdoSAYgTp44
pNiGYHN3FYMM74A2H6ekxfvZjtadIfWCmD+YY4EOlZgAcSwBWvrKVG0FDZ8BO3EAHVdt3l5iKuWs
WzKe3vZbTpUSkJJKifJxHLRws6HjWkSToXDj1OkHcGeZcGL88GGcKZmEFQ9Xjg/0ZuJg6oypTunB
kE3rvv8r9HwBQiRig99+0et89NS80t7Z+bKwHIOmf243UQYlioRyD85yqtKm++7xstLtwR0zvFpQ
YbgYWwFVwuynsPlFWv+0FjC94VCVmtoJ2ZH73UaIIJ/hOXDa5rM6Njp9k6qSMt5iLeGA8msTwnsx
H2O+NG3ygbsA+hLXIwrsy33yylqbLMtL01ZFvuPOP3XU6ORkH4d2ttohOPJ+zpd6dGWOmR1Qu5AQ
JLTcNB+cmdLe3VIeB/0LDYbNBS5rFwTfk3A1pPJqEwdD88V2gqsWNOH7Uda5fXLJd9dh3ERBeYfn
fAWEPTMSf48EBNxsEl4sukrvb/dJD3Y6TZojhHI0QIOxPv7vRkRjLMRIBZdI8/LPqaeuqVpUOuh2
Ofe1c+SYEaE18O88/VNIy35CWwUrovRxCgiQDmKulUCeydNowErc3rP2RdsBN8SN/T+V1e1e57KF
tenneICvnqIeI+mhFoqENn2kF7+1bDnRLTBCgDeqHRRgW+Tvz8CeTYljz/tzXV9T/IdqAyL734EH
e8m1sHYfJ1d49RvgwTvRlqfVe0WiFAAeXJ92OhQjWMNwy64Lgt6jnalC5fBBVKGGbLzkLhCvRwjR
AURDSOqUBl9m34DH6pDf1u9aVNlLsIqxdGa4WNf/r7TRJEe7kTCxq5UDGtvVSDNizC7u4ubyoBSz
xHubFlxXnhy7hBsdu2SwJG7SNU5LXFEBUVHiqLyT8yEju2prfc6k7ODcGccjtYA2DUF8X1bfQHf8
uA0BHAll4G1Pod7TvJpu1NtYliv3MSydYAhy+50LXQzJLa8RHmNR50vxv3L7HJOyOcgxMIYWkUFU
fTIK44PMkJntnCUQIYDhJXj4yPdFwh+bz8IAVntBB3PC79yb2nDZehHK9d3lGq2pOAKhVUa/2eL9
yJoI5k5P0fRBNckUQlH5WgrcGmqwME2zhUgP7XdlShvhZYylW9X+VaN0RJqRb9za9mGYJ2Pg0S4L
GrU3/y7mTRMUStFyVepMRnRq5ODIyMXfA985QKmsf64BMiVQAQCFFJoMLr2gjz7xbD9k6RuRS489
5THYBgPlOVxD8bGKRhjzMgDDMt5ERUeVAo8kzDhBqfz6vrkhn4i/TevyKt/zTB+VboLtpk97QG0u
vDd99YhXFooW3m8c2z0v1q18e8k4yOUDCeALKMZgPcf0KOsAnzXaAG+Q7ArG2KYe/F6mf9gA3/b8
wA1Fy/W8ACKv5hSHCv0e/6WBnRvuEcFuHj3sN0nJFWRwxV0NLFOUdvQ59TDLxrKEW2pqPJo9vKOm
XCHK1ImR6Mi4najVxQxkckEhRCZVBaX4uCCn/c8IlaANCAYoQQIxt6M4i1zLbbiVM74XpxESBZwH
stLUeledeIk47ZtVVmGMCnrx3peDMgY+mjSl/iyBFDG8RIttc6a/Zi/LTUPynChyaENjX0Z8a+Mm
/rd9WN1eeFC5ioo2i7EZbD7qnc7/56HgBr9L+BcR4CegyWnjnyzM5ajVRinwGhyx0+UCcTsSbksu
8w4yMCTB+Dji8dfBkS+mnenXDu7o0a6eqDqSiEv8qjr+VqCHU4pat4TAqlHUFfIoGuYI7xQHHnDY
JhKVF56ktDX6Cj58uIObcDEp/ZaTDYM0hJPGeucBsYPZU8GTr0eByopuDR6+QFrarZawE4svJL9D
TYH1PzBNi4e84WgS7zuU+uj4ait4/rRpCC63NQjHBMzEJK5Pek2i+Sa7dBqOelfUx28WFZvfGJvc
KNJ1FAj4jb/5uQ9p+jqY/dSOPSsbNd59UPiv7IYDdPHRPDr4iW2y9+bHa4Xnx9H0rZAYBka4beeP
QeqDDR+lYwiJJpGEFSaf/PpCyrMIOehe/Hzj730SPN+RWbaWxH1rZDmJUYePwez3H0BPEZQC+ZMy
7fk3Z0M7/TkpGK9Y4S78IuHoYmvIXYeEbz8+gLB9SXLraAJsfdPLok019YKr4Jcf2dZz5iGR3Ksn
RqXvJVpPBbrfUENTv0IySv9c1vHUCJ1LK6yrdwlfRae8TC7klv9g8uiFhoE9qeatrhCoqhce0lxS
gV8njTP64f9B4P6pLJc/OhbXcqFJZ/ujR90kAYjUyTgafrdfHLdKJRwkccHkDJ3vyEPYqnd6r6i/
MeqU7lKamLbCJ52i9ZVpXq6C8JvsHdlCMfTlve2N1baapzWetKiDEhZEaEDQr6ANyZOvAWh6dubA
qwkeA8y+UcFQf7p62slEid/D7bfft0XDbBwnakkaUZLxAUVexDer1rglHf8B7ItumrhS9GzhEvI0
yjkfVw0/F5h3jx7GWhiw3w2ThK5VPZs83+jkucSj5hpxIBo56CFrlGdIsYY99IL7leG0mobM6DvQ
MhHHIMouUw/PC+RDA8lE4orTUyFDn3Q/hhvEHYp81YmKXtdGR0Lp7rs2h9WX2GZQT16UY5NgBSrp
vkKd6prC08G85lZk1nQA31+1EtKIBVe5MUJi5fEjSsIxshN8x7EfxiK64iwQZe9mwbmgUfsxeuyv
ysr6pY2m0678u0BMrBnx6sK2od1h60dMkfMIQ0TMIRVtkRlbJoZoN8g4IM1SGApS6GZyVReb/Z/U
ebHtqLFmLPFfYw+xeo7fWz0nJjNhsmU522MmpSCbq0PA4pOOwePOtblAgkgb1KvoqZ1f5wk0j1F9
uglu4B0ererxkyuYl6Cy53aFcE4u2HwWXEWSawyJb+OnaiZLPqGnM+LprJesjHZMvVGshEY5yH26
RhKFc+S7MgMcbuHsxotGNN176pNg+nmW8za1xQLYuObiMOO38hw/o4lQvbCJGSAFPY/r/M4Ru+8j
PQjgo8AgnGHCj4Z/hvVBGSO+dp3p1/3/7t0T1hIIO7GvIUPuVSdfTPepRDyEtXr0dBgj+c8yPwYT
402nUqIuNX9laefLtSxptusDPzVfGI2mboAI7Q02H6Ckxm+sPVO0GGVBu37VlVByu33hEuwYQNan
qQl32uPsQC/I6fYOOVt4/12NatdP84lpoL5j9dPaZOGyoS/Jl3Fnqal+QJ5jss1e9+pd9r28De1M
1dljzp8YNbVL7Qz4/SKpeS37fhct4oWA89eihwtCH11BzazAzOL3awEJpKEs66Cyx+8/5rmeu1yV
bk2LV/Jc+U9AuHhloRWDCFwYh8wJGMUiZ1tLas9DvucG2LqiKzl3ce/UGzqwdS9+mRDsEG8flyEw
ubCycd2HacsNdECvy9+sOzOlDVktHDz7rOg4DYa3wJFh35qS4NQdmBxmOg0Jdv+RADvlgGEOQciK
75Ds20XgJQEnxSaO54v0jtX+LQez/MKzpz0vzOdhP+Z4IS/Gz8oEYmqWGQPXTubIl+UEjDh45MvO
ASehJTRP63iGhfZBgiWlh4FHFAfW822wwSxpUUpHvi/A1jpukQg00qmfPf67RcDFHH2X0kK3+89k
l1SVI4KifH9y8gPhnfBaBqS43f+Ni3/4pnnyJfIbXKpUHTX5j4y9XBaks4QRzjPlrHZNOW/TFHN/
jmujdrcu8KEyobc/lvoW/1hIcRN0zNkNI8193hp+QnyZxWbapEaCJlirmyIos+VMvdJmpvJtxrQO
fKBYbYJF6iWsUybCXxbXL5t/eK7gLoo45jTkn66LS5nKJAzy8m/oXvH7+9NDOQwaA9hx5+337ds1
E7zXywjngC/7wZuDFO79hhKYkVDJuDW5Pya7jbyWByVlLyhIqSG4c3Jf4mCjzp4Q0TJW2vOLkkOe
ffU5LI69b8hgqklkg8w/MNvz+la1M5iKUqtJaV7XW1COaMZGlG4orzJxIA+8L5F/TpCdsOuZK8u9
dZlE9IGhIlaJ8bPh92imbKdsvYOnPwCAuEQfWx26pr+YzPj4VMeCk+4Xnvjjq3MqLhjtHEwFNqtS
1K3p8G8zFDXAGEYhHtLzTKvqX1urAHzPuOgJtT4lxEhaYqZ5sClUH0R62AjhhICr3hqV9eqO9Dbx
c11Uo54TjCaFFkZg+1NtG/HvBCCaED8vXxmGZNgNqQSpNEO8sNFafWPCjENNAu2zBZZk2U2QJVb8
46RjZcgJMsk+2QfsJDNg6m633B0gQGHuoxYB2aPSl+nM03YK8NRFRtm6CTbBJd96yeTNWXNmyRAK
RHLq//UQyxOJUYG1dju59Wxk1cHhvLK/Me7JAFxRj2Mxb9rOwaGoNlMLugurC6g8FYT7UfrsAhR8
ooM4dK8fYSEFLsL1utZxnxytUTjm3VhoZycqxaLq0X32tNIii/EciQwIWYyOKpCsU/XzDrZatSxv
PjXSoGNR4pdhfFEGY42iWJmra4oQIR4svpaVcz35Cx0ri8c/EEYAFCqJNtwnXjsTeLSEpwdZy4Iy
0uHbgCaiHFhATN64Ilth3tqCYM5u/7KbiuMYeYWa6P/GQ96fljqayjjwwTZJT2A8Q4PU07+jDP1P
SovMrDih6rs3q6EYjrmMmH3+SGc7NCk9tGAw7GBNVvD938ieUstIJk6wF83q1u0WP8iRhpEYGecj
U+O+4ucxoe/YFygag1UOzv/skcncbhHYDeze91iSr/URX80CrlPdHi/SIaMGCVtS8G5SaC7Jdb/8
V1JQruqT2XNF+QTvceHvhZrYwSrRDscejxChEtFQjIp3rjy/LL136Cxf1fqI6k/C3iZzIFZMZ4wM
+TACo4U43tq+1NT2Id1nUbXjPtelsEtw2lWqaT36Tiv9mzU196rdC8fn6Dp4NSFvU11qMjq6Nk3Q
oItXOXKSrTAdoob2xJcpu/IpBGfS/lybY0XqcFTnPg8s1EO4B3YckxiiQQSnfaM72LOx1KWlUxvF
/1REBYt59PTrGKmrCzSkP+4Jor52FKaBms4t1En7oTZ20Hyh3cb4EzdyQWSDefzG5c9iBsJtG/jt
wen1wNjEIdIA0XJcM/yusAWyvlZ4ZjPV73MvvhBusUxOrCFdE6pmsqUJNA2pcDfNh6asvJ/jorPK
CTnf/4mGcR/ZURq91uhQ5Wp7ZyLG4icsut7B0fdKxb+pDmsZf9U5qlB4llQ1qd6n6zmEyCcSSjmx
l7pfIpTh7sYvUQ5cKX6wFuyrXCCj/5DEIVCKQFWOPx0hC3dXvUOc9b6OfbLtTZw0MHLiNyVhTzld
4Q6LD/0R9z0JshWSeaif58+MiXLPeCHlsZkVxF7VpUZHZK30BKriNHfB9OGuISy/sAxe0S+bNkuB
PmrzlhxMZk4fK7GG2Vu6qoFZSqOVCCJON+fy8WBA//Ugkp3TfXRmPWzO+EYp59dEiY6XpmP8e6V3
O6Lp51+HzDR5eDvAMowpwjGCz4sV5s9ibC24ryebo++jtFb+2cPmmi4eE/IZMt21ZLffv3YpjcvC
9SMwPpDjNaNNDvbq/gx5Sjhw9Z1h2AuK7uVPVdANuU0ByqSydS52eI3KvirX+22J2axIVUZjay/J
7cQ/97dgRQqayaOtVhvmrD2T0rPgxz0fJe/UqxxFJlikS7knSktMH1qk2TIrJRTstLYsryVmNmXg
mN0NHsKP1bWpeAS5yXMEBMZE8UlpDWqXB6mKc97IFm3hYeXc0KAuSk2vS77ZEkNrA00BLP8F/lZv
ZWJ46VFHVWRBmnVEOBWxHg7GMJDhtymA5UA/6lccMfRnHWjmkZV5IaZ2+C3BbOhdIt0xRm/9+wcG
6PAODqdKys2PV4XS7VzqwxT+IFvVFt70bTEbhIR+xGwbMEUYL0D8YUBrgicyreblIfkTIAzIfx1P
zLcMw5I19oQXlkgcJP6wBQ6L+OFGnxEYUo8xiwhibY9NWkIJuiJzcG6fi/EIY5Fw1LarXjI7XF3B
SlO410kTJuwFwXlMV/b47ZNvOKB70+FP4MxMLGCagTXOEayTOGWJnXQVBpXeDw/r7j0ACW5Tpqdo
X0wdm40pnPCGlGo+xBgrhoYqFAIXKFf7Mn2NkDiYK7omzZzKYLvr98DAMVGCCHcSQ4CsmhnxOgKj
XIl/6GlIoDhdffQTYY22/jyFKSQmYym06stfpiiCD8wIHJ03AhoQYTOdkTStF/WEca0Ugi8UpEVT
mvpBg85pKwRH+gpTxSyVlBFsO+AMiTJyHBlcxLW9Yfdw71klVVfPpr+RNba7Mm+EdMHYoAYCVAbh
sqoOe4BK4pc/pd9pVeaVsbiprW2Y/wbHPQIsYrZpXtuyKO5BdVF1zBp/OJW6RPWgaxOF7SZ2PsH9
bZX+3xTfVaUYS+8D7MqnnvfLyDoeCE/KCyKW+Q05bhf/ChipRCszjfR0UloD++zIr1Suxpnf1Sxc
K9HiVvLzctKAT5TA+NlkNXbWREPN0eLJMRgGxKYp7+7e9d2UnA3BVcpCPwgw+1kGGwpVEBLw2JOX
o8WYg43U3kzhfrd7bIqDcXDXVAhzMdK3dk5YGmTju6u4XEqaMQlrvVtwxyphKAkP3iUq7Lus1yi/
59atj9KxjmPo/vURLi77hwjB/DsHbVqD1omRL3ZWgrLZmPuEM8zw7TTwnu+ynxahIWyyttVykPSI
q9wOLAso05iQW4krOV2nWA1HFApTDYt+WIc8fgF0X9axkXvEsu430h++GG8zVH7oJFH/yiAucge0
LOCXQ8RnnyNGZTFR1CRCBKFdsdUi7jBCYp9MFaxoxpWKrx9SOrCR7WxF5QACzuJlzunxs1qsHcwc
e3haVi65iSoFKHJ3/YBxMKYC6bz06pgqeHReA6hp16QO4rsgdlgZhsorjuL26PxSOVZOJVHDe6EF
SDK0Xd3CsU8LWKsO33ygnD7L9QZnOuWhUNMuCPT7z0l5cCPA3YVt1Ijc/Zsf0TZPtvOD4eTrzaDZ
Uw7e33H/Ucm7MlZFlsq3SArMrQIgZvOaCmoOdqfBbDGsR4qcGur4uX743TsFXVPhMpQVnMz5Ba2z
ukrwxDARBIhNhMeW4/H3YtJCs+5z/pocQqXu3pGiksRf/Dddtr1UXdHQrQ3/6IHvc67Qu6iRqxwF
BxAruMiJuC4zni7HXP9eRDSXfpT91HllSiHtgK6iCkspUBvG8Vu66A8o/pcZDdLC60TQc1fjnHn9
K1L4Sj53MrRC1PgkovqH/66wxPI/ZttJkQ7MbFqDN03fjUzh4LUeIO6R1sM0PXljkGT68qrYWkje
tv82Ldkb48OQ8MO7nKrVQBDPinJz/hOfKvkyBCvfg4b298ApIsgP07BVgp7OyruR3rNMY5ErdI2c
/yyPIqTASPgmgzOHoqUah3anyRDuguaoETwnRL0lRZw2Mn9C25kw9yB8NIFsuei4FUgX5mafzcoz
PspZNy0LXCjneiKvpsNEzLfAIkbZjhrVtHKnacOAz2Bdix82AUocdycamOZYv4LxqV7ANIRfXqYK
w7Rif9AixEQHIW7UktxVnUyrcewKrRMpoWSJPlpctN1E7wAvZxZMkXcm1R+rrEYuImB3l2U5o9g+
NlbvnM/S7K+yhxMAbE29cQvLVFi/2Xscrh4TyXQivUDjx/CZ3rjGQuI6I/bKkjKGyojxB0ZZNGMK
xGVOx61/pqz8PlkUlzawFW+13MsHBNXYsIhgEK5MPydgBHT64b4ZyfCTK0YHD9RYJaH4WlCsswW+
RzKcda74D8wxHqNj1A4e5Rc+IT1LTmW4upZJSgaJGAezc14H2hODJUYoJPscQ6YrzcL740xxDLVj
iRhCxHZAGk+2KPUS/MS0azVITyFbLTGi/Y+NnFooN7J02sXTp9zWetOsW7ADqrsxN0IrjaF51eq3
k8h6IQo62WdbATS5trJPnjl0q0Qk6yNF0abUqUy4cTsCWfEKu1z4srZRKEBgjw/7psujHybOlYGt
Twu+hZ3+/J2eurB2mzFqi4zWUN2125jbSLof0DyEnjPJseV1DG1zEL8VtxUH7Q5B4PNTKYZn1+hk
/7yA9xYgOdJBa43oAfsjrctYnLJgSOXuN6AKhe90XF7zcp9Lk3LpYd75bqg5Xr534DA8vD0OE9aA
v3W8mIbs2lpDeGLDytc2R+lN094E+zvDsQZTytbws+UDoRNNtxVlT/F2fNt1f87/olODZCq2kQg/
jlb8oq/6vrxVAILMkf7N+vPJUTZM407026/4/MZ+W3ysIOwIy9nRInE03JLbIMSTTGXtJljUNzBf
7W/kjk5Y4Un0k3eLapwdn5/Tkj6OSn6qTMq1obMnAyOIG+QpCziZUGwQv8xzMUxoO0afgJ8ZK2iV
GoOM9haLAMXJW47gWkKu1RAWQwJuivILkruFt0hQsdXXNV0GuYUwWehjsa4AWe0KEKP01kcmMQkb
YDAZdzZeLVywmr8JM1tY1Gw0Kd5mwc8B8GLQAm2h4O044DbAvbetA+q0wLtiVDB5hKH2Z4PfqNr/
phZlx4vKIVC0JA/sXChKK6vvut4Mp3Kf1pF35WxaS9ZH6+E/0uFlMQeSL9hrKv6P/xxyLMuVM1kU
E+ReqmGRAp4clHI+TlUfrp6FJ5X0+NPWXrFkAjdNnKvhSqSmxeGlfrd4z58rX4J567utVwFFBXxt
xbazn3VIh7TSmQwKgtQFHZdd/lvN4uQ7EMxsGy/VpP0CPTZitnAVwxTNNq4FDCUkEjbr/5OIrFI8
5/O3rnCTYVCrjX1ggmam6VVlQfSUE85Er7TtLfocEXAAJErMGu4IgfGd0Gt8UWYy9QuaHC3yEj9M
XSml8iLmpizYvOHdIHmMvI5Hb2yuFN7MfdT8kK/aNQ0doMFBpAGEnidD2r2DzoMbz97+BDioCh8E
ccm1Vcq8apyKEGLkblhTvOQg7EcsrJEfJXRAWi1AoUY8n20I+ysKB33+XmtUvyNFnhq0TxcXByyH
WF9DvN55MhSGLP9XtE/pJfiMLa0byRKm9y/rjpPggtWe7r28UPs6MVHgz/2YwObe2TluB+j3kpNJ
xmu7Jeb0tSGWcR6E6x90B5PBQw0S1OrBAUlLlthmCKzrK3TcwWtB8O23oGAHFFCXVJcHBIwOK01S
dK4t68IuGxdDqtDdzC9wp9uZQmPJbNLIt4n3XtUJrOr36I+eegyYMG9L71Dcw1+PKqkvEPCoCX42
Cn5By6hKUnyDBgi0ZnCH3LcGUyxcyiJ9OIzkqSNC04BcMMo9G+ElqxCS4Q2rv6493Rru/PzPbWZs
zugk4JhBlO5PnwaoI79cSM5EgSkmPKFgkea3xCjvLnjW7+3kSiiqTqNFC3QFYuNZJ5ChregyaoOa
K3S2pO1GjCqDnZPMM3ljGeYX+71GoJ6gKf74oGvTkBB3rsCjksPkefPPNSMfvRxFa0rrvVvMxmCt
PO1Xrz3tCVfVUAFE7ZL9fVY8vespQR4fSIeWdwJ+hc0WIU45DLK/c+BMZNJGVv5KdyQgSZtlAv+T
P9buNJdM9n0DgZ7v5rntEgyy/RMx5lTuP78C1Lkb37JJZX8wfl5TXicz5QttVi7vv17+4918VgCf
Ym/5a/NKbj4tq2OmF6iFjWttBcUDJ2F1irR5Me5Xs8DsxDfiEhmOFFf7TOlJR9otBaenol5Ps+m5
ex7ftVi5XClj6S3KYBYAXjpmlLjynb5pQ/Y+v72qQKSdHKO+cXffY5iNmOtDu2QLLkUREJiME0nG
N8oPkg/eAKCvdya6CrIyM+J/CtGxzwEEAvcqNe88cT64V1JXlx5UIfpidaOT26gy1gJxW/4zmVHS
JDmW7+OdcaMQHswltIrfU1EdmgsupyvX38fI3kEPowAPyoaDIyIseG9oOg+7IB7fvKAnKu3gJtBx
V7eYYxCBgs0Qh8CchyouSLfg0x/qmcLhu6IxKGa5wm9d9T9MVAbY1LhgkFyJtiCSjjxUkhcRoLsh
+uLovEwkgNozJ1fL6PbYmvRvTzN8ZLSQt0iLKleuck/0dgpwM4Kq1lSbjDPtZluQNGnKm0EXYSEs
pBFHuvAopEmOaIXkYKIrwrb6TDDVRKdvu97xs1aRTKC6PBX/V0yE1sTe5IZujvLEFDOd0Hcneg1z
lnCIJP/C5lB6e6ckLhDe/f5lujAZcfsVGtmpRr3FQCjGyqFhtYKRiGQ8Y9p40mo/LmpTC82sfzxe
bHE8FJdx14ximtBtga76uy8ru4to3KBPaj41o2mZ3iPNGtLz3D+KcjuyLrpSCHtkUxkyqVJkvANO
kZaEG/y+vcSt/op0YZUMZub7twtjZQ1beZTCghGbI3Lz6Nx1mz/G8KiAC79/AbZF24rWd9RoxpZM
ZjTcJUVj7ZR0+1uhLLKyHiZGsOFNP0pb2oIbnso42PrvUHo1r3L4UKPqVF8wmk+V25ZNJ54nVrRp
JduXf9UG3Ks8n6+xeRrI+7uj62PVwwalfDePJtADZa3Z+T9a0txfNL4XfgwnjQBbh8nb5zepSpol
4iYItiTMC8wUEDkmLyY6931m5UJGdC8DESkv78kFyEHCnflkPjoNhWIDCU/B0bBN2OgiYHYCMqgu
3s38C39liDWyMe0rvMV7x4zf0nfwFYgftlV1NgjXJVxCeJ5cALcUZsG2bMaazNf4MtZU4Rx7zD0z
g5dy8IiT7Nyt/7tfBQ1mFEM6wsl+iV2A0/vuAZIZjZhyTQR48fOlt6lvMgsckVCCcURN/4pNrNQx
fKtYHLcYCwjuD5HYmXfbAuHuzQOUtAbCY3sI6svYlyk8eSZB5YmWlW8iKdpXMVIn0qBZcMShiBSU
f47E/Z+DN7NWD7GO1CdAMI0NjxOxDTarmNmJ2KC7vSBHLY99jhDMuMi0BvYxthNc3Iq9jBBLQukx
GhyrjCmiN6bQXH7wc9ZzBbWTZ+rn/8HaZpOFsB7DsmXc4CuGWJrDMyeIPDG0ay95NcWWg4PdIjaY
SYLuk5d5N0phbS4XXI/RU0zObG2YB6wuLLFZqf4Btz6sEjeWP3kZgFEC3gi6PtGc9ubSXafROqDM
NXi486IFDjlR4Pa3zXPsMOmhc8Q5925LHPDoVM/IbZZcAozEU2Iyd44VJiwveBjp2i5FyFCOg5qi
+IKWuB4Rk3BAHILbaR3j2Oe2QB8dvQLPmJt5AJuTptK3QxBuBalCpPL57tB75kT0X07qM1IIVX4p
X9iREglVJw8Oi0T3ccZYbzVNlLufM4HDhSWpwtULr1tYaEnzkTQOD4HQ3u2FUzggH8CJfOQfuC2X
uvp5IShY8yAajMXu4bShUp9rwsfCnD81+/PebYuWwswyy+i15Cag4xyMx8mr7QGFjekFA0zqEZFY
58AXajfe4tpCRw09tM3lhm46Mu+uSpMlX0ifoRDUnAYTr0BY3a+ooqsvno4H5aKQ1XXRGiSVmq9R
GIpwOgsNcyatg2MUruIt6lq2EHx6Mk8pIx58OLf685nNCOqH4+Woi09M3lDZkFcgBgrFfCyZOiJw
IK1K+NIXONmxzjiI3+yupUBUkyGN1czjxHNDsP7U3ymVt8gVmdYD0Jxub2AmuvsCw8ZkTOE22wwg
JMTeKlZzWxF3EVLmIxToZ1aKtyqYydbIpUmxqnKVAeG0O28IM/Uaw6LyD/TtTrBfhMHi5QzhRxa6
YGyy+B0U6s5O4Opqd448znhcInNeT3sguE/Z4Y4fu4320Mv5w+/yNQlp9S4UpnSuELK1iSZ54evL
UJKRhEEHB1+12wolkoNJLOk6M4zzpmga3Xir7qe+thc3AynpE735G8FffvRasO/x1E8v4bYv1VLb
/rKGMVDQwUCnfNaUQXaOIH5QVxrVozUXaWD8iBHiq0XywkskrUlBrxzktUamcOwRn3mvyXDfYfE2
gS82g076QlvULvEbP4G6FvvJS5sSKLjSmKM2TdzcbNQfiNX12srf1wEoW7Uu6GGPXSy9evBtBbQI
l0XR1ubTsYwy5Mm4KEPZbshnv96yAH4MjoW4ie1HaQ+8n9LI3PTDex+4oWU+wq6SSnF5+5kbv+Z+
0L0UkADUZ9oo7O1J/WfT6pZ6rqjkq/ISofbEn4sz797oiJb8Z4IRulRGIUjgcAtWvRM9176If6Z/
2HAHxn/rCQYekOEVLxP15YVx0elR5V7PZOcPlsBM465cS2VhPVMKLbVippXaKvjRUpPqGMbJOO75
W58RckQPg9HpO5G4+p5oMnxuXX1BpSDUvFYf0MsVcW45PwPyXKRZUJpzGln9DUH+owIQc4m4/Sig
EPMduJXxXzNIHfqbjXRmnck2/BVaGo9QuJ7vx1IUlWXsa/c8aA9SvgBGFw7FCdOkvv/NSRGmPhUH
gvLncA7znf4JLGPVU32/WUov/NcN9kf5ZaYUH8OFffHxPDebDxJ49P1EgZOaycM043ZXki9dJLm9
hw2g3xiTbioLvCW4VhSBntgiJw9STHxcVAjJWImv41XUMDtSRTBDYUquwPkfFwwm2WOimWQtE/vk
LIpJHtkloPME4IpvxwvQpSiCvE9zvIx1D7Q+Wi/IXW06sFEZTxtGbc3pGon50drX0XQQo2PflC6r
/2D9JortgcyR7+jD/X4Nt3Xg37uKe/8g293LMxaD2EaIuUq3kRUdDqaPnCnrsB0OQ3OTzhH5Dfwh
mTtJRNvcut5chtKVqVCL75g7G2zf4lgKCAwT9YDcxQn4rb6VCizKZCrqvgKrfxqBbJW2DX/Q0w2C
BYaOWyzbWA60i8gvQAN/XKTFi/Ysj48Js1RluFjPEDDsP0kvo8g+b1UUq/WovDbQQezHOfAZreiq
Lte4FCjdMn3k7cCY6eDS38kNEj/kdduRKTv+3JnyoUemEGDh28uyEZeMHHugqWE5sGNajcklXq5x
gjz7GrgYx6wUxgGMiC1Wj38Ht5F+agMboC3x7jhdjC4Dvx5qvUXCSZxAdEvH7chBrGSjlFq2jupX
hqILseLTJ8VRZoqogI2plxx0HT4BAYR4pBIYW8e19KO4k5792TK9yywuVx93Hh4wfCd8CSnzc7nM
ETDtluAp9+O3RvxZrMHp4XAGUQg5yqXedT1JinBEpVtwx9/YZQzIcDgUeZsmpGfYh+qbEZ3KXcVe
B7T9O10oq7ukQkhFaBDMiA2U3xjXM3vV3rI5YQh2dTzJf/nngr0byypxhSSe6Acw+OcJ9gPTn6CV
getTXloLFy8IkWcChEAssl9o7PSFIeATr9ACN35VAmFu0DiBqVtAF3GO9nuKAS/T83rDAOoklkYJ
3umtD/O06/N5iHKAnqQ2MVvrRYgmGZIfPJMWze+BS9yROs5zrnsYGBhlDvxSJv9MRmhb93Ys/3wK
VY7H6RJlnfNDc37AlvpFbqgNwOlO430oE1lGEvk4sg4nFPu+TGvxgyO1YB8KCwC9lw0nNuEll9LQ
famR2xW4TuuYXqiye+59ClHaZKCTPUZYoyGUzXmelAEmmRVUaEkweH5YdEgIjA5uuJGT47tt1oCe
82dwZUkkMW6FY+v1G+nvGz1pIvCn0Onml6GJZjBL6jmlGzTMW8nPttEQpFkVqFG8QHpZCSzT/fjq
fQSFl/6rtH1JKEkPyid+t6Y9uPnuseiX4JiqJVOxSoUtKcwrl993l/k3Ce/bZ7I+u/3RbntPwjwh
uWVdKox//5xFIzwmKO5oKLJ6OfMaP0j/n5CK86qJfm5pUdoAWZPBF2ePs6q/MlBHU7HED4knhz6i
foeiz/q2Vaz+QNwBNW3JR/PSzfVly8TRkq02s7XRoiPdDdXYRbeiC5haRaGqj/ho9yOQtt6WGE4V
qbyu300JnVj7p++tLGwDWONsQfHXK5EXtiOc7+f8/vtej0dSzRu6sidq242EU5Cim/ivm7pI/IT+
J0ZBDdV8YsMLxmectCeadyvD+EVzaL7Y7mqtA7ncEY8bnkGd4I9AwNZtrV0VklyeoucHycdWdn48
NK2+9xI6zttqkuXP+T7EsZIP1/RBiOBNzQFaljjbc4Fnsi1wK4pnfbwhXzaJ41BnW80RKCRpw+8V
c8oybxrhFwwqLyBh2B0RgyL76vet7r/f6AKYms0MwZe4eN5fToxS5Isz0oKzGYF0B1/c5BYmoslU
I8MkA8UUeHhGIE6mqiu2iKchjYuCoUTTTfatjOGyaWksiO3IWKglfwoVHfLH7deUpdNYYYINaqm5
6GvekwqQ6oDHi6wVkZe88R5mL8XY0mlVtfXa+QQe8y2386Z0Visso3nXdC63yFvuH6aZJnQHA8ci
z+DwZjg85sHUe+uddacEatcBL896BfKK+qb4ITeSyO6zwOJ533VOL5N9XAIBmbdJtmKh/mMMw++H
ndyMmEuIvoYonzThxOGdlA/E7w/EJDgGnc7k2H4lZMtkewy04zQMMmfmXEL7tjPVi0zcfNtftnhw
z/MY6Q+XGBbxtP/nOXtHRe1Am//XKUWHl8es8xCdKva4VzFrZbudN3u71YwaPxWS0SaFpB3nlceO
tX9T7VuYv1/+CYjnH8vNk0te+diirFul1cbu7/M6S6IW1PXDEQR8Z9ed9h1Ij8I8hXTmm2fxRzMH
EUPLzkGBWL4eI32ehxuQ52sb11z9OZA+gk5K0kJwImidnNwMZdBTnxLHIVR0YhBdeiGRp8Tu8SeO
T8I855TDy7NJgkO6IvqCEwoqkqxdsy9C8o6HZ4CmMx9Jl/rup4AX51/m/2kkMEbLIdLaP1jTcQu/
SuRNsfX9v7rcVtremzgPmRk8G/wqeBysnwB5BjpHWmM61NTA/IcLZP6fFNr7t2JMwOKv8aiD1niC
mSFPpFvj1WpNrHGlfkSHYNw+xJU8e5dMr8V388cL60OsIxj8Io406+OOACljyI6tU0rnaE2CykVO
q7TmwCsEuLkbEAVI3GGVy5Ba27KkwSftWV46qyAzKrp+r5h8XkEdoocmChkSuq5u9XCbY9dto0p0
qLQqm10lo3kz4jM87yz4h1XfU6wwAyAp08D8wNb18yBpGbRxCCGOuKb5N+8cdPrCdku5esqI3MZq
XwCsbiPjdAGbtDWr9Hx9PBYoUDMC5JTqUsZWHSDyC3FzLMVHEtpmdPX7p5vtwyJ0CVvK4nJelNe1
8ddUZ5Xhg6pI+Fey6tO3XuZtauUfELjBAe8C/wXOQm7L7x90x+A6l+jci4nnVEH/rJQrBHmbELGR
hGhsDsH7eeblZfnUYmCqN4nM+3YH/sqJ5ohh9HiZNX+ODhF3SZPZTfBKKTd9PDMV3kOJxNT9vj0X
6njEn6n1C9/ybW9Vj5twqBafPvqnyKBXSknpiaX1rUBpA3YbDTLjgBjLorQU8XA941JimKpPay3u
XF+IlVuMhvlhVJ1UvH7WZ2poiGs0RgZb7Y4jDk2WFCG5/XobmYfQ+ycnrnh9YCjA1G6HH85q5Mmk
XBJtabeyjj4k8f17ksxXQus3uY/4BlNewGimQWdmHA4DIZ3oJWU3YEhTdfR8tGWRnh1ohzjxUmvH
5leoiw6MswtRE+5avyDksbcWK7dfmPZvRXfhk4XKv4j540A9h8iXc5KAvWOqwpe4Fcmd+hwu4QNE
JGo494KzMyD8UtLdhLO5aavm8i9fUuaGE9OkWZ1R9hI1ZhhedHxy9szXDbGhRgRgSXPCWQ8++vaL
7kD/d2U78iC133e+q3SfcqC8eDIdCklsCEJ6klxdgQP/XtxLupo8hOzmry/OZMFdDivzpWDfr6uu
ut4GaBkU57U9Zcb+Rp0WmuleiSdbKvidOAT+8UFgsJmu95lXA5ONr0dBhXAC0WnsKXxKUWWbDXAh
JCEmqgbk7q/fDRSB0HlWBmw7rR9B+BJ74Swj+eoejoJeqCjCW3J8xJnSo6lPzas2eBM1R6ZMtWAL
BWVjyWKvT69lyaUtQjgGSI+CCMRZV+Tj90X9OYoSnnOOWyGsvgv+51dXy+zhlxWkwC+tb5ffPt00
M29f48G17mj37CeiCVBAfcLtu4Gz4ydBEJQlbYfzuv6xJZCEdJHxVec/7QyUJEi5xdlXdmX7PAn6
gnWeFjxys5UDlxdCLBl+Tw0YMnoFb03nORhs+UpYeMsZZ6DIrWJ17xTuURaeBM9+RBKegSteHjga
JiLT+IJmXjYKxSHaQ23YAlbjPD2BguGvArz7pW48Zl/OuhEFawcYJsldQUkoVzxcG0jz5K0ArUMO
uz0JG7TS/bFNKrcrBxYN7Q6knoYucj10fRU8Fp10ZJA5mZeR7tdSnER6Ho/7Un9ZMgFJxvlnPgUo
s/7+9w+bUrpEpkngJAlgRqHqioHW97rNS2ZfHRWxzYSCAmZz4M0CgVscxFIY3JHDEqR1uJqBdfgg
KLqo/EpmR3la77t6ZMVcboK7OSqQBZ3z0hCJ4oZ04F/0oJxUIZcFK8V9t+TBZWLzfJT+6uBrxc+D
Gpn/77qZSz+ct7I9HcAohqFBcwElYZnaAp0kRa+PdxyRk827BntboBi8tYHPD4bCVRpU3o2VSj/n
IsObeOPYfCUS767lCwooGBMuMKtvQpyQdPD/4gIFqGoZndHNIe1gqAyWqlMiR98TZu7IdY4jRA7Y
2mYBsQEuL7SV0u31D4c/Ck4i0SXFJQxw4lB3OGWcmyDxpnqAkvHtszteCXYZvMsI82uRKskLulP9
Zx7Gu/CqEApx3dyZxYBmdd4zo7XOejQEbb53Q9c+2LByaZr/ZLPJjOCO52dcX4KBYQw9hApZ9ao7
RubIpna7aGpZBhg1neBBE80WvYKW/O1KkfzjvW6UX5Bt4OB0+DUoCrFFRgTXol3ImcZwKhtQfjIF
BpVZQo7C8qpd5zJWTbhKM4w9qkVj1ALQTtOU6GrciUBz3k0/U6EPYq/Xp8KLXQyDHb3JsOISYxeW
dGLreNsvxIpXWwLrA6wKE9d4IILf2iig2peSn6/0QIPgXO+9PG7e5GSqInAStfwi1AE0o4mbfERd
avZ/YQ6wGWygZfguXxmObVlyVOGjnzVr7xTAxC1U3QwMaLT2SXyqhg+o0+FQwrsrFCBSAC3fyxDo
k+/ik9d3kCmfpucL/WlkpZw3P6+1BJ+kIeL1Yf80U1GHMWVF+lFmj4aFuJIF7puWmNzt/lh5dmgL
6mTYvBS3DfLGmxvt8Z2/g70E+W4KcWBA+0ngdQPFGemPpE8DeU2vEDazcIy4kmioDy6iTV/ttnRa
XS4fm6kRrdKf0GZ892uX45tWcMCx4ZVYEMaII5u2vu6Q8Rcwwlb6kHrG1+8Wq4OamtJSuggagjm3
JzdYDSruKnIzRACuqGfBQH8g+HPvtdTI7QHKSUFBS2vnClzCrk16jSutwSKr/xAliIjzebeqIxb2
8EQQP9SaK1UQNdsK6eeDmWaF9s7nv6FUtZlikQPUXrCmtZpidwZM3le1VkzL8tO8mP/VATMijcFL
1aDGoQRIBaKeCyPTorvIXig+ulviQdNw8Gvi1wenNJSUpTsyrVWWo941nvliiHieXly5Bsp1jefS
qlF1DgzPqbVRMMDS5MVjfg9tCT9uwNp4hrCHWEBDDJChAzvpQ64NEQVyHrEen4npeqOMwJlYP1Mq
/lYtLfD4rlr7ulz7djp0Zn7gwnQbACbNMKskxrIQ080/Z1AiMQ2mW5x8EjU/E+prs/CdTWrKKVgN
OmtaM0BAVoc1rEFaiZAaX0LatudMph1q03/ooMW+RPaWzEE5WSr3Q4y30cXFg8fY5gvuvHJd7ruK
1Ul1uYAVj1Lx9siQGjHqgjKpZ8Ef7c61R7TC/G2OgTV2gU8y5I/tC0/EBZaEvbY9Q9GdGq07Ri8C
wig9smlBBrZyBdkS/BwbOK9Kw/pI1rL+fIBEVhjR95CKS+qvmW4FpqVurobIcawbcZp6TKnWFwVt
oUGJp0mUuaDx4uddwt6DHYbQCV103Hq5/DgTeDT6N3MXpz6OmE0ErAD5S0gokOdP2+tQa2GYg+7K
wmLfm4Udnq1L+WH7vm4/eZYRTEb9hrgpbpJRr6fEORLWjeNFf9o+X9yRitd7NTRVwr9dA2jTK9IB
0i8ZEsrFt1P2p8b4uSnWW3GDLyyi3NwRVBP4pJg0nTZGhi2vjfGFdA6nK0Qx0a95dfQXVZG0Ou6C
TAK3010QA88CGQjHoxNRikEdP5r9XMv4M7ZladLnoDLp3PFQst9NZ+EwzddX+lB5yzu+zomRcUuo
1rjmUi1j1VXTRW6xx5MFHIsV7+VagEIkz7LhjsotFkgjKWz5tsmUSbtTbpPTtEsUqMW1D4/Ydued
TakxvDKzaH3XnE33CsK0VCltQ+JhAC9McHrlqI1yyDfNXb9YPvc+HZ7qSn78Epx587Dx2qh6g3OI
0q8uESTLlaKhvO32EwoLXx/QGIV907eGHbQ8gjQyYq0ddidB7JOStnaXi6hv+6gxMfZcaGvGQK6Z
ERB4HcbuLhFlQ+Tbp1VbUAQYiQb629wk68NRIOKo7R6Y0Sj29s+T3o6HwuJ31hY4BW6N6IzfJ++K
HPRKLedXSqUESES7mlcY1/pIE9F6E6lsAWezsSuskZs6sbbUFSHknEx8nQSJ6xQLSbocCwv+0Ph8
Rym1Au3V6J+rbwgxGqZgx9/hd5vbaHJC6OATtA4u1/9NJ3KjFlHvDUiqdp+dInLh2mYZMtksRqr+
5pQ357229X621h/nzQWKTdffGNXk5bCKzpMXBMgngw2HWLXLM2NM6y53gngUGPYUt2gIakNMqzvP
bInkloZ6Utf6pkGW384razPUI0HREa3m2a5RRqgR67w1D3PEpGjlx7acRenebxC3Bv0AzQIWXp4U
dgbGOnLr52ZosBjWxgfkeYY6kHsCBRojJTICK6xK6yltdH/Bsy2sdVrcUCtrISK7E7lDfBC1vvdZ
s62MzxRHUqNfq7VOxBuMGnhXAKyq97bm4mfAV4zorMhNMDALwhht0b/m/1PJi5e8dVs4q+81i5fu
xPpvShfFrf/ds17LQmWlFHX3oMM4dy/qQtOyCA73P3Ip4Crd1WTE0+piptn4iXMIxGiE/SVa/pZE
GHqZPatw0kZpfA8l1JsapraMYBPjJnfajthlijxxj0gd3aStaq4Q3Z1xaG4dWUJYdv7GFRDxdquJ
qi9RlEtIolHcD38PjtVz7mn7JZNi/AHMcJ5xGIvi2V3YIKfUToL3SItgYsw8uhgnSsJoMgroS/Jm
QC9QAb+KGJh0r9LilIYR+OXNVeEoRIz2GpKE+5mucUpMwoOfHajZ8PaoJSGiTy/82jsYfqFpcFa/
ly29aN9ph/yC3K2tyH4bMgBh+BBoAHw594loW/RWdfitc27Rexnx0UhFSmEhBBgBE//fk6zwg4yB
4yae0trLBZWjCmm+PxNnAaJRlHOP55P9yFOFMa7HnbqIbFfpVDOXi3WpR9N8heyw1L5AZLfutnkI
8pQmfd6v6N1vUfKXWdOVOEsqiuHXUHV20NqusBmrB05sy/3J0giqJwieJcPbLl36I3EuVNO6AssO
aXmJzsBuwDW/ZDlzw1jLVvCV1NERtNL4s4TYyv++DGQTy7WNF6G9HidYHLFl58Q7AqgSK6u9xHTN
ZBL5uSjJcsxcSojf6Dz3QrK5QwpxFL9LgrGTIH6VBOYqONSqNxVgSoyc1hdU3jSBBpRBCfHwExBU
cXp+0b4SekqVThw7an3ZRXdtN1jpj1FedzJL42RpjnDPqkV7EzKzMUQZ6T6HzO5uXLAgOJlpC8OH
BUgKlIv0InpW0MDgSXJyC6oNlyt8dyL7PVr0oNUT6DyfDu+hv3uHu5kilnPNnErNV/2184vmolTA
tyXXcs0VxXUduUYeXd1e9IK5PwVbOa858WAEKBx3Cn3DtDWxGCEeETGVSG1c+ogJiTSBBB0d39LA
eTHPf7nv+k6s1CSoICMfaMA4NrEgqPmoXrU+I1t1wcx4ihYGTLhvo0TeFj54c0pD5CjkTeM15EmJ
23OzttAQ4qe4whc0q7lTAe6GIBq4cjQZiP8HylPvWhSHMGfBN6cBEYlTI+zadkSxLPORRmSRtBHi
cDIznGZhv6oEGh8HYepa1d4S46C80OQVB3uWFhHkgeAjdkBLdutXBLIizCv1h2yxEwQ8ns+2WlPo
+qvb8A2/NefDfK6E6AB/2ySiiRAec5fhreDkp9UyDMNU8PHCbXN463vW/zyTWlUYDFJrbcv1gIeZ
pmCMsIiyizZa0ixHDXgALdXCAAKP0ed8h2ukAZ27kHABCeVFBD0RdRMyI6L/ITlhjn87wE0Y22zH
UALmhLvHtPPLlwdmVtPuG9xGe+VtfkVlR69Os3tCdNyszvoK+yI1C8ud/ECdqCHtZbsDZfa7Rn7g
xyME3Asd+sKaquh96AOMK/gEboXZcZ54U0SAFre//P1b0isvkSUbvWEuLeSgQedftxZOxxqsdG5j
mnkwST0pxTaPVwv76pRs1hCRa9kTtDiTTk1uOkDFxEhYmW4iRUGF1JG79NeBRQ8gw9xvxO7HNHa8
X2ohdxiB9Q1Jhy2MUeTqgzvrPrO/5/CeQ2En5b3h6BaE4EH6HM+3YoCcvXyY8cKDgmRnv9TAt32D
7DKGb/KaH+PxlTUypkvBow0rsxC+So/Y/n+Q+OVREhTKlo2RjDtA0oQUhTYHFc0Bi3TUdL61XdQO
fruj4NTl/B8XsCC9UywCTz4QEqzXDfj4RnUSLvHXq073I4Ju1otOT4qfCZDdDYScmKD+NDlYW7gb
j0Stfr7fT0YKvCBDJnz7OvRnxivkq7TAizdYVyy5UHsE3PP+NU2i5pTKsrBUOFmgkgfk/w0xcZOJ
5PxTqFzlKE3BfJ2WreF7OZWDw0pI/i4Mc+lnOnmTVPGRL/Tqyx2QnwOsTi3xsMCjogaLGJh2jseB
SnSO2cpoltA2BmYXM5cbZXlN4t4h2HiWDc/Fu/zTH3mo3uABOrSk6bWumiTnPnk6oYuDjZ8xDeR1
kWy1xZmEXqwqdVUZ3XnCee2b6jJlwgjUJrL0IW9m0A09nnQiu1ggF/n9yZ2FoSr4HnpJwgkKUNSz
JwE5wszXmwN5TRsCZpQpA8zyZg3eEWMyeAwmZAlQHfQgMs5KScMjUsJxpRP3IlMXL9kPCT1aBNjR
B5sGLZh2XvKwThMYagwRIOSGEniFqjldSrpbxu+TR8T0Jgp13M76E2Z4y8BO/Kuj1oNWPNEA3/cO
139Ih5N24ujh/dhgBIJGEIhZLncEYKj7dBqwIc8zR6+dM2YJVTuIj5p68hOJly8aHbGz/3FLBFeS
MJU76Y1UJYPtjjKIFK8q26crybyyS+nRlUgSRS4rvhM7fQddC7lM0CGVLX1ArUSSPT0VaKmuroWR
6mHRoTCS2W7hgNNwD4DAp15CMArVF6CYwroIxBIL1bCIDoQ9SqSDCmGd50W7HUqnqC8E9oJIPZXu
dkiSP1+oRC1rnjgVJyGORCVNiIoGGHNhsrGmZgA0Y+Ob5wpnJbbp6uWytLLEOOAFP8jN10Msl8An
mOVSYxK2rm36G0AeBcZEa7nHPZ06E7sxDCcGJ57ubNa0j4HMSBn2Zk+5SWez+AldM3oEDxzbUwvY
qS4NvYk7VZU1QuxJUgf25kJZtReBF4H09wqeng6R73hAscIRc2WhwHPoOf00BQcKWnztHPjxPPIA
NEXM2OvVqX5iBLCyISgZdS+cW6FYekHPzijBdMWqHYGVeQbSdziFl4M3I9DBg3l2kt2Z2TmkJwRE
yT0DdCmNLBcHS5AO4IZk/CrqHIeb2LXx6ZnThq9ybEBEVL0PnPlqupdou8r4eNUN4nGDD2tDHPgw
3cqYsVCyTCLDb9dseE/f4yDjJy0IQ7No61nR8SZR0NM8JEb7ioEAddjNP0zO7aPUn8UsKTDUk8JR
z8FxX5enOBNLvEvasEakI49JJTMlBSca/8cff/U7/RuXx8WBd9PdZxatB4Q2ssnG+wDSbYdZyS7X
VNjaY+EGOLHLNrRJdkizU9xR3nmFGhX9VjmB5WjfwN0lXmN3WqseeMs1aLokCErNGEhNi2XPiaQE
ayHGsvbsF8qYjxE/B0Z/a+CnDOF6MUk52P+GDMLXOHHAAz2oRt9DYZZWdtSTv3fq/xM+uuUgs3Cv
BgYAViwVkT/kp8q9lOzHEI192Mu/NkqAA8CYfuAAbLU1ympfa9k2+juM8LXvorXkS2tF0Bj2Dizf
2vgidnzAMm+99B13rxa/q3qBNeZHo5w5XndtHgL5R3PVimq2jXogIeHdGE92ILYP7ljPLFEkUC2n
btuYHVhsfwU0kraekQ2FsZ+6YaOayIsTNsd4kNf+pbsIeDRiqslB2JiPMoExSqVSmyUQU7gNLpNj
jakE0IG5UHwYIxZT4JQY+MkhuUr4ejHhqiLiU0vwUd8uOVZB5aMTeft9P8yFTFmLuwaTSKUqC9qg
F1F81jRKwn/VTpZwI0+hHoNpLeIiP8n8dZHr84aV1MfqLlfjHEOf8wqtCqSPDVQfuEjTxHtZ7Iwv
9kWaKYDNg3wjTSQOCQBZKP8YpIJ1jqIlURgaryIll9KC1n0VGeUJCTBOTwoLpF7apkcq5/VCTZwg
mDzH4orwdSzBlJRPaBf9AeaF/ZVBWO3agEPVKOjPtKCqniS7K6ZRXLyqdUVLXQJpjwk6VGh6lynL
JK28ELjW7YXZcVP3MG2ON4WMAFEpPK8GJUDE7+kC1rwMJJGJ43GiS4VU45ltSmCNgs1R0pGn8eUd
I4Lg8tQP20akNYCzP+EDfx0IcVKvJoTWPLaCsV54zQSAmnaeUc5Nwierl/Q/Qck4clfGjZrdVLRE
f7nKMu6ippIRmAKA3bQCZ/U0W/Ah+NmquJ+mEokBKXJWC7QAyks8GyxOkU0+69eQ6oCFyvXDgDQm
1bFvP7hJr2BkX4pUCjtncVHNWF3bbySJw+Pgz6LO6OnPjoGu/AOgakD7av0sU2wtfkizqAY+q34D
fx1ip9MnCrKvHf9s9I3U3hiPoDkqTtGPg4GxHAU3grLP4YZXkM5AYjcZAce37/y3BJL81D3q/pUr
3GRHgfsHWpl/HoF393yaJLoGX4mPM+KqBr3GIg/iRB1TLrra+w8mJhmaZ7my6RJAifd7hUGc/lsH
6aYHkCkkO4ZynyMvjIWPVS+NwB5/nY3Hsg/Ft5vCXKttSqGycLlSCX1yf1Et72bnxcqtoNDRnjrs
0jl+1Gn4SpwEuYjWUb5knWPslKquOqfNUZ+ry1LeJV+P3J8rgeCPf8fal1dD2WMvXx79G94aDPAR
6meSic5aQ2GhIEJoiJM4Nb+s8OTlUlxrakTSkY9fMCxpeRIFKo0AWBOHRHBYfc/0f3b4jT9zl21e
kIg5R1dhxoxZlEZaSYQUWlvouYq4IYjb+djU4oNu+v1063e/m7IT2Yeb8zK9kkThldKrsu0Rq6yT
LvGK9xit7+l544t680AHNzBXPGkXg6UTi+RRkDQVQtYqlAY8/RZFDA9r2f/CitzoKpQqLZcDOHnZ
rh1vZQ7iQa1Iepo9uaT+CpldL0/8ngk9fPEKxR1JNzim1f/vC+nfS74jblJF3/Ohsc3W0zRXZYzc
joW70p3cUwxDBeH9piBnoIbM52T443NlN3AOVYPVSXnzr97kfcoCVDVuyXWrVpRb/D+iAoUWxs/m
33L1aL6bs4YGjL3nZ5Xo5sLpxKXnq1Cj8+xGIYKpAMtJSKX+gttkF/38fw4R4lh6DkL3X4SVBEjJ
9m09YQhR4S4Y9FaX6ZDsTaQy6E8LWzwnZVBRWa8jQtK9l9ZokHAD7uonkE021ntENJOm8P/pLyuM
CCNf+K2lKOWQtcnVbxphSCRbEUo6kA1gAj73F2rXtllHumelUdY83IMXDdhaeINoJWdoUAYWefBF
l+mJjvCrL/fTk5zrUo2Dtjs4pxFTtpqiyZ790NsW/mpovGlzBEVXAIlrVxm1j9TQnGca54fgyDae
NoKww881xlZRdgGwVURME6zxkF3RvWjTnZGdZwUkTQAGELa1dg8gb2tgV0/UuzUGdIKpZvi0wM8p
aiN7e+raFmPtEGqJn0gV1hrBxO3seud43ETsPJK4tbJwl+V++8XD4VsCkJCZgm+wWWAbXx9053rR
JQfUvFL5PKPU1HAf9C+46QOeNYpKTBgNO7EivReVSRSVZEBE/0C0OE6LwtYaY+3j9UJOwI/xo937
CCkxKYVZw+kzcK+JVszg9ADyETtkthGeiczUSpadyvECq9YrlHyQpcX+ih6TGdR2UWzRJ1BmKcan
9STMlhfJBwwVLAzm0jSNi7IEIt9Arob/OaFee2rHOVSRJlHfWytxFsULUo+k91B6LIaE77q3rpmp
IUnNx5R94RlJJCjKtskWU6zqiruU4GAlGb263T8hB2PY+qRBL8SldYywJdQ4P8Y62ApBtRz6vc6D
YfhpM6esuAO31rs8EPdGm+BCFUcafwEIgNXNNOD6HQCa7yQkSVNXUcvjsAiF2SQtV1xL4Kns9xF/
qnwukOmC/5EUZBNQU8XmqB/dk8HbFRg3szRC/490FWorl4dCzti9XR6E4wBhyQ2vEiED12lcxGML
tLSRgwDT9ipXiIOsksJ73z1U8Zk0Wsrody/t7nBeiExEA5jLOlFOQhijxv1b0m3E8oupFR+D5QRA
MT/K88aU25qSMUNt9pSYxvO5F3uU1q+l8msZh0rdE7sy/2dObxQ2YlvNgM2Xkx/YJOGtcu01h8Z2
phHCt6mlBzpVZ8QBieWArWTCWGwjzerOKZEcgEnl0JY4e8lHjE8/AePDPKE8JlhV48ZTeVXMnThN
bpe3vW3GYK2g24serEBkVU0lpk9C5NrD36widRVRkl3UG8TysBU3NYdvjsssWmlQYndT35DumpKq
N+27BM1yQh5/dHfeKrSRaKRoE4XskBPP69neLkAJFH1uQdOEMHUyzRuZRWbGJpEavcE+4dvqHUOf
vcY64tQQ1o3y6TbrUmFYzwoI6KVRLdtqN4hRdpbxNPgs0kIR7pD9vvSU6xniHSXP2PblZiRoF3dt
bQ8x/7FQPkkolDvTzUHT4qv8dlPANVo45FhvEcgcJrsDBrdLHEveQuzpIsjh3TnaNf+1KCvYhwLu
nUiX7L2n5CI5YRR45lFFELT6+aEsQQ25079cVwtejiA/yhBW09vSg2aulZKw9SxSG9dWboQ9VOxR
zKXdsciLPfA2KYCQ/wcVX9GB3SMfVTB18NQaiuEwyZVql/ccn6G20KvU8EaPsivPaf1L4uT1Xq7l
YcWyYoQkvYTeQIRj6O/hqwZfPgZrV/TxQDQAy6AEwvMql6A5+OAzW3CtKTmAhKkkgQ0KDVdTANPO
VZfr17Q9oYcYQXC89zOsL/NzjP/9FoBaxcyyzY5/AOw8UlEYUbBZCPg1ISWTHtn4lRjLlKJe26SZ
F3mLAAtXHr7HHfX0UhAtD6pKrT5aWJmgn65UBigITVoCB9b+oyN+mKNvZA0FkOVsu3v1pV7wm/53
PnOP4EpZgM8UU1aHPInUPl1UiGa6v/idLFh+oD6Jh4y4n2JJi4ruTzktXexGAo9Y0dO1w+VHdTjB
zDIjfL/1JukFydOq5Z1py1IPG7Fk2CkTIpTRNrl4RdRdcG/eg4PZi9ghtF1vW63qZkstOy0AiVnn
JTnt4lfz8meb2AILoQOhzHho09M2+Hjk/8WE68q7sKcx11DoUN76oO7Y9qqwW2Yv3gt4O/euwOK4
ZVtB50Gj2ex/MrWZw7QCQHEgg222rjbCZhvMUxcxGPP6EpcQKBucMMpu0FyUhxZqw9TthKSta3sm
vXnhMpySvqMq3VmHOcldYvIVHPCVeWu5qFVh8WF1dAGRH4oFF5IFEn7gf//dnzWiV/37cfqC/jPS
Drf5s7uYHZeVtDG/XNj/D+kiNH5hLAW7a4Dw6qDmfokKf1zx/KbCTuioGMqI8Suv9/uxZ4KwUI2v
t02Mji1J0zyH0hPDFLm07qHdR2f7j5RLOadyMzlaIIk0HkDY8wKG8RAfbyubFyJW7VV2ojjecsKi
BhdKiDBZKnyTtOJbd3KKAafRmTMzM2IIJx0XX6FRULufjfwcbNKXTVZjA4mCc4ppsUGjQW4V+xR2
wM2yeSreHJ5sW/1TUQWiNKtYPvKs2sN2VEas0aI9mTm2VlkFhwiexKLCijsPFYREEaoU9giz4Ecx
EQo3qbfMi4qMYs1SYd3TeAqZLxMjrMk62ombLAEL+CuUnuoRlvokdiYRGw3sWmpkox2k5BWAmKX3
12nsVi7WxPFzGLXJ4ABo9cTbHJeSHv/hXV2O0GVAGG5/nFthI+wWqWKiKuy1Slk1QQ9gc8QNy3Rq
ThIu8KI/2ORu92Qh6eIGXtbVSHqigpGVb3rZJG0tE9upiZYRLidAMGUa0xGVe6Rbc2g5UBpwlFTx
BlNbh4ouxbN23ylcHLLCsICw1APs2PiF64jHbbTAJrY+liecLwc1AG/r9PeFtWHWeTW15b0QMM5D
YNrbQew5lI0D7SXt9jPS3GXTy0q0rYvZrOqzx4q1IPrnuJGZuoJQCWtro1tyxrIobrSZjKy6YTJ1
f2Fb5WBKMIEwnFhCNepc1PDAeUQwtOagfMA4U7PleLWuF+3CO3xmBv7bRMVrJNg8R6ocjbgg6z3v
Bc8LK/jokgCSYCTBWcqu2MIn9q6So37Yrvwke6wd2qKC7nfV7nVor1KMqufFXgWVgKe2eTCICexx
e1gROsBO3vNvO0/XnvrWbq2zKexwsXn/hAqWFbIfdURTXMUYl45CH+0Iea7BarM/ORzSgvmXldHl
2gM48G6B3cUzo9lbr1WuXKOuN10VtXDkNjaLKVyRtmBFYFVEDHEYxR8Td2ksMAYbw3vSre0lPb69
SuirqzIFrXeReT+80AbRsepX/D6tlT68wCvuhcDrmxSKX5EDqbOPEMjcQuJ9xdE7JVkPn0anbI+c
FhOqEsEChBjsnLpDAwPj2xdYu6rYoZampu0Cqh9Ml3FQTR5bPtSdfzdpUczPF1SG75BI8iU2MvyA
cH3d/NdIdbl6ZnByUGubvKXDTXJVq67nC2AX0RL/H5r2RbezmD1Nyi+ibACifYru353TWE2KoGFm
HawBj59puyjuqiCtLXEdLnb35bpAZaAUOTVtgsOz41k91LAPt9ipGh9WFeXB9k9o7UakbLtcx58w
h4bIqtVAzJkE35lQ/YCiwNp7u7TZzAu7SMM64rkhsWq4Kd4AB05qmMI0rZdIDnlulAambHXsXDYc
mev69RVFvvwJfAYyA2EA5F0fWjEXTGmcKlZtsfRYpx0UcKMG0nolgnL8E8Js/ilx3Ark3gANweqi
v72rCltKeSDUGrhLitekjHHizHz2QoPnvhp3VcSwBrkqC7CPzddy+dlwt8MsDbOkgcd3GDDj8pSo
N6IijimyXeeETsEUuUNFfJlXM1f9ye0+3TeHsrIUOnJtGCwvrUrfk7PEkSCuyrBDXbyl7BHtZ6YX
P+Uk1eWVi52U46ZdPO6jrf5eqaF+bFNnimpOnXfxxSKcZ4OGZ/xfbvaPJHjEMse4KUJPh9alkUGh
qte0l16hK1xWjl7ZuIMSI9GQ9rnW4sBrMw1RtFmmMg2YezJefYh14qMlCh6i/0xItQEmO7FKt3zE
0m7ibFx/VXv/e4Ie8Qzc2T3N6vlR8rxXRPOS34CMNpBBzXDJ/ilM2IAJje3obk8Likp6/eZ0U1Sh
plHbt/R8QPXaWAJqVdR/v/J6yj6wFULNv5ibIlagXZFqyX5a9AytIE/mPJxxOx5IymnnjNtCsko8
EEwF3RjZeEoV23DRLsymC2axfKP13ycXd0G5/bd/JMYx/42yUNzmCU1/EY89gsa38DRjhGzGKwhq
5/hzVNqxod6uiBL/z+I4mPCP9tY+P8L0EHvxkPiVy4pmE9jkK8Zprmw6JzL10C8IPBgmM7nk4bSI
JLP7cflNfRcYEMFJ3U/+H8hZEV5q34nE62kzHFvB5G1mm6hfib1eXZlbWRyJJs2YZiI2CB1NXTRB
FGUd78tyKhrtrMgIxPygamorjRIFYYRwdeR6PkZVH/duPGPr9APjXd6w69HAKTwjlGaURg1FwgK5
Vxu5eQaCNLILX7+AOe1XcTRK1FrhaBmUtwUJc37VEn+76M+oaR/knIUhv5p2GlBOI2qM63bQ8T5N
UQr4b4UMoAOid45M2Kz6fepUpbEdodrttfyFPr5dzk/zGDhvOY6bbL/bSAB1P71hbmwhS5akrdJ0
Vn1ClpVQTw+h7a6PgQfSou1R3iVMGutmnlUKOk4SQv6Rf5dLsqD3Yy8WpCoZODPVCSevj2BmgB8R
yntILbOK9D68Hi1x2VMhH+NlOa6u0ApRMvFGYIeMppJIh7I8lW/JdIfbNs1N7bOnC3M3cFG6iN7P
0jCzjsRGSlY4afTlbD4Zgi/9Z87Bs3pLLcihy5iFZZBtokxpEsgkYyY8aOHWt/Vk0PuEI5T+EHmo
caYIIk10SwB0VW0Yvqv6rosw/wz9hgK562DrUtCKlp31bZ8ym6nLth4y+qpP0gu99d0EdyePZkHm
I8mcvnOsNarRJppMS9I+9o9XcnrUjUEhmRopg87tFcWvDInaqTcarGEI0154JYM0FovRre+tHYin
+VXsMesuwRHQ8wMjOqUksJGEfzWHbQR/idLPQlfJ0KhvE3T+LSDvSm+0KkJy+imKmOsiJ5q/pwPb
GJ+EH89cmzVgF8DK6TXHpeWVLO5FDmKh8uSCuubpfGLYT4BKlt0Gyml/N9cmOOicVNJ2lCWZBnCo
fN44/K1J1o2JbGUTTQ6z8tcrj5G6GOUOZhjSoTt+xdNe4rGT1/58hBikwRTWy48hd3eJEPQ5Pype
tDVaZsf4yOX+ww8Gg7FMjsKQ1sEKnwGLE0JJ1TstAM0PkknMhZtAQzGW4r40SNZHsM/Ut1xOTzUy
iPbJ8mvfMKMZKrspsVu1W9tV4KIw09Ev9xhWSWCNjylYlvDpDJPPwSLdI4Rt2AffmFOwEK7V+5M2
c/ZV5CF9q6CFdfM4XdKb6lq2T3FyBtyXDzyYTOjOCiES8ibB8Gmt6ivVICNRkCqjF41AhQbeaaXa
VBgeo735oJNCPqdQxCDgnlnks3ClEdGUckfpSLR8AnCXFWBSBG2+MK/BCFGQaBHcThSB/6KIPJEb
SAY1bUrnXxzZm449hvbq2glDk/c22XNqgvcGtpMmKwyzZ+JIcD5ut80xcw4ue7GEFobF6+0FyBHa
Plkec0GiRenHXDYa2a60XFdwQZlBAFS7xuli4mXwINPZV0O02uIEct3Vpk79JH9DSDHY3Z5ZvqfK
zkk6yCHncUjAoUVS5aqbde6y3HOCUKv7cH+u6CVMVlLFE5ZyFp9cF20oC+UfSaeQ8L1fBnNz6A2D
yGrrfdRvyZFtbBtaQ13eJ/xYflWmHTj6lRo6Sc1i1GDZV7bqDaxCUVsdtiLZWxNUk3RZzcGrbwd1
t5yvjNmLLHwFlHQtb/dOWgQDV5kS0KCxfWw1qidoBqo1W7xmXv6jU37UOJUoJWVJScQ1U0dy0MFP
/6X944vg2v/sRo+y/Fj6NXOS5BH/3dMcuxcdFvCaj1Hzn6lZs0tLO0f4KUja5uCK7v2ZLTN6NeC9
RAk9EimaQDC2bK+/bsN162RMMc+SkqiD6gjz36EEg3kNdLqFoFr3MSweFU3pwAw0aBmpC7WMHgjw
5XMprrNkGrsuZnXuhoaAgmd23tPVvCOCKLCiPp9Vt4FqQzHi7viwgmpCJ3HnbjjshlFlr8LbSEPf
lqhO1Xh/jfNY5C9RiahwlWOoK8XvUgAXDEf0mga4XYcjB89cAOoTbooA/36F4dB0WfZV6JRtg9fV
JadryAmCm1+trjYFjXQhgRYu3H4Wdwe3+PwTIDTJthHbiPoqACHObLgeKcEsCaEi+lO4atUB2vcV
YrngsVF2x+2J7jL60r/JhBjnznZCyCB5BjPJFNL6t3reRa+Scl/bN6J/Okeb5DvAtSDnav1ySFHX
3RljU7BpvNK9s+fr/kfGSUu5+w4vu0OZA97FServE/D3y9acP5f0zds+bQXNOcv9maHD5fQKSBTx
hTg+eNBXeRmWLCmNnXH3d6aMeWZL9SbFIP7O1MgfN4oYyUQTxH770X4V4Yly2SBhNRCJPc/TLXBg
lUAoOlUeULYTAvTogWI2OOFB00v6Pjo0Kwbo2LMgCD9SfpfsHRyVHclTmvC6s+8GumxgY2AA232u
QhVHiInhtofRs1hjy4TC8Hn3UNIEkARfdTdv2fKU0zv1eOWJsAYbh0OwikXpF9OuUlIR1qXRsl3s
14LRfuti2GdmdrpM10Aze+UhIqS7lFnEeSukRV/YZZaJYGaVs1/1aGj3nwLnX+EQE3jHcJaW/c7R
czthbdpG2pj6pdi61XYOO42wEh0BPR+PkJm+YZ+//zmWu9QDWAKEKGE+UrITVHO6MutOJw5FVO89
ZHh+3nDQz1t58Y/KwyKne8VqiwzvgEvz69cy0q4y/7uQhgLCHZNjfpXKRA8JMFwXT0cCt9ozkLqR
+w/09j2K3dFLTRdcOChxL4urQR7JuO2RrPpSN/sXgYh/rE+AUtPJGofJceWo1LCHHsOwQltGow8m
iDkQKbiNAC/6bKyMkW9Kyg75e4IhbWce9Z6AA6dBwCvs9qyp5svxNEQihT51zTBdtorksQTEuRJ2
Liko9XTGreZgULq9b407L0JHvQsXypOg+EEM7MHlwkrQN51FFviXlrpae62Uz+I5xnIWom+SIBSp
3Yl1GrasoSCPaLAN6K0K4w8rcBnwwVZpQpDG9C79GMMqMIzYWys4z2kFSKg9ZBu/ISccy3A+B+WA
ygQj5Ms9i/Fk6XfqJIjBeAvG3g100wMcNwbTKHgoiVq/im2wuHa9TwdUAdt/zZN2+tRyVR4En0OY
iOMfVaizrHyz2Tgjy7ESOAs/jQ1BKS7z1nVN5rzXxQlKlDqLgrjd2cDNhaxewHY2FtmR+KDmK8/I
Jco4JDpErhUUM7iUmsnmrHjUiZVCe5fV/+xCrsfhw5W8djE81YtY8ILDzT9QBJSePLlq+dh/PkFj
lA3xHSgv1YiOUuGkVwF8f1FPMJE10RSLjuC16sWrq3KlaaZL+RX4Zoy9ptZA/BCpdAmhEz+/GvfY
ZNlOKgTwxN/zsImQptzqFR9uBYdr186IXHJKMCMJ9cQfM8aioJ9F0FRc6SzfwHSDNtIMJMvAWIzv
jTjZT6Go8Q3xfA3Q7qdRx38JBfHeOkbHVUtA1TqMGd3AQPZxUfQKdv3i9q5sMsyJpcoiKk8mu1xg
tAL1Zl+2B/IwPYX0M+NwPGkCGrz+UiAfxhZJk4rmkPxHSrMRyGFcGdTMtA80733UliMEuvytq4jS
AVHPzYmNRdEtyXiYx9NUKgXocfbEmwZ7FWJPQZ1H/Nd3X3Qs6td4qp9lW1YleXZw4HZc02tmxLZt
uK+po7l5T2MmKN7kYEuFNp6BJuwPlI4wb+nsM3HOPZEqpZ5Q94dOL2uHFtO86PA/xDf7DqKl1f4E
sMuexkm/eia5bVOmv9ZqFjLb7tu8oX81i4ss6gFtQaBZIT4ry0j3XUXhefohQrnguy00s1jfNgaH
yYR1mYYcu0MzNOTgCnOE2Nk7kmWXR+KVgu5TBf5gp3AVc6iLETx/W+tgqB+tCcmZyxIpGpYffQkx
ERuSj+My/3M8oUyPhUWGcl7x0L3+8/I00LfkMgKUu/jivsOvjuvRkLyvA29+HrvBMlIU5dW7YXLF
wDqcidPvXYGdhE51p5JE1OwigT+ugwYLxy1OI55FLb/9eDYUvgt2S0eRE/O3yUmT4gAH12tsW/qJ
Ru65FCXZJyrD98aAoUVKoHgy7LuzKXXhJ+PI8Q/q8WQ9rfTP/ThsfgNC2IGUCP4MyEN6lj7OpYUg
tTEQ25CbfGnbpYVWdDhpEAxk6GFS9BODmUDaQiuSrhCXeibS+O9BFKwD42OqFZv35nBENdF70iLq
15HkDqOCHqqnJER54fpqNI4r/knp+Geco7SqXL8BPcoT1dDO8QsYkgNYyLFd2UV27XrUbUMdSt1w
B0+ioY2CrZJ1Rm5jtiPmFSWNuzxCzomS8be+vZXH91ZGz5nWzjBeYM6OpTsAXnVjQzobbOmuJhrY
QoA23VUPO/AL0lOo4fVsWYg25zCk3fVdzB+sHhY5fwEczwyULVHDjGuaBaZx38fAQde3RaXLBynQ
Bk8kmT/X2Mk1Z2r4poG7R/m+t/FLbttYmYrX7VOxyUgIH5CuXk6TdCdLRhL+XdkJxPL3YPkNUeRI
S1g1goMScoh/MvEQq9j6K7kkhY58coFlPyie8C3K4e/4dl4by93ijHPccFVY+IBz01h47wuEe87L
XcoTqVvBGAocZWCLSSBtkLOX/62cNwrn/EkUaLm4kbYctCgaj/yTmNsmX0DatcrMFoAeQcr91h/b
hOAWAB7nPtJZYFqHEo1d5M58sI17Nopi0Rsf9lORMVbvcRNi/T8+9pocuP3JZuQq6Udxv0gd7vVW
5JP0//rcIBms9irtGzkbx3z354EE6Lc91fQ7pCao/zoaaC97JZ0WY1duD/M2yT6dOPJ46j+qGxFE
TVFG+X0ZboF+w8f9VBYZRT7Iz4foaZ++mGCcdoWUCeQq4oRI5MdFtF7rT/tZw7LFb4xduwh9bfWI
1mEbZoCS9iQFQsLSAyNlh/bthD4fG4SLlyd15mb0qUG2KPXqLCCI65GfjKvi1oRat2kzAtbDO/Oa
WUKdxXoenxEc3EgS6zVyFgezM314OARvj7HbydP75SNDdW/f7Qx8aV+JevSR0LQHCdPTbQP0xkMP
GJkkMw44naUbRf00JiUKwiCJXyfNSv9CeOjCtWVK4ozSMi+PWgd5H8T9H/73EbsHbsUv1UkqY7cb
wYmngfA4k3tYSp3OSopU4uTqAJL+xo+lLpnfHXwtwKFUAXix1PMCprXhCOpq0SXaMaJHtNotUxHr
zZCfPXVE6ursAZleiHowDayetQzn4GgaxEoNmdpsZ//S3Dq2gqGpKmWmyIdYNWQ8UH3DRPgF1Y+/
io5A5xNQD8iuxMR56CVpMLEY2TmE9qEAKo49ldjUFdvemR+CSlCaZoIQlRFOvgEkNbKkzoajN/Yh
PZt3VAIWNNesqqnyZE1XxYavSIVHCrwJhQf8wSy0SfowF5K2Ur5AUqp/QDy/cHv7sF8SMv6YfCAu
mFOsqedxxOZfYk3zWnsufwlqzDZC+idK5SS5FhCSfZJw0hRyCT8bqiooF8AnfdycXOCxQ0VZHefZ
ymdLVFi8RFyi8K1EQTaEmGMLXaAZLfkS3ilCJ1ipm2EVmyw4aueLhB0gG5s+HOIHmmqLFEE2D4BT
ZHYWztJ2AQ+XKw6qEfxIfo3Jonc2SghGPJETRSNMRH0RFbgcl2WgqaCEsXx0BliAXTtMSsZ1i3pR
dtz/nXzORsM6ZlblkQFqjU3NtdG/Q83EtD0Bx19zS9RMJcrX5hyRxLDQCwbD+CT7zyyqDLGj2QIY
AogwRcFSlTvWFvzdiC0OLGnvvJN34udKJffP3MwqiHIqYXKW4a4s9zxxvmmi8WWbiMEGyZkHr4g0
93WDXgo/Mhe9f5x0OsWo4uh/wLtk9v5e0paYI2b33Z0Wd3YkNSv+o3HwRcuprTppnJotLUM0Qb2w
BkZMKVHuJVjylQsvkC8zyYEwvF7NIRcUQHZ5dbRNQeVQxWFZMHzT2SydFiESfRC54l5zQ0WIfhld
wq/0bRcKE4IpUvkv0qewpaG1BgmOyBo8ZsTcUa79vvyf2I4aMUH9ktW33onXPGIFzsQd5ZlFdORb
CoZ09CIEif0jOgWa5M/QDL5okreUTkfAUarsLtgRKeRnE9K/olHbRECz2HIKlkocpt+RqqfcjeKL
E2c8Kku3v7YAIdvm2JwwFFJodMZFF2ElGN6+BAWTVEWtJw97fTtXWgaZ4srvPOv9bH46jIzUCn/Y
AzGU0Yf5uObaITYuHgt9i1mBRiMZ8HCo7llb0cABLcSUaq7uy/Tl6LDzSwI3Y15/FZ5GT2Cl3XRB
o9STQIC2Zz1jJQRL/sFyROo+9lx4yKXHWnkWxzkGb0X+Cb+axWpxpSj131oaCoIfBYk4JjDVvdhP
AFr1yB4AWCAlCi3ogtK/Sn5t/a/Qmo/I+CcLIZFBCSkAWE9rKl6h3ZN/RR/kQlzOyaApgoe1AkE/
aNa+dZ/31WG4ljLIpnEt1/OxqaA9pGVWbKwhN2upn1P5Pbxyah80hnRtA4/klThlE+tbeA43dRxR
zQxnnui9vPr6KD3rKUFOO64mDyosu6aRDX6/zhP+q2owbTayZkfelBwGtx1XAnDloUkb8XFnbf/V
8sjX5eDZmBIgbFSnXyx71X064bJtJ0MUYkCUgEqnRcSAZUfSJhRAFzQTuIJVaMvheykWKpGQf4fx
hzORbSpEyIpQX1jckdivaxC4Fj5zpx6Adk9HSAD9q/IdwUT7eW/LdsEmItRJ/QdzLsFO12nGOaGo
rBEvsaxIgPXWnQVuDgQ2XfckchvzA9XEQwTBfgf8jbgEPzsdT80eyQh0USpnyEi/I5vnihq+05F5
4DOLaQONpiywQcVOl0m0aL2VWHRED5S7mI8Pd6f//p9Vb3DwtXlZx8JvyzaaNDv7JWVicNw30WuQ
M6/z8zffazdhNfFmZ+J7Z9+fEFWhu9/6/XCitYHxuLLCY4KANW2D8odoMRpfKGEGmQ3IOWlPo3OK
qc7C1nlVM/7TowIYtIFeqLkjrjYNaejcOYTSIk78l83VGwGG++Rgx/VhBz3auaghLSBN4c/ytefO
s3VwPR5EfMTG90h41at2hqf4cQQRN8xLCckUtFQSyKzj1Q8LHM0Cu3psUHP3F2a9TGKymNMRymC1
06PRC+SPAuIyZyIXrqzFnJuxZCKT+ov28NAAKY0ZnzMyZLp5yjHqcSuRMXuU1moRENJD28ZkOMCC
mSanOAajoa3uwL9DWK5ECo3wWMCaa+2NEyIeFq408Gz8QWZdGvtF7HOV78X6s3VpMZ/tr9Cjfo4e
OlwPfqaVbUqaUSZlzA/zQtdXacSQ9SDn0NT8A/IzpX3UEEhiAH/MElnL0xhRmN32Sn9FvbyO2sD3
6x46iMvOYYPkrMmmlWRExcq7vbmcyBnZY02i0UDeyKR2TbI/5VTavh1goioKZy2RQh0cW35z2Z7g
kgMfT6FgJMRzcJjrIVLuYz9Dmo+wv0zWAmTPUo3I+HFvftXfdDUg85gTabAIRK92CSvGuuZ5ueO+
+3DVgrSrz030hr2jYVzniC7GMKviGJRS9gWgV8/jVuNGsavlPEHjWHNrH0HKnIl7d1R8MsKLQcwO
C9YJgUUe9jHRovEKyumGJqPBavZjEiWv2ezLKDl9tbDKNbavWiFtQ70IGqzCMy9sddkikrj1Msy1
GyxzLVPz+Skt7hk0AC6ENBx+0hDgiPcdcye/uUWCOllyWyuJK14bdBnel3kkuTkbApQ0FAPuZMvq
1uOmBjmYDjBwtJLIa6MGEo8rv6QePGg1tvx0o04pwFaZ7ANSY7TNG7yZCXbDlcRDOGwRw/GGvTII
Fjs/PbPB2nOSaVuG0JwJuSZElW6ryGE4pYYZrOYi2EbPFdLSG+4sAQ6i6oJdYw/V5o1BxaAAis1V
UI5Mm5Z/N8OH+4kXG4icvpLXZO+NNKJwbPixpCBBCi7H3Ymciql5nPaxjXXV+2UZvryfDQFNWzf5
MXcsi1qx5xlezjUQLOd7V7NzwQOHls0nkR7LKj0q5xzvsq+XsGTXjqLiW0TVNziaKLftQyhDOQPg
KX9ntkvyXnyhOfKBx39RyyXoqod16/EGe5Uiny62g/rzle2UhUwrQ/nz+051Rd3Ddm8lfXWnnAif
kIgW6l1bdZ9y/5ryvMkULtVETzImOrHH+uYC0TV24xf317I3AZi8C2owA/9/pFWWb93Dy/9Akfnt
764g6CnW4JjFF/KTNfBelX3JdUSK1mFSsqe6vZ2WSfJ2MG8d/hLIo3t5J4xqDVgzopmEnIJKmgNU
yHELdLhF7YxOLdVausndFZbnqPX82NSbQligmnyr6JkUe82v2NDSdKzYOAN3dMNU61Pc/3tRblNG
XApKZtxrM6r6V5DEGupdqFeGGPUvSDKZebCNorEmFs5yt2cWV41CVTweu4ly0zU7vlBA8Imquxt2
Gy6NeHTW1ILWfKVNzVgur4nhm/nHg/OQEmSJlklgwLuSHlg9z4Z2ID5AaQ8F1YhuOrZ11pyQuuZ7
4bCCaXimMtzmSq7V+9iYBo12C77zTVsdXggSRzdXKOLkRN917GfrCogYPfIvavp8Oan4H1gvVB4T
Jf3iJAuv0W2yFx0SfsJchRe1ghEZjrdt4ZOuViLw8pGuJ+uJf0k9XYxwAU6z/+jxU3P5TUVQ2pd2
3rPapu+YCLPfil6U0idglhcj7qw3tkut1lZA/SyCnohIvDmdtOb+x/p9cPvD5jqE2H2fQLu9RcKq
UqZwX+e3nq7YN640hIbpDJJuFDcSBdyz3dFmndc7qUe+XgzCIiOHZOZdRq+AXF9Uw/YUxErw4HBq
GJHOkkHGCuAicN7AemTIgx0xDJ2wBn4rCAlsUAjstjJI72ZqW1uKElx5+qdVLjH9qB08l+rqUfQV
Dzq9bCDAlK7vf6gMomkol2JF/aSNfpLTYdndJxlX05s/TdTk9q2n7EZSDkgyHZjq2z2329Reg0fH
RdIu0uP6ONpmYmRbtRUPZgWVNcAJpQoK28XrkMzPmbm7CEQQ+D//vi3/8c/QQZscpX3UR1bDJc6X
fvKIW0QFC3ISBKf0qVMH+NULnkIb7mmnQCGQvS6CYAvOa+kEhuXuaOOuzi46AD1L8yKN7J+xOLtv
gYRDlEeTB+xXcd8jBnvFf8jWWzA020wKSkezUAJGur78nZkBF/MIYW5QsIwzSgZZe5VvMWqW1v2D
w7teF0xKIC8pval0XtcmWRaYpqC04HYdS+rsPgK+EC5NB5B5jGn30GEnRoXGzGPxj+9nl/+988R8
glQQwbhte9aoses3um5VE/Q9RC7bZsngmsWc6D4BDQE8KUvNnJO0IJisAfhPn2+XaKM4qMkmLW70
ZcPD+rShAG76tCTnWgMEV8NqsWJoUUvmjYbCcSUo7Oy1x1gGFj9olnUv1XpXPdFtU0tnT5OxADG7
Ltot0L43S69k1iQXjG54lGBBbSHSh9pS6Jg0UjYNsx+VvbPjJTin0DFkrjqGHltvDDO+dvEwu7bU
GroEH/vb0PqWbKIH50cjkAZZmaFd7Zq7eaucQgSe4zT/c62IzcYwoHjXYeIDpma5fPWnsG1En/5x
Yxu4aui19g7OAAOyqra3CrO8JEVL+0K88xa3Q4ZwAk4l+j3lv3geAIJz+JXETXA3Xt6ir75eMhps
majQ99E8ZDb8E3ztB3zWZgZagPec7haJRNl8yqrTHV9KYxQtyNRKtrpmllFJd4m9GnTj2e2Fgl5s
pPqSsBqzyTrsHqHh6dDodzCwYkmpCHPKI0QGJ5hiFxVabV326Pwl1k+xHsxMxgzr6OZVEbrbjbdI
3YsEkvVt/Gi9DkbOPy/G4rnVpftwcPck8njKzUycqVAgcqpe47oR6L4eOzl/YRFaBzQb4euONuUJ
oVKdgVSskytDQrOYbZ6UrXZeFAGvgFDo0ky+45mH1eLkpaTL30GARhe4miJJZiW5cdc5ozUAwwaj
0VikGW+/sFK5ri5pZhyiuU7ZzriZICX+6dVmt4Wjayz4fiIutuxJE71Q18XMnDBrWHv3xmmgUDBw
5mDDbW/ThHwD8pvW6AccJjWOLXSHyVFP+S9G3bgiQ5B10v2rjnsw+Fs62C2ER6BLgjSvLYyCAwWr
2HNBxYo2OpfLkcjQLQeRWz39AhezZJn53K51JchwiRB6mRHrdICmN6svi7pbpy4/OP9c+DhhgYTY
5zrQSWDoN/CHnroYHHh7SpMuNTkKS4MxihUAGaHL4qAqWdxQBqi+W0Lo6ERxh+mg022+vtlxxmqe
hs7bP8hPceFRm/khaZ7k3xfYjhgiEs4xqnOMiNiYMugmyujChS07I4W4n2hubkCH2pnKaYz+q12U
UvvmyomU8iqim0ydszXcBiXhzJxdAFkJQQWJOa+lKU3lYZoJn7ageqQU+7d0nKGoDKGVwGPTlKwY
CWxA9sk71JfR4sECk2QJpVscIF5pSMkdL2Az4yAtxEJSGhIK6LRGd+BeXwhxeDwdEbYMAPS1kQ5U
76feLRRbHfqG4E+kOxxmn9rWCZLz3u5hIbSQTkaHtDkOWMtwMh/0HKsK/syFl1jbDItg8ZM1SVMk
6jZBF7MWTJjIHb660wGkFYAM2gksxqv309R7as8+FqkOCmzVp0bqTENkWXfZ3hwn944QaO5uP4cL
4V5WJ9UTDsRO72QKt/AY+NYPNj3+s/S2VX/L8lOZHDHrQlSETGQaif30NAUYClP+iR8pVu2heXGV
Q36WQOjlLlzC3J/n+l6GuMpb34KSh3sOV6wuqn89NlUzRebGJWnNB1nAE6BBVYClFGP6Fiqify9n
oflwSGUcVZBaT3F6fs7pxbrMpc0tIpI2u6qfkiNsEZhJ0YBZCJ3JiMicj/oL5rmTOTDef5tauZrt
7CXnjutELBUQJD/pOLayzTfdjRIaviCxQVBvOoJqKbjHOr+pkN+WpC4dheXRzucFUp7oZ9BAkpTT
8DKVXdIS+JnwvW55hgXDJLWlAtwVmvPkzhyvhX9v9Ehd1wZY0kSH0LcxlIonk7FvV/4MWj4SMk6P
40Ez2oPWWCZPBD5Y6Rjs6LAjh6LKRkR4zGakNJBvHvjpaHthwzHzGj7xx7jPwJTqZhGLNu/JUHhj
V/xv0VnAlfH+YrJtc2nXGldvXCHr0pv2D9pTTausWBmduyr6knHXe0XQW/98H8x/aoWyrOWhqbtN
oUJXseYld+UkeHjsRVg/i04t6IE0LDUudcZDgwZC7+izTdyRlT+1rZryF/dZ666ha/HZIQj2qk7T
84fdkg7Y9v0PA4//+L9HEGgFNZgxO6d/VTE2LfQN4uMxnIR06PibwQL4R6AwCe5jhkBDpA6bOGr4
y0y9uNOv5nCWHjumJEEsJdsM/d+jeO1C2gR9xFN9MlwKFg1DTu/+wsnN6Jaumeo98CoDY1Y0XKO4
Xdgj2QvpL9D5U/5rDbbKD7mgGmMnFHE/RVgwbyIReKCBjEJd3QnHKf2gS8zHdSZT5qulzqqvi8Q2
415tTzmsgqgo31Ybrx1j/9+QmLLe/KWsR1hfZMBVoG3Dleuq1kN58UFt4bCoPeaF71SRoQghmzcJ
UZnn64JTER8B0bTeKwfntnvouPwRVCTjVVntcECDvbcTdfDAuTjirxNgdeWN0QZExiEdDk/XO9sk
PPzmpeF+OJKNU+dstslMs8AwBgG8ZEF99qihAmruMpBKETdguRNzK0lgCeslx3GDsITBwyY9TabJ
KuIwRWirR0V9sFh/rR2F60l4O1wkq1hBboJj1n65Wko0DSltjx/+lf2rv2iZZzgG6XXKNrcgQYrV
uAUZqzmb0646SwDg2Q4GNKwXFbhEB1hXhzUZK4Ou2evgTB7Li045ExzIHaBqmKlNueofTCvPk8cD
R3ojgwHCiyEtvXSjiGsp+sbVx2tIluvC9KMmuN9idv1o8TzimHF194IOtuTttWPg28waasWOW1Y3
dc7/fE1P0QFbJ9NcsUkmx9zEaj2rwgDnVigLjEOoUjjnw6gTcYW7j3mx/4wUg2Rh546e6tt4zQ4+
adQ5tWmEJG/LavR5ODzqmZS4CiUoElMfFRi33+zRQIokzP0VWoOLSmhneBU4Sn86gL1QXgr9s6tg
6WVs8iKmPqhpTmK7Wvlkve9NZEbxXAiR2gSqOAN4XfXHxf96bmarPv+cNQybWwJIg1WEWLaSR3Y3
vevTZangjz/plHQ8VsLRzDwH09nGyjFXCAE84OQJkYy54gqGGrsJ4bO6za//1O0T3ZVW9AmWl6ho
aGUnPSgi5frhjoInMo/sLQ5/+DNDO+8QQBHWl6ybbh3PLSx61WZjqIzWGEUVWlLV/ZPQKyaSrVdx
0Q4XkMEMoNLs5OOYRuJrNy+RVXrzmUeO9UY76vjsRBxem2PGFn8qmXkYEAn+XfRi8K8f5CLKrjow
9OSmBijiHX8G8O1xQAcMpyzGExW+74p1deD0z3uvA04aTbdYdJ9QaUDerz5T1a2fKQ0wi3taUOyo
RXLDV9Icq2Ap5ySqwAFs9Up0weRhET3Nj7xRTbK6tvbBeIS/MRvo4izsbBFYXQesMwvCn4cjDKHt
Y0w/1OWuQadunzTDe0nqBOsmAKMBPUYAnxARvFZWDIpyKWn5uAcDEwis/O5n+MSJRp/nL9FSMeEq
GOrdxkWB6eiWY7g9LpoSrBQM8lF46sWJ1KBtUE/oc9pD2DnoybML9Ich6G2dKIEnc1cDiwB/9Bry
saORP6L+nKLRqSrt7B4DjnqZwonkM6Qtmliv7gycK8FTNPOeu3WtchsuWKvO6ZBeohCAlUZ6U8jM
HcO2UH1CLcwKljDy4HYeQQToiF4l+/SHsw/otCRKdfwU5hPn6idNyeJ+Y2In2DAMdGUmw9Z2/6nu
bIKP7eKBE4sknxSxKYPNrbaOEm7lm/TeUsPOUGW03q1jC5y4r4Ij1WkDxYy8vyT6KzDcl61/N/F1
iCPYHcRwrrOQjKvyKE4X/WuG7R+tbjnh36txlFUmJEvfRof7TuDLUnK3d1EGuKfFtB/vpKRCIFEt
EtMAFZDjGXIAcSb9ThWbcIayHA3QVRBq8pD0JIBJociTwUUBAPfssYbMu3pcvjNFxh8oY7fE41AI
gxs4P10KcX4Dpay70cXMOOyI+hyxXWI/SmdC8xSCx6Z7Wx0rJCisEpH8GZ2ljPjad5Ez7GBNN+75
u8yArmyDWxwc7871sbUP3gF9/r16KTxDkp/nuGc5UeoiIGtp/NAJZM9sHBXPvHdaSbX1cw+kTHUK
D1z5FKbozwTMysfpFyiSyFSLFq+fbunh3sP6eZmy4cjoKnVlUx5Ls9doNGVe+mHHpvbKQE5Xdiot
gbhXT2UiryXL8LlWQGHk1D5NK7VmGpxp8P6MNag1aJ3PJWrzvWqsq6inCerCmB7aOUb9iZ45IS7/
eCjmoacoKgVoiUzVtRCNsWBHTy8Np6CPeLGtVFWgMoeQ3W1x6LowP/JsDT/ZUKMhM83lir2hLF6r
wdweZVQA+EroKTHw7dWt/u93OR9o4wGE+WVjpwLAq0mkW7riUKxZ8fS1HpdVAubvyH3L2y09Pvkj
8HP3muFN8yo5scgCxQPJoO3PgjZLgFcy9JGVev15VqzaCUyT3S+OiDjdDMw+idLPGI77UKkmuC6L
nRMJgw/u1Mch8xwdzLmIVmApjQfsOko1fFHHGRwnm2Td8WZyPbOPQVqOBYYvGRw4mRahBKKhoAaV
lYl/I/whuapzrcfS1n2C4E88vQI2fViDkSvRsJjN3ekC4cYgpVLYy/hHTQpRzNsu9QAvBuyx8Nkm
DJ0rJ7XxQmxm/Qg4kQRiiA9hBe2vvhfU1GCeHy3PRoFxeOVUssRmwqHjLfslu0Ohc57jsWS8eexM
wxz59QYF47Wh6D/cAhn9zYZSo/qGrKL04OG4OBVw6QMww6UdaHLd3M7DD4h6OVUoqmD9tK4pTRYW
pBlmgz8Y2cpO8/OyuQGyuOd60LbevOs47d5yVDoh2Z6uEnJas9PFvsJlq8iDZPVn5fEUkhfyXSE/
op3q9IBQnGutl8JDZNIs2n+OBf+VonT51kS9T+AAIwgqirWrajQuJAo1dxp043d/6ZswtrCZk8CZ
0m95zWzvLCFUcRvROqcWRzqzOzxHc2SvWCBEa0Le2px2cEby777GCAuvo6l0ua8NNRpxlWuhOGzp
bw7mnunmoaPimlrMOqVFeZGn8MkyrY9TJysU5PDZeR8k/lYo14c0LaRNY+sAllNY5vwOXeRaAAfB
22PUObNXT09ZVdZT44Vl9kyjFJ7fwHCISinVpoT1U/J5n11NeuJlDeGQsmd0R8b0nwMosZL82sXX
WkwN+CGrFTOt4KZnwguY6g5uTJ9vhYcH2wLTkw9ZOYQs4AWsAGRi6FIM8J71Uj3gvCXSaG1hAkbL
wxgHKbtZp3g/NvpmpEEme4mlBQCMqsmlB6DVd2J/C/swEvhh6HlgQxIt/hEi7rQSTMDEkkzOUwj8
aNnvGwLJ6VUmyS6968BdZwpa8umbjECbKTrGy1YYp3gbQNDEeqaV4x5sCXXMerWprRLp12SSCjbn
NCWvUIEqBEri2Oc5Au22dmBpSoEYRTw/e3O1VoJyJQEq4kyIbZ3ooatk99fYOsvvwT2IQngXTYz7
UtDStQWTSL2VKaCeCZ4Ly9KS0pSo9TliETNxXuoeTxGVPUIV0S82JSM+kpccwXrF3Bo+mt0g8YGy
Z8VhSoAfCLZCfcUYGekeaQs91drqdUgX23AjDumQgxc6QSxhCyDaPQtQDdMXltG9zk8cDrs0KAk6
sI71IrYvY1FCsQ3HhDvQlKD/khLnKpOY3nUKrgtiSIMJCEB7eGvBU7ZNp0eWTI2XgBcGHN9YHhRb
gKa8fVl2QvFICtll8z2ym8RXCNTYsXvWHQpUxVkk5T1Zoel8RDC3zgxuvEPn7iKqauyeOQXwwA/W
u/YZ+xIhYcKGd2DpisqFWLRJSYqV83ysvV7+6SG9L6cS2w7YSg/u7v+CdnBXMPgkaY58ctuKfS8h
eTPwhjgPL6k5xZMyxlLxny9OmAj8VjLAGEWwQF81WWN54WMYMxkm9rOf2hiNhZEJ6OhJVn7cwmNR
PAF2WYX3+Q+IvNkDCXZBXjEkFsZPvbWozp6sqUMvP37EMju469v0XOH+3xmMxUFfHtb++4FQkTz2
sO7eyxZJfNyIabaqsMddKnAaELqbON0pwTs9Kt7EnThhwWB3XfHvStSztHQzzQGpy7jHXT1/062m
zpTJIbGNg31PRmxmnpPyovlYswv7XxX5r94cJtuVAx5QgXJpYDuNeq1xcYVxUGKKJgCGiSog+bwu
ilJFSAoR/4XQXHH1B09CJW6LDKSO8aNCrWF2MMgtMuLF31u3Ya4Xf82/9/UDvrQeLyr6mjAWrt9W
SQ7wTcxOhYuP3w95fjagzig9BlaWr0bCw/EJuJrhh2v9Tf5wiEmg+mFDeQ4vdhKOpoQcVInVBjv/
ZY7wN1NhTQhgA8Ou0cIhVA+Z7okMrA7caHAITzoA7lHrjrPZpI6REJuYhyqalun6/2birA+jHhF4
LHpkutal4hP9QfjO87tQFVtyIukbDKWAQfMf60L2pHKsUB7zSQLYmgU6VxjHgN57j7wMod500Qvi
irHJu9CQPTZGQcUSOssFFsKwUswh1PpKbXroAM/RP8NbzYbwVufVIYilrgsO0T4gQCPDcVszgPG7
jRAcmSk4iy39opuyZ5vXz551VIfByshs3iuafXHCyBt3lc/zYm6JAznOYVa5yUkW0doGk92qwgFb
B/AFwBOxmspWOXuHHG1nHQxajt510X+8l4woTtJF234Qjzv3NRgLWmIznCzaS+dob1m4dsc7u6V2
57g4SHmmDvRft3hrTMUdJWa2yVtU2xkSqVxpopalLhpM2h17sujtt1zXQNutBedg3O88hrlpYZa9
uXEM/9GwB2lAoZTeee6E15GXDP/eHZ9toTidNqkeEh97qPfxAGpaItWX8YLFhgexCF0LMf6mKcPF
mHLF2phsuCozn6yNiSHVGdiJgMQRGbZndWdKwlGLd07Qh3xvfGCOj8m5W36sXQuVjHXp4Pkj2det
G1dgNKEJ0v/a6DJhpdLJkDkGf2rNkYbflUC0+bRpr23jCzl8ps9dNzNHPes1h4beCGT9cNOLU30l
djEw2uzi4bASe9TvJmFa3d6dtA3io3f9ls/vWm1QsHOW3+i0+buX9mKGWA8gzpz14QtVFwZvY6W9
XyyhXhI0M5ZI2DYcQPXd0a6OhkYg6Kv2lSIuTPB6PbXJiTsRG2gi7W5dCXsCzyrFAegR1mHbEomm
RXsw1WojiAHEVeznNhfPAceU9HhbHXMnHOzE9MVsBMKG5giSoRTQthXd0jSXh1jA3IIxYth4EvRj
J5yUSIRqkqzErbTWrFXGwOpVcX7T+o5inDk0rwhUluQaCBvs7EEmI2q3i63e32afGtOIUV/pdAMq
BafHw7W4dNL4sstUMBfqQe9kLw++tfyI4mSYos8mDQUfPxufneIL48iRbzxcZZv0HqUs1FHjtU9C
dwYskx1ifwoefDS8294QvRUzqj70oUjwpNdRtAuDtTC5jQIeo6ETDn2BU7N0vGAX+lOy6s/AeGyO
T533VJkWjm8eLm7X3whgf1GAC1gNpic4kh9muO8isFvZddoq464C3EfCn8dLCCca3THAoBWNtgOT
t4Fw1vSbMiPnQUzBk7YM2uKLCvXWe3JpMAYUDK5MjeNSBD9AjzsQR60BrKTjlG8ce43AL6PwHmpG
HgW9dzM2bZVzeDxkKe13d/rWwKAg+PQ8xSTrq0SIMpgNbOcEw4vpm0Qp+SIU17fvTmjVmIa2030j
v5sLCxaqIjkSEnHTOR6wqNsLSm4tL2hgRdv5/T0m+XlxdtSSwuaZY4vzltWlQ8WAAWv/HQlmOobl
RFeqJTLe2rNDyXaEAcqH79lS/1rEhvcAw6pB5QiKNWmogQibA+rMt/oiTd3OQk/zZlvKcmk4oZqe
OrYJjmTWziX57HuRW/IZryVsX+yIcjA1zjK+48CLDAqks2iY+Y27UuRYmJnh2RcUVeIjL8/JlZAN
CsqZcB+qyKIWe6SWB4GPtgs7H0tOn/2YuO8c2I/7u4X+vCkRHXCZXwm1vwJXCVi/0eNrjIEl8vJ3
L/GzT6aqo3P4u5POvAmWxjyxJ3g3WltZIZG2kb/pQRLo4dhQ5c0+ZlkI6Z45AyyRPOHC4ZrxYWAx
g6rjazGpMOvHpG4Kp2mEPLypHB1CAVzqtblpEUY1+Z+sm6rtjavL6rxEV4w4aNVLt5jpqAyuaUr9
0jKuY5pSD9Di2jTmPsKzTpIsWIAP1WWd9igVTtkNcEbuHvrQMNps8s+lS785TBUNevgrZnEBrqLP
lCVvaz92EKyzZx0tEy25ASBSMIesx8hzDN/o3Kl+lVvzYqD6rF9+PaUVtJXKVrptQBZiGljIq/Sl
XbIDb6udjqjJ9I6sGhNI2/fsiDXkuoFrhLq/xdsK3epUTHm96CERG0Lx/tm5wHgpkS5o8Yz2GpAk
Xg2i8tUG7KNBy1YeGyDiyphxU9sarRQXsDLi/63ifmYmrUNTKYlu4C3duJ0A0MD7jGPg1FQyKHaN
zxIs0ZfU2Ql2+F3MB/ZXRdEmvc5esLQNGYqtbK05TWfys7YmT5oetesqfg7c5ZTPYLIxjBK5ZEFQ
khnpBY2/d9vtQiB1dzJEJODwtS7bEt5XBoqHQoaWlGwAGcLlZZnSTpbQ80lmHa21fyaEP9jv7vNP
m6kGliFg8fihrL+9slOv8KJbxhqtFxIRbD5q5ZJwBs3bxlMcZzBUvg/0iWt0DF+ZeOf0eChXLqVp
PsDYiOkya2WQaM3V7GeZN5EwOFRqHmorgqC7fT3by8zRB8uQdYKo050144gg+TUPSI6sYQYSIAFS
8+Pm7nkUj3nezIzmHnnTWvjXO28B0cWsHll6aF/2Zcczo2GGSojg8gkgj2ydJV0WC/6HnMuV9HOn
LeMBYV5kJUpTnbLel2i8JzwJNkJGgkYcbOB4OZduE2Vb9TIMv5cG09XceDN4h3JI4iyr0NGNchKd
Vit1FDP+51Tzua5mmBFr/EjGCuDABXhaoK0mvI6MGUbtS5hsBHFQw1TnXIGqKWpVhrVolgUBXReF
H6kzdIvH1yZ5UGhmHtKI2uiOvn/xFW8wsdL7vTurs7ETpo7bU2QPiY4+oC8sSZAA8lRTKyQhLbBD
JCeChdmWh2qOmbkA/jlr13M6CFysBYDnQmzMqSkJ0/mg6knGsn1VPLEaDzgB6AjEgIF2Hwgs+DaG
fSqD9Bz6BzaQ946y2DdgNbXu4070B0GtnIgl+NDdu51nCtSlV/JG45OHuSYd6aJPr4rDNqp9+aCO
t1tl5R1d4uIK1BCjUrebJMsGz7jjraHwYjzD1q5vhPYPjcQ7oG8J6y0ZtrHnrOmLLt/XnfjvuWv+
RsNZu0I3I7eEyfuUhj+NdCkbeDGJTZWqs+NdtLtx6j8suRXIRm4gT89JWxdc/iP+mKVX81FExu10
yTq4BfVIAqkpyylLjkYtAZ9O5y2LY+3/rMj2Nk6ECg+BhsPELmLUP+n9KJ+QfSFy3DpSw4CVVHIt
+8saAbzry530x2/I+5ZDgbTWPut70wANiC9bgGg+rLRaCjh4FnqszE8Vw/Pl1isqiV9OFLlVGnyV
AQQS0vXx88fvRPFv0hVJ5AJoIPJ5XwBW4+QLuwFPO5yn42G/LTFy1Xc3QsYr9jUoRa3Q8BdOJBpb
u0YRv22+PmyVfZ6La9rRV0w0AA6TmDsYhsmm1bSsH6NwVW0tpYel+u4o+OZsPB8MquPEiOtWIRg1
g6qq2QcwkWHmR42EBew9UkN3ikIpDICHmKZRzENwRREo0669V2UBpf4njiIWSO9bwGsZPU9Cjv+i
PtXX2t1pyoPFZFIeaJKviO7oPWi2jQ/EV7ORI/A5QsRXp3x0YV+JyhRwwsUwWReXFM9A/T0YF8Pc
q27i2qA9mYtFyr0Gcl8pLCjG8zUrgfL1VlVBzxsb+kQ1BbWef4392GnzZb1jd4tbiHMdvcxJdCQl
ZgX9JyeSFmcyeR41TeEEOGgHDGUQft4kV6JzWx6ssta9VlM8EWI7ANyyPE7qv2dVSlOGWkE8Xi5e
+IDEnhDQ0c5oV6DYdIhMtL72M0qa3lxPaJfRfCS4EeMZMj+dO5wGhhON++MGf3a/TZvVc/UbtMuo
cR3HLnoX7npCvlfrSWR7rIDqVptlggfkAJ/uCtbCKHlGjUUrFejl1IjeYyQCXCSKLJxWJs89Clbj
vWFQXu351iPZll5fYK8Qrp/iSX48iTswHxj5x7qNbYBR5x95veNzgUF73b6tKc5AzsilhRWal9sp
3J8106FdgPqQ21oQXP90PeT7KhmRoWjAwAGu5cyR3X/DLfLQep1uUMW33bklP32mV+lqrw1fZvZW
kJ9xwrGCdQKnEOV7RZKRD338yUZhqSFyWZ//Tb43ZUg0IGdLh7vo/ngLfiXJckR86i7RY6pzTDz8
qucClcp41CBZI5EOjpY+eYo2kpZqCGasrLj3LX3YgAdh1pela2vyCNYWVa7IIV8Nx8+I0De9Qcg5
XQnwqbrb+9WpGMntM6j1E6OxZswnGALPPuQmpeiu7CjOC+wBxw2jRnpXKmbymjAgw7LbV/4eaaoQ
RvmCahHiKdnb9eammXmJld2vP/WcKBVoygK1vA4HHCpLF70lbb2DwkjdXTWlJeDK5JaxOaWRRRGB
E7Y5Rk0tckaOWYhX9ON1vPhlVJMbZHaqz08/sFpRTyHZ9XY/MUx2bHINVLvRLI/okQBS906U1/KW
XlmQHqMpWWV8EE0p7Mq7dBLoI/09O9sAiCZvM9i7itt0IMdXq0hSXQ3X/+S9+U7e4BWnJKz7AEEs
4Ss5zQ0TBQLklvjJ71pLB6ZgEUd8rvFE2gu5oIRbEguEezrOc6NcmDy/edrKL+ONRW+eSfVuAeuO
dbj4TBXkfqXfX4sjUkFxkWz25+FBcAdDLbYCwWNVm7481GuKnBe/X94mWPdeMBtzXcWtBcs6EJb0
5AQzU34v9AdtcsyPeEuDe54e5Zpjdez2GE2JLlEjwhz2HCWgug02gGdRKBDew4NbXO3/5sCWoMvi
33k9YiJCkcboeQdDh4IOOGfnznlmb8xuAM9Sr5dXn9cSY+UU/tBbLDLTGcUR9fuEqvFyZueAPgy6
3rV1x4C397WPRFzj9ljwd3xinnMgz+3uZfEta48mBmDnbv66gA0EjvoxrrWeuV5OOiX9G+SOhj2T
Gr255ba1mrB2JnUCT5L56ZaeZ9F+/1/Jk0bNqMxoTGET9RL6QSqe2ib7OHo2U5umSiS7EluU4mWi
6l1JFIZtDOlFfxSGWlRi+kS/uzXhMqoCRNCSeOEhrxd8fPPn1w3A0YMJrLEhxr6Izx3rmTIfx1nM
FtOjZfZ/0Xj/MqnoGHDy65yGVaBTZu1aXu2fZ9B9cBlHhI63IWNS3JkyqFTfDmi2i0pZQXNuns4k
bMfYXr2eHhazIGjPZou8Y69Gtk8D2HkFXWRm5opMxHvxEi5PSyUgDLBaBVTH0VMOIgw/+BYNYgX+
fqyqqgO1P7dNRzZPhpJYukfNPu7t1R+O1ZWB4UHabW4ZCr4wBo+HXOFsbQ4OVqufRL8vZT2CP76d
69s8tgDR4ubmymdxk8DhCcfHghGh+zOugi/KWFhyJf0G+JxpIZB915ehbO4PLHk4emylKijap3OZ
1tbsg6EtW0uA3w8/9iPpv8GW8SWRgubLu2FsrMo5GfgBvvK2T9AXAUHN0iXBdNu5ETQh1Jwo/+8M
WkZtxoRLlsiej+lYz7XFqiMYKYX4oMkkgu52oP1zN+X+S2h2xYRYYbfxYn6BhzdaGfKy76wHUZGS
px6nEHwRDXL8W8TPfuDwl+cg/KVOnT/4x6Gl+lGc4AB9rwyntfJEMdcpWL6LnIrEVsao7fVAg5AY
jB6WSqHgy2wtiyrbAUmgM/GXWdRpqL81evutKbhUjZYvRix6j9D5aaDMYMaCiQEqgO4njKWw/ccH
optGeY+7lr2Bj56h2//IWtoJTFKA4795IlMEgYXQCnCD97UJqprwqSod8KorFsTU2PxLG5Q6Pt/n
AoCJJ4S7/QkhCJDbs2FrM/k9h3xW68OQknfquEgbKFHEUymb44rSGWbUD5/kHb6+RBDEkbXBN6k0
lnt8o5FueqL1iP2EdE6LvzbNNFlkkK6NCtDD6ysEAcnzBmtOQexeXXNwqUcjWp9FeiwhD2C/wva6
y/iJhma/icdsDROi8iHUPJX5Wz5pKKFhS67DGV81gZe4GWvaqN1qmZ6c+usqJfWrOnmRPiBIbAw8
3MoxYbs6IQr+LEYkCIGWV9ITFAw4PPVaQN/J/8ZQz9w0OsaMMShnNm3bEUJzoJYMtBZqOLXxmDcy
/zvdnlQPT1TNTNhTkhWXOFT2W4tSRVGRXVfVhTYca9zukC/GnVyXJr+e7ENQSELZaRuqz90yewhP
Vh5obFs9S2h/Uy7eklEmss6aHPVSHhCEvaEw4odFw65HZ8Syl6S/+UDobn1OgnyOUpzvi7zhQuDb
bbtR5BYyUK7ISYs1bbo4ulbob9lplF1IyANPFHeFOadEXB5320B568mf2CijLBJ+FwVkmzZYSB7T
erUuJltumq3nPhGqgvWOaBd+zEWN+jy3gjzAfLwrxn+azQJs9yTvhYfmOsIxD/z4BveDQvaYmjSP
gKDe9QbFAeDpbWXPTl5BPpiFFp6hDh5VQFTKr+ReHrIWVdGdf0ufJbKGJiBZfNBxdPVtaq8sJYdY
thgUkZEWrmNsnJARLm37+W9+UFg13LJZt9c+mYzq8p3bbQQK9kfnNE+HkoxTALyoYtwCYc1DvWNC
MVwxNJvTD/gaFegWg9zSP3wNDkXQ74UL0O8fG07ZOckeGBSz31AKN5FZwP+8D4JpX+yHlEvZsECw
61GkxXWinmonLIU41xEj2yBTit8ngzPy8SLLAeBVmdTgWRaOwxjxT+ck8OSQOwJ8u9ProygfCujb
klPNVa0iy06I8mLEhv5pFN260ypf0cigX/Gekk2yzgW5zfj0MVuGFeN29VBYdj2zAmEk84mbnnbP
9TocbBj2dR6Th5xKu3zfkXL2lQU5Pxd8fEzdJ/goUfJpiYAdoNOms/JeJKBtEg4LlnwC+PFIQn6E
Ej0N1KL8BIUu0ct9q5AuZm2agQWUo1yUtx79Tw7vlvXw1zFGn7OlIV5Hqcf+0U1akdbCS7AVxI1o
qsIxco+YtOOwMsfUu2NRfV7a2iRRdwPLdoVbZanYAg1IekqEDKXUdNsuQbXCZ8hQOTeLzPPV9qMA
8vq8F0iHYt8vbbt+ZLzPVroWdLkjRjza4zQReeNaq/PM7rK/Yqpiw+THCDaI0LT8hE6ELYFYkM6V
m7uYmj4ROFULZ9UTHq74z+rLvPkacVvEIQM7oFoBwXRtaXzFZybbMrL2daAgYQBWlSDUD31JFzP9
fzv2m2S+UVmIvQ6ujkIwW6HbLFgrOQdeMI6uR0A8M9f+YWZIjRDUYYOlIWGjE71zM6aUXAMR88C9
eHrYUbmMJHqyts8dF4TYNlrYKYPYg3OriR8lmiHSLrb0Qimn25pnh7y0vXfCjrTsl7Zq/CqfzKJh
OccVoJw15e5XJWSSVtehNkjcJrNZwVMW7MFZSvvEk2juhBGrwDeznbmy0K1SN+sNieXt5hfbsvyQ
tpe0PYuW6uVN5dbtVY6JwRAG8aoWJIHrOBS1QuS/Eml1E1lrnYU/2QLX4w5aBQflOtfHghWdsN6L
L7oyQ1Q/gA9xb3zlhJiIAf5+OUtvSeHiR6o0JWACvXhosoxcEX6bAhaXKD4upc7zMuW1NKNSO1rK
+nAWO2Sn8g1UjudDu+JTztPbWiaUkTFY0+gkeL8SLu3vaaaE0oHAFqLp29Lbf9lcng4Sp18QHq4q
p+JqcLogKxsfVkE4x8gzeBUBJ1Q810YL5TPITkR3Sag0VW0UxGay8w2AevkhLgPGEk1q4S+OwMuM
BJ7tYaVHdadgqySDcqccuT5t9NlMZOAaFvfmZ2dVl1C3BK5Ae5jEWDpV4s/bwlLKwltMDddxPS0G
oVjlJrFPu3Hgne5iwSGPBYazk0n+LYYGxNQ3Hb1mcd6pcWm/2QJ/IZdOBP380L/EUb5+x1H43FsW
ZGxjioEbxf0GNAQY4lEf0HTaM/4b6ONoDOZDuPqY/5rpkV8TByuqWfFrLnGFAUG830Z7jqwCXri9
M0bsHL3dyoCHBgY45Y9Si4WDBKJQdpgZfubBsp46a2KMaVMdZ+WdC1lsvROfkY8NLO5x9qcZFfKt
YGr7Wq2bClVAH34RWHewk5ITwTtXwgwjILNsIbiMDpuAgTdw1srXovP65GJGDn00Pq8RiNWImK1K
fDvWkGrFhjIVJOcF7Tdyb7s9mwIcsYXy0N1ZOKVjfMLCFkbql5yIfRDxe6wrYiHzea4i5zEG+dyR
bgMZ0qm4E0vwUvyZBMa5bpWVLPvXAkYfUSVPdsJjzKUTVhywpLAnINkTQVpUsPxNsVx6bO+yjFag
WdWsXfzFVm4D73r1vB4KceUPrXVYQL76IcGmE9VX4jzUD5bvJ2iXdUM5fzkfhx42Mmj29FWrzu9h
ZvdpBbks99rn0h+DK9duOju7HRpH6PvJM9yWiP6akDrJQiiFMJXuLeaCXLkQiim7RO2nu7IiGZsA
/3DN5n+AecLo3QDAW0vNKFulrB1jHgsAO8Wrydusrw2snaJfqwf0I4QAK9kGhKN7IT0SL2Droq+U
ktUisIX5hN0Xa65H2vsnIh5ZFXrsuOseGM3XVcHt+vQv1hCT6vtEas13qqkywtd1B0jwi/CModl8
EckH3ZE5EAYTncC102jz2oosK+5Q+Edab1dv8IUBYKF0kYLS0vx76O/6rHrGVft5ebds4gX78P9N
8J/WJYJ6rtez8Ql/cTV1wqhu5jm+ExeTBX6RiphodaIPd8OI7Pq1X/KW4jcx5bLMH7UtKO1lB5gk
OLYVpoIs23YxMmlxkfxggUegSiYazVos+QNLYkOYJgbu8/TUG/83G5AmGdBkFUBEVb/gFfYqGLcI
hi+Zdf6Pc77r8/1cUNerW2ei3vpfZeASHBfvymZNErBa6RKiRNAwVRJiz/YqHT8w+yYSb0K3pbTD
y2vlijLOlhzntmUrkVmBIzPZ9HTe/sGxnRvxx737GncMlQkh5C7h9SDqOJFbfVpL2SUa9AqBfuN4
Zu+2szqTUaUBlgYwzc+19q2ji+q2UNgJ0+eoVSMUUDXOUwaLXMKR0Adpx3869yJheTe/ltl3+yaK
POy8HEdUnMAvQGyzt8w+pDZsh5x2I1IAQMdclHGBIBtetf8wsrmCv6npbZhwzXvENCFPCMWTOlGA
M15GNX5lxFzvV/Fg2LsC3jJmxWVNZPZ3DciIkTg+FcOtos0gN7qtgCgPYsLRA4jtwkC9KJNLRpQE
DsLW+qXtk5hDokItGKqofBJFmo9Sba4PklAwugRm18Ja0+MxAgrcPdoem51QNpKh8Dgpuu60VCI0
LwQRK111PDiv9rqDVd5xNodU+1FIWsO0k7wj61+wlvjtiAUA0kTWHrD2oPs3Kb2vZzN2dDAr5fEN
SuWUYQza9/kAGZdr96Xn3D/MMztVZQRNRirIF/fkKwh+hJWzQQKZnzBKlmJ/iNWoNI5ZgvaGiOfz
viW1zwwx8g7I9ye7ZGpeoWJU4EvPBiaKRU7hhoHi+85RBT55YqqHCzHSf2WOQYram1XBW3Pfh8h6
spisIeTLb6KOmOUAGgsmQNQynOZBGa0GAdLz+Ezik+Ium3Sf/BOQsPR2sxB+F6MOPE0Myoh9QvB7
Q48K6NLQOgsnzXQtTlh1YNmO2XxYg9IG09GrHfJfpK1I26ToOWwmQrOpUWRfnXkSoMMHGpWz3LxH
KnmIxnJclaXsYWWLq1ZUgVGxWHfsIPkY/inbLKByRt5A86LtNiyhO/NKasdIXWrIry6liUqygSNv
O3Oj84RViCE4rNYtxbeRMNwioA3B57uhu+2yCfXee0zo35hqzN0jZnxxOIbyamO8tM1SW8OgwCJP
7uMQRXEmmlx5z2NWw1YT8GHyIymHcxOswj+y7xM2Dm8TY565bP933jlJ5uw/Rdymjxye3c9OAJxj
9XfJUTJp4rcb/arVNbWnZhNDHoJ2rlGxpo2igua8RpmieGD98ZDE2HPwTOqzR8Im2c8g3nVDmgnv
Fzcmc7fWOhOeWDIZyW3EaY2AobxLmfrqd/iMxxhUOXi6HXdRIjuGQFeXqcLtGAoF009j7I1zJ0n3
NDABckti3m/zQXqIhfZ7HdJD9tMNTGwcWpNfK7QYG2TAWpHI13JkTIYP+rSoLVnj5oVpHskOeT4b
CeGg/H5T4oJlzpBfyTp9IqpalzCdnCqZOaVOKYUrxmtP9sye5OoQGrV9Ia4Iq536W/yaxBjUf38F
zM+XfI1xxXyL4Z4aCFJdqfEiQcR1zH21GQu88L52em4rlopJdjCl+UE8kvCSlNmH70ICo0E8ZJVM
HGIOeh+gxfWezOTMuA8BFfZLxIBFdhp23ASO7c/4m/9m9gUXaqImfN+Q5z0utorSe7ZelC9h14FY
FNIVxwNzWx5mSRQ+fMiInHlGNV7OuJh0uZmE45mvf1QjLoZ569QqdBFtk6U0Azp4uEpYd//xjqW4
2tOWe2tzQdI9xY2ttWiJt02ZFha+AtjhTYwrEF0RPDGTdh1rlKgnVEkyvEP/P8FoaYTWXcC9qtH3
tTP4S+11JiqkUBkmiwDAwAhYn0AIjsp1f0S4NmJR+kVSJIgiO1U/urJevWwkibWxkuVV8gVt/wNn
fK0HONyrqaa74XmNG9aB4gPwAVVP3c5218UnnYEhN8yuU5LtLHzNeNoSEl2wSwMxVR1OFkGlCVD1
ldfbapvZjB8/4IPCZEFN5/TFxy37lO6xquHl9yB/aPLG2NDLtzJ1g5+Q16ZeLmV6wLkvgaAQrpWk
n3t5ITv6hfRaxffqOf+oh2h0UIc5GXgqdShavUcYoaAtVFHueCXA+mkhBLy2QqbxbueAQSF9nvM4
cSUCDDC5xuUFle8wrHIc0eviBLfuoipifCWOaOKjtfYObTezas5+F6AsPa6lVCiMPiVY1U4hGsdL
9S+TDBwwW1mYiQogqJW3yjn8qObkLOToeEC5Kjdq3jc+Us85r+4fhBmwuiAMQhZNDtubc32X/5zR
OEubrBSjnDzUQJWDzEiavJTd8/TQFlgFnNv2eKo5J7ItW+DO4QMt2bt9sJweQbq0Z6BqPEoi+L5C
t/9FIOQMkkDexSworVRMyIko1GulnQ/h1pZwzhC6TMTnDHvh/d6bz4ezw0pVfkrOkOQN+bWMvPCq
NmE3Kyafxdvo+jxx5BD73IjeXZxIe7v41OvAXZGsRdvq1ciBg9XhfVDh2wTQz5kUvLL4fNjEsW2H
UKnfNkPvP14RIMbEOnEfEm6hA+0CshVPkJShh6ANowXBwr5CVgUlmQlqsktjjb96GUvL8cZ7BID7
cI3HLCvzWrBeMPrDp4RoHiyrx8+QxRur5ppZwCes5PhTHoayAaJcJe3obsHnyQeJm1uUNuPkMzBI
Sqh5N0k+FrxEZQaABj4Vm4p+gdZ1JXJjJVzVZXVX+p0AvS+SHCljUv+Eu8v1/qgpNV1hVemcerYk
UruqTPL+Br+RkPj9ByhXAmLe3eq6Pq4QSYMXFesv5hQ9MP/mdvrNyLcHlWTrGw5/U9F+Rcl248Nq
z7KfzQkLzT2lHHPjB5P8wRxxuGRCUrbcgwYiDaJziUZkcl1vLVrAbDYxlOfDGM/iae9qDtT0SDoN
mkrwZtvjpG+CYhomAxrXYGE+FuKvcgD+PyYb8/lzKTWcaz7Z6nqOjJJaUnIVHT6x0iampbeGc6Oi
GHLCaig6SN2tLcQUz9kLe6auCEV0MGQ5j2e0XxfGastKL6DQqXtbwm+gYBS22O7qpi3BcQnWku+O
Zc8nCg0ud5ZrWimu20Jw4Yc+soitSa6+XyoQviMpdWyBDU6pqEO5wNFer4qT/I5Oy7mhiEWbDN+D
nKWHvleYGOA7ypEriy3hfBSOF6cGMzoOCwWhgbMz7aDysAhyutjLFOd9b0fcUt9UCePzHENzcErt
H9nwOw62OKHjbQg8OesLEGkE/g0QvinNnS/4eaaKCsAqVDh1p9DZjolq6BKNrfHyED+QzOx/6ml7
fAydfxe9M/Z6rYrmg6uVdfjLkbvAaxhS3K4eFN5pALWhisP6SAeiCrAh9HbSAlYf7426YsGPYHgG
YsZ0q9dwK5noWIYpr1U29OH7d5YwJbR93pU09Yg2hGfuPJd3wnIRQJsDKcuoDbQV/x0BVFoH98/V
ABBwbfslYzR8xQbbiUqk+POkBBj2NRIqWddWWxtzoD3HZu3cZRY36rPbtMkvt1ZOpX0wq3vgSlbg
Cdv5H8joedPEjqNH8v0hzj4DWuvLaLZIstFPE7XQLaZmMGdD7stvrRLJoOo+rWj4bP1kJ9o2V9iz
OMA8VrWG2o8a4tJtfZCmnOmWXC2/mudC2/TvxWHYloHc4YwQAR1ekKeMQfGmBB7BC0Ox+4Fsi3f7
fu1tyZeOyvUYsnd/LdSgVGsZ+V3eOtesUFgsDyHRwiEoiSNZTfEWyHqC9czTXnMUgTigdj4fPUKW
muuJdCZOBVCX5qL7C3we+CRet3jvceAyxTAn0Ki71ePM16dDehbnOuDQ/yKXkLuIyApc3nFfOmc7
FkujYz0bGwGAS7Zs3mQtx64Qum+vZC8wD9iWpN6X5FjB/6Myy+cNyVFCnhMaX6hvTAtuxVvmgD6C
KVAFJ3yypC/R2Yl0n8trQV81hPWVI/j//nNpixmE2q3aMGuICvXYDTP95KdBtAzPhv/9jHLwsmRt
0G0gxxlmoMhsadyxw/2EzLrKXnEUfvNYuuCsUBrPmOAIcVhTGvt/9hKXob/QqOBHsb3i45mdCtgz
FSWeSlC/VOjhqFkEuv4pzFU7Ohoa+DKVk/blUFKF8o3a121t1ZzvDOqlmZoA8H3VSh63pfaO9T1P
YPXJRbHMUU2FQcw+cJJ8gUi/MF9nojEy7ILEL0H+d55NgBZ3QfGKtNvQlTopzfdSXrqX3+BekkIZ
dC+/t79aOZgf0ScbGhXyU3YcAHtFcanlCFY3Zj0L1ryxvTgXMkO/+yYtH5IyBArWksudWnpqWw9+
XkbUUxD6onReoDAX8filZwMLfHrSnovibWpqWdGCintLUA70euCrur8ZEqHChpqJC/dwvMizueMo
JwzXGO3HOT9eI6fBMM4MzoSiF6uPdVhGi8gT9PWCUFIcyftjIzIyQt3+gsUKdDTMADdafj7Aw0FB
9hbP91A97wynNqDcZ7+2lR2HS3qpibn6/Cm6WQz08Fr87Yv5bDoTo+foA2VSsHqjN9HAaatGsome
6lzo9BaGlvvqnn9ztgdaXvvBBJtqF23RQgMhDnF/O1nJFV2efuaO7IEk8H59H5UMWP6Qish38iUK
u4Jw5Kmk5CcWXge1b0fUgMm1YcYskFJ6J1YeZ7WsSyhFQDbCEsiJ1YDa/yp4WpODr+itFMIhcvOr
lydDA5Jp1jweb8+WcmQJfDoQX3+3kiEMvOZJm1fdWvl72UvytGeWqtQa+Nh1H+qIEDvTSiWgChSJ
g67Yp7sp/z6/MKmAwXEXvckfCtG3ooFPYobUaULYoaCfrJmDazmyjQCuVrLel48kEjxUevx0pg4u
94eqPk/G8+8FkpYZy0Ek59zC25lZ7Xt4SXuQjQ9m/sisVlekkyhCTgfvo7FbpOpXsyXHFYFp1s8J
q+KTd+mOb91nSVr1sZ4FYWXbSY7RQWCxYEwUMKhoTzDXP+FwKW31d0yf5QBXwvzq8wwzgJcUEC1z
jIlrfOoNHwhDuifHxBJtpZMID8HepoQBOsGgjla5nT4eBNvGY8kCooXGe30kjTEzFITfTpKcDDXB
S5hmuK1SVhqzP7YPqJZULvv2rtLSYbuI/AnpotpZBtow9r1d4hnjRKFTIu44DGfR64o1KvbVXzqv
P4PUqy2Z2Xc1N3IGR+qvSM8nObHzmbNwtGcpv7/AepUfRA6hfqP7SMqr/pj8e3Uu64oDi7qUft1T
inqSi3RvRP3rW0pdxAWa8V8QCCKYqh9V/iGfKKRfiijSzffGEKq9Tkr/VhZesl381uWAz4+mIj3i
aQjpLcYlANRbBCZX+ZE7Q+SnrOxzvzW8Qxvx6k8f+50GBapxQ4flRQ2qQIRSkuybJfUXyNVUQdPB
M669y4wL4oVGZ5eBTDkshTOTdJckj2xKc/CUNYlYXc70r4z4LMmjr2+1ei8dCuTFBKWJLlL7mMkL
NYUrlmqI15eiDaQ3GtTUoEHG8zv7uBy7PO/lQP8fhO54xicss/v14M6bTlQ6aiFQxmSjgq7H0fYd
buHxo+mTRZhoCMSmkCMQS7kZpcnOzRNRjHSNja3eDtgrrwCe7zoE54Rv0aBl/rzFIj/e+uo6ulsx
AyL3AS+5foNIlPeKOpjkO7KEQIPrw/jf5/txi/kDvoLtEwouXupqUzpOWOUnAuBlNwIdHEWxZeiP
MoOe2SgnvL83vSjXlF/bL6IkVmCznNvTMU6JEE3aih7WW5mQ0aJHxOnoa4EMwPraGBrH7LdTYy3R
z3eK6kT3ic3iY4j/fikgdQ7owOB3wnedTYk+bDNbp7WAEHH7tB/OOan5+rdKxV8/xT/9WHp13cuD
W8rlB1ngQ9y18JSDxJaEYVYrMJGmc3YVSnxRiKDcz0IlluO16SBlSdY8PRdQaE/onvxl8NF8nEsb
qICUAGJMKEKn7BPNqS7ie6AA/61mWVjNyZYIFi2LKdn/wJdRAxnfIJXpCh7mX096imM1OHzZl5vw
r6/6Pbm3GB/A4CB3eETm3uSsY1TbPQ9FHsL5c80xegv6ekp76hDi/Ii+rXAQruH2FJqP9X8Uj1fa
jKSZVv+o7+3im1WeQnvV3W5AeJDAeUsoHx6q82iQo12FJ9uUPixdGWOi5PO65UGtjf5t38dFtPpK
zBbYcGo95groC1LUX7JhW6PoGC41eAzA0dvUsYVtoR5MoZIQqF91o+g4Yc2wxvPEd9MBeOvNtyqg
QXmorrLIkvYaOhNl9Fc1PvjdxFG6Gbn5r6dV9ZldO5PCrqmt9crQ86c3xSGlPUZnXn9MgSuzj2Ap
QJh69WepI1iKTjyQY/q2JsWVO5Bko3a2Q3r7eYCd5qVWCYKQS5FzsVNVlqGNJbNO3WYWC2GPhdxl
QKLEhYPpMgujxnYWt+phHWmVNoBjyLF6zqNFmpf169atm3uuEPpIeqWnm1/tglsvqAiTBwfL4LYu
bD2Y07XQ3VSoDlDj5jEbfONgOykGcsAe4L/91wpNUFLyYLR+VgKjv0cKDyIZTAD9wZkjsn4Fm9Jn
DGLx4mlk6A7ZUguLOqXhiQE7fzFxF2nSKd+iFXrVL0oZGW8gznH/C3ic3kkvalKab7Zbncb2BhCn
wusTQWQTxVlkMuUPtbiT+1J0DDWy2rvf+1alRgZm8SbSefKuKvXBCgVOFddzPveEhTOcM4EbXDzk
wvg8R3Ijqv9f5WwgRgSCBbxrJKXRcJRcyZHIrmidLLCWQqPsUNpL1zCo7f/fgTgazawhOY0e1PVa
lL2yMixn0KA/vYcAapeUEjNIUFGqRYB54SUYyT73a0KuVklLUcPLjOkENY35qHTpNYiDNqDiUogZ
asLG7fzGRkjSHNVCIbMOnZUxWEJttt9QdOsQolrZoIZP+Krf8dijvGz9mIFdrwAameu3FOTItc/9
FN63bDltC2nKmxtGOgn84p0b6z9f7UDb+iEO6KOTk3R2GzuL7m/GdvFr83Em/ZSQ4B9g40Kx4hOL
NjzEzEvb/DCkbaWDHMwCT7h6bLYFqE3HJ0oEcsGuHr+hf3jLpLEGLWK2WVM+ZBOsP/4cT0X44vW0
7cCklshWzQmvnhTrCjUacv/uKpIryHqFogZMrpR+IRGOcN1thXjorndTW8sfYVrOfT+D7Zj1qte0
xE338xsCPO20YuGxlI7fLpfY/JEefl0UW1xbr7fXtsaPIWeQPVSrBrUmkvSa5BBUpUyuQhFgTCvY
MsnmKxysiFMAp7NR5S2KaTer//Hvxscry5DMiw8rK1utqAwY5sJOgc+qtbeFoQ6Hbh+wVePnzFEm
K+JfuepMXvNjQWMPJH3vlHGAKg+mgLE/xynib2YLZCdWCvlc8cMiO3c362BRHQn/eBerQLogyciK
RxDAr8sPUv71gtbXWToPBsRrwG0ypY2xzZqsaruVtOg4ke46sH0FPvmxnYd+jaQ3m4QzQ5AVYlSI
xRi/ApIkpli8yQcQIT2o6sFlHZduGwfXYZzx6j6L4lk1XvzV68iYW/XQKRfDy7tfQIgpZxCe+Gz0
gvSXnEt9TOwE8iKj4NvaGUix0TEba6KLB8qbhKQ3hC3yf1Ih7jbAfANxgl38S8I2cvgAmyoMwKnQ
EzUhYe4bomXG7xpJTbQ16CO83fQsnYoa950qKDZqP19cUr5iUT48m8WlBVUubHf4R6myVzSd37LU
PUzKbOjqwui/5U7pFa+vnrTnC4OOKo0Ie6Fyh5vbLOjKk3HqKom2bKLTA/7pvSkKG+Sk0c/7ouMN
I9d/1yVdD+5Gt6tmTCBV/w83Po7p+HV8KYuT0HEv2Ms+vekCu5wWnNWTC5NxGl1J9DB9mKvgTvRM
fqRPlT1sBrLK3lYNI2mOdGCmcgNn+kilDLJO8Ekp/VD9JwgHTNvP+x3oA4BS6f5q2+Vbmq1CcpBS
PQqUz609K5ZBsyYbDFgXQpiKu7xRUrXToj3I/Kuiz5VwsYt8RERFtWFZgpwJ4dM4J6gXxy7u1mdu
FA6prvUKucVHzwwhOaelsvjZQ9cKNgtFKwIq9yRSiZ+Px27tHrbhharodq7aKleQatFhVBHq0Zbe
xWEHid1HT6a6OL7JkRhMgUAC1k/YxUm5CulDgBunJQKIm7Z91aDQzqXjoEuGgitSA5iGgZLs7bNS
FYDdmVBIzjSSF14bnnms1vA9hkjCJ7ptP3gmtLvTsMtrD9ij3451LnSp8+/W84DuKphgDFXYTH9v
PBsbsjOd0xsCoeR2M0K8HJOPt7RIykiwZmrxUtmsUg9eqg0sS5dKreBWch9Na1APvFCwUd/mWMT3
nnkcsf17w2c2vx7wDl1wOqnMsh4vfT+xwmezIprLFWBrjGavgmIItgdS2mksRyszLRI42kTAe9FB
GTXf3uaeGIQ7/e+9ptLvt6LWINPIOOT8RDedMAuiB/5dr3PRe+rTRhYWRAk0DX0G/GuNHPB0iqEj
2lFSSeVlyGp9112stWaFHL/y/zpOhTBXzrN2ts6b0bdXj3XzLwUQMqKx1RslBDxa1TsJLXUxw9gw
N9DYhIyiv0WfWHHJIgXNEmub0nRlIMmwpwaDKtoOOIg7D1ku77Xce7/2bOJkM+nI61PhpUx9/bIF
BWqI90kDBQCPXm0QC8kp85+YnQqt3EONH1S7I/1CKGrdinB+C4LpQrgohl3Mw/jJCkJkfzx5WG4e
l8EXdt1M+135CulRk/MTNNDiflR+YWQG9kfLvbYZG3pelpu1JtPfXhdD244efuFBIup7vR8iOCYM
C+uqQLADRQY8QM6TtTQimLEwX/hgV7vf/6OWNkCZWd7XvUa5MYYqwthxpK9zLKqfYIutz0QavBfM
LV/BSE8O7CxydprYcZa7kGNJpSNb8pXxfkuZpWcBj+VTlQE5CJh24A5XsrxcbODmiRVUXgAQrudx
rGcyRsUKdi3dTLPoUlpS4ubUtF+APH3oJnadMWEuJ8boVwAIKhtIEtcGAEeD4OV8kWXSRgyMfrtC
F72LiGiLSO+lpb9NVSZXnExxh9FemtBvT3RFBJD2lWehugq02EY9+p2rLvGebet52XhUw4ucDDOD
jiY1VNHAtlA9DxrC/1g/5pKn42YhGet03UBNReXroABpoztG3jhTbaZzGUyFC3LZNe4H9Mh/DXNX
hqt3m7mfymJdZ+Y9kkz6aTcC7MQCdNaZVnsuO4S7IvBszyz78K2TQVp7msh5i3yBUI7ob+bQJQLV
iWT8xHPnRc6SQ2BtLiwM/M6I4+TrVP+/TDMOJGV9qqqc5h4258gbCvFgZ/J7uZNo7+DJOCK/zXXx
fmzC+DE8rBRDkYQ9ANjdCVu1I4Ct1hfKWIN7Lj2kIBfeotttZd45HarcsP8x/7USzqcMcgQzkbyz
mPWVvSV9wHpzUGYwP3uo4zK/k+ahx+OQqfpI/nL7e7PjKAQo0XnE+CgcGguV8UT4ft+sZJ/p0jfG
dXtqOHvZz8+vBRvyeae97h6pvmNBQhI+8WQ6dctp4LVwezSpt/5/5nufRJPA/WD0I62kbKgZrc6k
GTQzbZWWtkNBeOjj/bq8rtynE/+a5KVlhtuPmJY22eTbPo41BiJdKA7stFYdIPrQwg63Ai/iorip
NaQlbdHgw8tskf4MEd4zg568i0G/v7/eeoY03TZmSPF/r2Cweg+GP/T8Xd5nfotZ6Z1QnZtd0aTp
qpsVUeaM+eV9WPwxvHfGO3pqKvbAfkrwOwfmujVTFkrtfdnhT88j8MeGGh2kQhzsDS58dm33+ntq
+Fzv5AEg1DeRS4AzezPB8engGcC99CipERsimhIeLUsYZOT74jEnqI2CjtL/d23VX+UKR5rNM8Wk
clrLh2z6iAqHBs3iqZOy0bhmIXwocnIcO/btOSCHVkmfGAr0KwVCpH7krIk8Xe0phJebThC22g2W
+qLnKDkCVlsGrFQAE4hFdIlaJtT+yyCpKo0kp2xQMP1uxpTb6LBVxH9m/yQ4UpFKcyFczmJhDpaN
jm1bAjBO9NneahNB0LJgRxd94tWHuB9WUE0ZTXghj/NSlnbhUfag7QE+ZIZDBuzlKpurIsRaXGjf
BKCOapPC7aza/nXyki2ImGJVLN8uk0RzQOQBrJMkaIBz6KNfoRDJhrtollQnTHIpLBtiUvmEwlVT
adRsqxnC+NUqvT+iGsBYLrMwKya4d0IEcuHSVztTsnbjoyFe2XuD+yMSpxCY6ejtXDft7FkPpEJA
0v0zaYQntl73DZFvl4MXkdI3bMY9XePcaSk5jBWxF2rldb2qBkCgYfhJArcBtG7Ql4SUPDlVNdjD
0xs6UZf8gKqjrOXo82+D7M2P/qxlb34Uwd4h3fcxQ7WqYHZP5XenEZ0s59mMr3QgVRMTcvIH2bzC
h/c6Vc2JLuHKvdtDo/eQZ8BCC+AtWt5TzhiEphvqS+UWIGJv9w36fehfo+xkNiCCvOzZAZGYasFE
SMgot6n9054sT3cYcIR0cXztJAvlw2El6C+f47xdKr9gkf+bXTlkoEQRk2q0Zi1L9DhTiM4BPwN0
3XdzenO1DY18gpmIxOsM6GCSXGJjb0SgPJ504CXvG9FsXRVUBQh0NlQX8xOWCGLRlz29cvaPujEj
QjIgVelytWeEzz3ZcLi2v0iqUiO+Y+E6IktFRfalaYGd+lwhfj8c+FilgdTdjNnVb/Z0SpoE/1do
PYvM+u+025OTON2zYpcHYOmDG0Gk89JyBS8SNaWJT4Cm/Td9YO+A607ASxoRY7BCk8tBsaPUOm+t
gXjOZyODpuicN3DCQ7TcTW3IKUh13YhtgZc3SdNvS0AHRU+wag0vwqdaLcEpEaJNdUSMXzqAj4cf
8ora2p4eDJ8Q60vDIRo1HNxKPOLNn5mBG8X3l21ha1bGqhNmvbXfd0KMWQU/OE0jfkjGxdeIJBwz
1D+8rpjGOh0jN66LifhsnsVl8NYlSGFKgNQqDNaq4BGgO921jhHJJ7KJ2y8iHwlUQTh2JfYtLS68
OhqPnQhHze9vgfRbNtwna9GLm8SsGFZBvPVCg2+QkiUGIPF/3Zex93IXtR0eOGFRx6LsLXrss8yQ
j2pqQKcHO0Ldyql2B5VfHw0J6LY7fzupKei05EHSjCn2Pn0NmMkZWQZtb8GoXogHa8oDHi1YoBT+
SvfWrci1APTIqwzqvu5boz08J60RWO39jAQhA1eeihpjB7JazZZXz9xoZdQrhJK/rU8Plb+IiwfW
klR10n8DeKgkttzL7vj0i9M76a5V2bXD2OF3ad5jGGY/ysZj4vaxyuaWLRYkxjnBnwFJzW/juNlp
/PspgUDAi9QWbP8ZG+1N6VphRsEtJ93WC48UrHm6ivtD8qyvwsQLqEqyrnwlWPXguPosdSlkkuCe
yuxfc9ZBcSW2V5GIQjEd3ydweaI6wsykZZZRQAIM7fD4MNhMDbbtIlj9a/suabfTYHlyKAZUAJVA
W6/H8/4I9TYM3E7aWJX7I8YZEIDze6jeFxypz+oxJPjt2bwJvrYfxeS2v7F8eJojrdAgG+cMg7QS
+ZkY8Ti/qHxCLgH2J9KJejqDIE1JkM5iQgXDuLxl7i7XZLckXKwfOa0aovOm3mHy+Sx8EWQjgmNp
13JTQRa7tcnGzDKqfCTc0X2k9Wx/nB3HcEC+pU430v6wjB2NrSf/FvLJQ4Sb/z568FVndf83bmhC
bijk6xWfIp34Bcjquw9Q0a9VNMSTGT7D8CxdEDbVBiKnYbP2W/oAEuRurSjZUcGMbgU22XY1JtA4
NOZaY4oVp12yGYk6Omhjpb0SmmoZZCLRjHsJ5kbkuPDFAh8wGt4Aru+z59x4k46KeyAvX2Z3NBoN
c2EQPnyzBXT0GpiLoQv177RRtKvGj1I2azrR7eBWTd6iR37NmEg5UO1O50WAkX6gtuFk8OUDWlh9
W27UTxDmksbf6HMKTi1mNlUvFo/YFQhFSpydZ/mR6AH9IDYumpa7HtqcGBl7A5tqVmWWawVWp97Q
K1CIZQIwGRkpVfZV9m+/qU556mwZflw12u+WYeoDnvKK1EQrAhV/gF0/DYLDQS2RfVhTO4rUKE1x
u30J8wk3IxHk4hm8Yft+e8gaqJD2Dbx8wvzHKTxVqFz+vrMcsPHJNeWBj8hiehh2DyHlz6fRlJ8R
POUmk9gr4iDOiQcf1IOt1r58pg1WZ6hiV6JfBGKmYkMpREX0B66G0y/UL1je8t6ErPpOdj1b+eUj
7zK/hCRhcCYPAH/ceCVobn8NojOwePP4qzzKFpQkarhwgmEPJsMv3jHSKVrOEAI97tN6jy/fpIU5
2expm6we7nuVOV5933oLsaJhfGQNlLfkEGXtfoy30GOvaiyUq4LuDlni9rT8t43/U3YwvVFbz4FJ
6WE3dCxDcvB8XkQvLZ8Q+B1F/FrwAHt/wjOpodAIjQLOmRpGnr5IfVTZFzeln9sN3ToexSsUkDsW
KU3eUB44YSyEs7VJ5DoWeKU3MQCjX1eGHfGhOkVJJpBFObLiGEc1/n9WjFEkRksKu1e8GLR8k7s9
Y5Rx7F+3QQamnJanbBBTm5eZ0huq4MRMJbVPkoanRp/031gg1xiGs0U/jtL1OTPtMJ2zripN07wu
MrYBevBkGgdJHovPJa1KIzfPEavIuM1XS1CYZApcmLEYikHB2ti19WfFCDnyxcxcPG7W3rvJGtSj
qIaLWcX2SdHNI7kmNe//lrpB7w/YEL64ksA75zbCcW4qlMk8P0LSWwPMZ7Wb67nGP49C94+EWw1s
3SCKrfo1uzLtBQ1MOPJMPDD9qdLq8MiEjDZS+N4ye6KQSNnZf9sJ2U3TJfcqQj8lcEE3Rdh7lFW0
I5Gvc/NIWrpT8gGNshhi+94bHLNE1yYGD+scKHSnasuXoafobll4WTmNimIsF4JXuLGTAF3qEhzd
Ll5BiCAHkewa7Pv+zxIizdH7MEun2CUf0YEaEAI0tfzbBSc8FTbIRpmzDawa6x6H+ISJF8iCP+eW
ZN1qmLz7U9dGVJdN6VV/Dl3atqta5XcA0qUVeyeN+Kz5ZHFYwX8O8f0Sx1na/z/230LatwX2B5R5
vG4V2D+Eq0gCrX6xJwPyyQuVMtTV/Pkm+vTsPjbajMcbmt0BtIjZIg8rzchRPyj6QdKN9bqh4BEn
jHMcT26BHrx123GlEDgRjfrGY/gja9ieg1D/kBfuxnzm/k6eq/7EZIp9TAaiZggDfX3mvGhlE80r
py7vUdl7BKL1yKrspxuafpKa9fzk1P5YCz2YN9BwKs7SJbGcuQF2g4WPojNWttwE54PLXNDldr0d
ryJhC7CZM6KgqxV6BQZojV7RtmDh8EfXr1MG4z2glIXuppp7a3yN3C/qEQCY0qtnZAF4ups65Up1
wOpIkieiGiNYimqWQ1t/fRiFBf2jjQhFPOGhNWn1qXhxv/AAt/rJKmn0FVQchaxbxCE7DqLmZlte
AdgA6XnFh+y7jpqnfjhKXVaWfyQbbSjOuP5+4w3dLq29srEgQS79C7z3XaNgrqtUAKJ5SEM2EHaP
bsHX/QApXYfbGRlqLU+2W5p1K7L/LZdfHQO/DUv1CEWAEWtBG/eRqQUvNvREsn0uByI5TmbKUcrq
CVAVb9RW3CezzFRh+6lF3S4av5Wt4tEAkIL3HXS80GRUgm6NvA8s/8U44N4JrB730zQpgbJR7p7U
w+Cj0qHQic/jMQAQZFd3ab8qA/ljKsY/grF4ayLQGzc8eBjp2xIptWsJHxbsQPchSRvxmOQvE1TY
7gSoJa8LodZpZ42aFdfziTv+Oo15Uysy9j6JpMuZoGk6DPEkbhR8Vsvt7JtSVaW87i50UbukrVDf
njmdflcsHXR6ZSoh0KtHbpWPAbbEFgYLZrD12mqMW/QK4ZadmAXL73JcGFfUfTSvjVeqQm9uifN+
/fyF8zciQuHJdoLx9AnW24igsbdiA91R3/I1zNX+IslDeKgNPdNr24AARryEpPVFfhW534xYVQ+1
/gG08Hs2IHWvzpPYP9rammIFdI11XzZFdjdJ3w4zYhX642bZWwxIsgXJFX5TZdVqQ4l/ur1UDS+N
HMhmY2FvXrCGo5tWbWg2VXz4nO3r3cMQpwbmJh6ZALfKmm/7/8C9cHmPBfLSrsQm/po5DMM+enA9
tzTj6ICamCBzJ/n++i91P9GyuoMNvxpxkiZz6k9e+WmdSKF1O/MN5Io79V0vPX0jbj+AX0UFG64b
Ijdbxj5plAp8BpxT/fRuIJtkyE7OX5VA0ymE9T2LZpDXVgd2VAxyg4gRE3qteZmjZAvb3ltE1CKC
FosMedDR9+tfGoOQwMp9jD7USQQ85x3mkANgggaDpbYRPpgyw0c/xE9tGhT81Syga4f30IGVo2k/
6JWTQy/OEIPhM3wQ5+EO8ED5EtsoX2AU9v9yM6h5TwMbjLA1rMU7xwoEtphAgCMmyGyil4TtkbH8
sFLnlHt7yzWUyqEHgAVEwkqp4vgzXpUxj7dPQFyAcDqNKwE1Inde4vJyc+MG5fv6Tmi67CqNhI1B
MLRarYXpTRNAZTxS9ZmiWteqT46EzLpBObreIusGGSp+90DdZ7FXSJBtl4YITQcCgu9DUVWM5slM
XgZ5bSqyJzRu8web5PmyNmwYsjSdQG+VMIspIVjSIfvGAyBhd2gwuRNH41Dc3/ctMwaOhiJzDF4O
eDtxW/CWVJs2n1mSOX+VesOfIDzT3bJOPISXQm4AtLjUKIQ1Y0ldXdRy9xbGNBd60celFWPc7aQz
7LdXlsHb0dOOdHv95QaY2u7M4aphmnwCMDVgCzGX2aPMcN0iM32TR+d5mSxw8QaBN3q0HOuPhNH/
y8+jJDasNrfx+/ok2RF2crqa9AR+5T/iMCvWU5hjOB6adi0wr75MIV/6sr1SqOwpHbX4r+2w2qOc
OfNCRphuHXqyu30we5KzHtuiXiTnpcdOAfsNVrWkjFaymgZQTtplCYy4WzxCWURh9CUhUGOFSfdo
Q8lmk7utsIYLwaj/ayINX+rOs8RYeTxQnL/J4oip9eqwX3xCQI5382Egs/jnKQ76AKip8NpXGR+O
/yh3u1D3din1CS7S52vWSOMa2eljoWBxGl0Re6G3vnK/imtdTUpTnWqca82n0cu++8pwbkTKvh5n
avtqVI81CFR4Qsvj0fbWYtPAue93VpRyYXe+JkVrBxZYTZCKEqny95XqZ3jmBFF7DJEUFiIOcYnU
gtv/gc/K9JkANULXNZm3/h0LgM7HSXJTdZHhyM+SgAPsxwTtAIlZee7LrBoVHaxgDIuYrgBxfxU5
aNM/1j5vb9yn/8DtxZd9GPIi1illAW4d4fJqokQsR6Ji/qrpuIquY/KCdZLq0y6CMjqb59g8xoFc
7rBjUgKU16WwsYV6KrZMaqTWEuFrJAkB/7LiCB0mTXlX7bapWHWgrltiqgB1NSn8SPwj1xrSxhta
2BbbLFQlVD4bRd9CDdPpAPf4W0LwVvc9JyTomoif0qAUL+wgy8GyEVUH9w2AU54DWPdzErY5BBgd
9dbPd/NV+oYARHzVLIwdFdaInfGRxXzw3hrUbiM0HRZTDq10LQPtUeGzuye/OHgEO9W22waRj1Iy
FWBlYVrucCL+y3cyqDSaIYKCIuMfN8vnQaR1AdJ1XglCuy9WIaTeHSoVWgx3bCj0Ofsp/Fmcm68H
s1FcYGXmi0ouLUzp0YQCrVFoNx6sv1k2n0wPW/Utw/R+OQMRJvMGelVL2zBKNH9EplTkCsx2tdZE
FVgldHSgnUCkyigsqP7gm4erE4mtmE+1niEm9DyXBMUXsAnvGaUjHhwDP783hN6yuUjjB6cSFDi/
9RIHsayBPqhaVRoIMXmAgUmMF78SUr+57Yqve6iS3wB8Pk4aGZ+eg2XzXYBu82tfhTnqppUKVhhq
Fbex6VOpqPPSx6M1gFJ8w/Hxd9cjY+pRCKCUQwPxtnf4iIzYYbAnjSWeTU9h9PNIiiAV0h/McaeO
CYd4b8BxRwHq79RKN8Me0qRWQ5wR73jQgTUjFlZiOwiKliAOxz4W+EzGCZLGe2Zn84NjU1t/8KXa
SHHpk3+ZiXnv3TFkhak0ODFGcsAEnDIpjyrKs1MYE1r5xdSJ9Xr5KOsC8G0xQ8U2bdaOSgwsqebJ
HC2JZZEicMreUo3U+op3bQSHb6VtIMBfICMl3Ovz2TBmpxlYkUUjqEe1x85L7NUCtf6Fu077ewpf
G4NvGY2ZMaRJsZcDoEjYFRjSMV8yuhLZSoVNC/rvrene4xlAYYB+ad1vqn4602SKUJ0/iqTZJ3cX
l7V3vvYCP8bFke5C95QmzzSTit8l9x6Y0HeQehurIgU26ukSvRpd6ISr1E3uw44h+JUqzx0w3yO/
gv1nGyN888XQiXgtiFnHZ13dhmyBov2yir30HuICL22kYSn3dUWXLWD4/8JrLhgJ/SWN/EYvwPhB
qrhiuMORO2M5uXRGh1lohoACBStsA4J3WDmsaeuTqQlob2YAqafuAURGUqgN17xk5Xk05ra9cT4+
9m1hfztOM7AtycZLfkDHIK2jb4zIsCeVK1H5xdkqPffZgXCxhTtnS79E/D6mpXtfdUT1pjKxbUdC
1/WsjEvRe8xnl8KkjViNS1+Bcf7JgZyMW3d7fp7qzLIGPzXTJ92cbXhOrkHsqHRuPTxCJr8yBgB7
WoGc3pjrBp6CgA+U0t8OmU4iXOghBAalXXxODyVVr6E7WOnGxle4nwYImVeIJPAkFY5QSbI7EePP
XRXJkSfQGDE2q8thioLDULtst3suLHLyh5sWWY/3kDKw8WaagXOgzYueIgXmGhsHY/RM0XtWJGdd
3NyM/XlcAqzp571HNoASe4CB7j0JDfrHz1Vnk406uC3FWK2x98RgSCCLwCeWIkOcq17F6Ty94HFf
TWiv+sKAV4FNCHWL0C0QeU5XR9FN/BwjHvYhyUvnyRbd193gm1FAXt6ZcNPghKVpfTUQbmB9d4EC
U2AEDoSefcslEGvbck71/E1KTq3gb3IOLeJdn0STFbS/Ik8pckTp1fshlznchBpuqJkZPe3MABt7
xKtPdA706kHaFazqAa7g7LYYcN1n9XUQX/Jq1UhS0VuFWIivoRoHobtT6JPqLfKWvde+UFbFIUKl
7BwAlbJIFJLXQK7dBnDZkMoKLpHnJOL/NgdHIiY7zTKxl3b8yolxS70fSNERFrnnrE/jAoC6w1Db
16p/gg3334gPMQhB4p5kUXjr6SRQAXlZHtFkf3McwiU3TX5eaGODSTBefTogyGpHA4wuZ21+APou
WsjaC0ka1UIGurpGNcBOqkugO3n1AsJeKaKrQq5Y7MyXSzrAbudKaOMcGdaFI6qbQ3cni8n+usH3
WK8G36vorOJJvZXxoXtxkC5uDMecLoSxkFvqurJlci65HMpOlpoBC+lOQodu4gHytozgEiSwkXJ0
un2sHw2j+CEB5ug/AkBLtZGlvHx3I+7I05YhsDcT9wckEyGkeEqoayZbSyUT/mWVvgeUNvju9r+i
mNddK/yK1RiFAhKu3B+mJt50HZpAKzjsVRkK0RhBsr910vs3gzYlwy9qb1HWQEO3LvDLtCOZUpw0
z4Onmw6UVjUR6wHfl0taDfnj6E9DOAc5CqF4kjWbgnCYCdMs9r4lkFelf7Afm/Nu/DEGG84cUN79
ZOJ1jawERHCBoMHDsJGnszvm39LZLoy0rqaCMQK7kpA5nWe2CIj1HODYWPwjJNsxmij7PA09mYhM
PtBLOKVx/wY3icJKhyc6NpVYXK0oT5fruZaorjhXgkb8n7g/9FBcu2cI3+HQWjK+8GhWdbQGuIWI
wLTW/XdqcAV0asQZl+SJDXUyeDBmk1Vo7d17M6LGqreBNMLQy3mexm7l8fLZ8Tt2wtY0GHFhEc0J
UdQ8dnzNA8pshdMoc86JEOrc0B2L0YxIoq1JwY/oCOBRpEGoFoJUyyrc1dSsBT12UHAmTnp7Gkvs
FMnrTZTLi+/KpRYbPBZ9SsMM5dB0PNSF/I4s0IH+XvihsQGE6jphkX6MrNKseg3u98nGgicJejB8
Rg1LwhD2etGHXZe6jnOAb4UxU6egNldRSIsYy+ebHliKda44aiq0P2ngI7Yb8k1TzAZGJuKVntBn
SFaIwF3UVmyZ/ozqgAfxPEoZmejK/7+YP1urjBmIKMpqnc+5xJvK89jZtmB9ACSX1WcRS+4CDlyP
KZhmF74UvqLhVpnSjBknxozE4IhTqnorm4J93DdOm3sjctL33thONKjI9i7fVejnrV6Lb11foT8w
vKJJiIi28PtYpTnTdOd+dLQ7QtYd1YIxH43FFW8QW3+fhRmKtFnLTkWDgFdO89Nk8P+JAkyHhH7A
jyOuQssaDvMztKy0a0dcGkmRuNnlEMQlCZEsFisGq3uwkCvvr6fa/xyXvTTWPRN72NN8yMlSMdMz
LNBG3ROYyL4XGQbFV8mu0Vo+wP8U2ZNFb4EkcvD8fMbMMh/puLggbph0JuXzustGYD05CodF2PmG
htx3nNUKjWlkmOEvIxi/fNUBhJtime8bT2NmtQ9AcfXMs/94RTxSTS4B0JeghyhonLWsMsukjBEA
hKfYZcbg8OAshTMOalSBGhtvREzHdLkPWb4NOP2EiRVYkZfxX99ckv4jwIpU2xM7SNDRENimGggU
JdX/Nk6z3flNOSZ7DU5Stjc5LMrT76IU+2jhTD91jS7X41vyuOSqc5mFYwoc5Z9nc61IEoq35JnG
OwEXJGtF3XmFE5vRSPueUO+gkql5dS+P+g6KloRFh2DdnH8GpZRxmC137RKtyl9c1tIW+K3+108d
8wDXF+EZoH/V42za9s7e71nbwGPeabKcQpZzO8DSwwllrIBSVwmbBul9LNcAcYStAeBwO5be5Pfy
2hqUEfWx+xCEuRrHHWoN/gfLJ5voVrsZ6hVqfmR4Sn0No9Mxg8QZ7bU5KxtxoZS6VZ124KUk/Ypc
kr7pg8etDBa6uB2vslbU0xRw8vjzQFOOIZoF8lpRykVRixcRQuTPRyuKYfFOI8zl8lU1N9zTvbiU
Uix05BaIjCcxOZPZgh+PD3XXW4LbNiD+WreEH+TckbFJhm2XjoF1oX89jFtSo24jq24ywTyvMSal
X4H4q0sNzrDFwzX+Up1ReCbxj9pq/hfeVBuacx7vhYWfGDqjgI0ZX7avvN0XkmVE4im0ENJTYCB9
p82MWg2AxB4bUWtUwsgVMAW+TAU+/OtavYgCEGjlfa2YB/6o3j8GQyF3l8Qg7h4vWajxy9Drtbuz
V8oPOmZYcy+wvNdWgLj1lX0YPklxMEYh2eqH92VxwX7KEDrhl35pzbVbaraYPEDyzv0IY3ql24hG
6ANu0vG0qAht+B9fIkzpT3O1lxosetsxRF0KD8mXskH5tvPXCXdEhJdpEv4ac2knseeeBfNiwMXD
/IFuoO4SpveAY60Tykj4hvh8uwaucZ2fs4BzfTWG75TvBhdzqgRUVbr+yTYosnaMOBBgoZAjPsrl
Tm+PSybKXgg9ABMfDPeAPyDpUYMIcJ61AuRVzSpzfvxpIZJpn075ZdtU+MaiPPfxli0kAFdlnLqM
CMNYEX9xSvXZHnq3vdUV7YZBmdm9SHyE8/8EbHlq02lkW92y8L7IpY1nnE3ttkKk70w1u0ckQMU7
TufJIJA/QGmHI9ia0tNFdkA8u8mz4sFcsTMMDRMNWgjxonFURzzICImafqkV/fqC2M6FYhI0yahA
uccwfRepiKZQW5gKn0rd76f5dDyP+P+yKWSu5Pri0d01I654Db8+k0EGictgaK4IssLy81yrV8gm
WBC2IdQ/HYxzEDoC2qXhM8/KuB6kF6sRpJwFglp5q2BDGn/9hDN93s89dF1L/TWioqr17ZEi/jQJ
YJmBo/KW0LHP5qD+m+MadFf/QJXZuv0owwnuu9jPrqigPn8Leqm8E7EICs8fsNWoRlXRE7NhaKYT
AQPDm9CdO/7YcjpiYB35maKJDEg0yM6ej1YWWBi7KIs31yIq/DJeL4wF3nIJuSTx2OUo8DHKVt0+
oAJqjEtyQ+k3jLyNa9ugRvyBe6r+t6cSourF2KJSgd5FDuGELLpsANPOz47F7gv5JU/ehPkcTznC
JzxiA8G6hponGEJnSLmCwLD/CxrYGEY+79+iPktHMZL5/cPps6JFLvLifNW6vzhtIYOlyuOSc+BA
yr/wXXyw5zRCi4+bOvbx3gbX+KZg9ug44FPtv4nZpJHO2Knn0j5k4YdvjTIWXEf7B/AM2/UlyBxo
Qg5PvnZrnKcLlDwc2jatNu2Eta1xYx8y8GXCxCAUxnH0yCYHiZW9xPWp4uv4Jh7BzrCJf8vXwpLf
JkAW6ODeOUmCdK7bw/xt935GTtE23IgSyDCEQ46u7p/STtfctoKryCepWq2i2HA9x9qDrfrlXF26
nDt4ssoDtlv5v15CrshjKSpIhiBbG9w50JOOVa6ZEraDB5oMFasTZ7PyOMlSrNWOxJTXqqV64qfD
utPgrxpk1vrnQkKwH7POI9wQv4dR/vgx3zDLaHN/CGFNSnIbiUM04AH4vwtUKuLgG0x5hIZZR3Ew
Vse/lix8EkPyApZbXJ2zXjPTlomWmxxv4T/oDpLEorPttJsiK0Av99pCDmsB7d834+j7LDpbZZHd
+Zg20TnJ7hwP0aesBCmRR+ViY2U+1y5x2XWeXaR4TyPq9bT64vW+3UImwpvbdJVwEMPRSUPzQNlK
MRg2jiZL+Q/wr0D4ju1oihiB00a7iqHl+nvZaPaHDJuwCTg9jt5b7bv87w6X310+1oemTm6HnG4a
KW835iUp62n4hu/J1w6mNojaYC13dyVoqAf2szwe58IWPhYkLvpIy5z6lSupkvUmgO5FVdIYuOdx
/LU54VRyboNaEng67gOteZ/I1Zn3jZ292nwszrwqSklk3BroSsLtIx5gypR6y30JSxJYZAiJrEy+
7j8TsKrEfEpbAEeSpciyGO9d5xg9uumMj7Rcru/JNMUiXzFai1Vit2usMAH+WmzoPQw+NsUGu9o8
6VLbs/zfNLNSRd5ipKKV/SCL7T8UyKavgz2qKL1pNhxTkf/ZGdt2hc9iNMA83vsvEp0ERwfDbayF
tq8mBYSbk3I6wPRqsaOo2X/BmE005MX6KPEVlHuRMFIzAInSBx35dyuVmxVAocmydWU45OIkUYQl
klvdS7AuJOryYQrdRTMX60Zanll4NTbUn2kB/+FWkajVNvsTBYdjghT4aAQPAPck0Htttm6kCFVT
SFC8sbq+mL0f+Zb7Wv/A/ZIckycKNbtvwbwYLg0a5ybE6Gv+0zpAY0MahBGTUxKJzihX/VACdPZc
tTXV+knJy5sRb+7v6gfTfwPapk4yRBYOFyZDW52kPmXIZPgPF3QP9v9E6f7yBpRsToNTU3Im3+WM
pqUjaQHth3UIv4iEi1FzcoZgMwdxlaRWSmYmf7hujfxW/Al7wRiivm4P/x5Pm/exuK155XlDJCrJ
qfTAfXG4mak+alfxrMQhYDzrntuRpMwV5lo8Zq0UPySKl4SfUR6qxXqRhDzCt9FswmZij7YscqkW
1Zz5Vo66+mxqR5qCvVWgbXj2ULsSMjz97Re/kFqXXXLQjbHreq4/R9CCn3NaO+hDjxEjJIlkMZEO
jwfkd9Q7F3ZBVpYD1MXniF7o8MPvuUjAuh7H6DT4gnQjuALQWVKhyAef1s24Ld2wjoBnIySHu+QC
cvpTc4FcSzaDpKF/G8oUMuxR534IfCwj3HRx8RVTCj5h/lwtIbmvgLiRNKRGwD3QF1WSulYXJqgn
Vvwb3zBRdPV8YsF7OyFomlZW/POBQ0H1EJ70RcECbqe3+lb5oiRW6NSTbKpN3OXMKVsz3zFBgNyp
hzIvIZH5Tc+58QClBffnJe2lISuJFxgebWi1jkZ3AsaIDSQr2aqYqP/qGo5d+Eh0QUniQzK9O/fm
ngmh1/TTQRsic/9/4/gDM+YPd/5YbKZSC3ya0PW6xkeguGNBAtWE/3pMpjJZu7KiHQBPZkxGG85f
GCN9CeUWi9kxtWyCjqZ1EMHj4cVnkuqpWY6bwNTtzMd2QW8PkSQxQ+RIlqI3sHxeYYy+gWJwLpyz
F6WINNIdR7cPgHx8WFx+ZQsSbJl/JjFOfyD5Ezd67VqgAJhpMc43mrbS/W6FpAbtULjxV2GrytQ4
N3Wmv3mq2EVfUOsnwBu1W8UhE1o/coEgyKtMRdeKbCJTgtqinkh8Dqp86UWPuqmSLp9tbcdQ8Ul4
Wvjq9M4/qwpThLR1ic33sxev6Ypsh69+CjMB98CjsqMPgHK1vLscqAO3Fe9yf3byQWqB4tF2ky4y
tzzwl8JAwKi2pa5uwhXFbLShqjUPd+gui2vw7JGwdm0vDDJ9rARJjbwGr6M2M9ceSYMcgBMdgtet
X5U/8JKB79/OZk1FREGhw0O34iqPp4ZflbP9basiFb7wtdrkXGSIo+0hWyF6oPfRZ8oZmztvUyHl
zwqFaRqpM4CVjDZyHYbSWmR/D9ErQ20090fZ5JeE8+eOoktV2/yOXvdEd7uLiY3nuYyMrenj+V7y
xNHEYz4vl4x2AsV4JDBtObq45O+1xAXbVOqn2WH0unFE4BMSZWEfjnHqXIPguLD5m6iVJdSZtljh
6FfU+jiNobNxzTEY4QY0/7dRE5I6a+n8hjmmr8eUHgC9T1oMlbBZuKAtCx7DRM7a7j9c0h5qBl4V
hgbm4/hu2biG86n+fLOJlyW4TlyWIVoxGeLlFEHpbm0W42vkWJtCzExzJxzV27L1A4Bu+V8AYHz6
IDmoXWWN8njdrEqg/3QPj15jkOmV0OgSmtiYWPpqTrAYjuAbvjF9JeTVZxk6QwLz1Ns6SpQIe7J4
DzYcz8ZxRnA00DIv/Ni1c0qON39syqUPIIm6pDDJyhPV+ANo3jsaK30ThA3obxT0sTZSS9LJ7qFy
Fj00HV8K1FQxoZwBb9cK7MCBaiA9V/2g1kUuWzswP2puBbLtSKa6/M1kDCAEZ7HYQo3mNcufnmCi
E+dAsoFVnOx7OHGmGdvQLdK3Uoqg+AJOVDIUOINWonN02sKvwM6Ukc93L3DoIZl2UOuA1S63NvjP
37QzrS4xIeJPQxUkmmEwPdopVrOkYKOOrvyd/+tppsiQ2iN3/TCJU9/4ex2IgUUwGX5Dh7MuRS50
aEauhDKMPaFnO/EDqZtERClLv5K7lZjnDDlYc3q/WF+7P5XeYAmZsZ7cS5+q/enCzrLI/npREGXm
NgofUNvwTkXXLIFd918zuoaMdGlSZPYbg0kYr9fNJzwxOusRg9VnEcqCACUWg6MKKM9KL8qGTCIv
yaB08BGgEaHBXKzkH0Uipg7SMiddGrl7qyYhN2aj6PfrLOrJ2xFiFc4MqrMGPXEnVy7KtqHFqGVd
ecwSEQTfxhyonuniq/vOv6DX/zr8Y8X0yCiQEaTg2XgBAsaxQd0lyUh1eyE4QJcWIzjQ3nWkQFR8
jL4oSuXrLZtyGHNiGEkDaI5s7jyxbYORv2FUTrSoovKPnCK37NBHrPInjx4qx9tJ5Rz/kQrR0SrI
wBuiZguE22EacCMwfbOUJ7d6M8u6U1fbiRYQKSbB2afj/0Z/ZOZ8IZPq0tcuBaBuu6MPDj53GP+M
eCQenICE6nMuOoHn5u79X1rBhBitYmET5Cc5WBv21ZVhP28uy5pOEhsj9OeCjFawpw2yXfvytCya
7rj3EhoDSiZUsJToYqVHkuPiAm+AMkAdt9S85DSlvH/Bc+7FAoy9W6Z+VHRubUiIfDYwh+gfpfux
n+WG5Y//35WhlJmM1WHq3JP4k0zv3QJ/6iXVFzzV3uAqNWr6DYGlZK0M9o3ILzfixKwGz3tk9zkq
HkfjlUsLwOTwmgVX7VlfUZn9YaQwcmvs/dCt3r4X+13uSmBUrZvMBFIpgGjQ8eMBKbNHMT7Rc+c/
d/Pq4nv2cxpHQEVO/hqPMky5RW3B84oIevbHGML7Ov85FWpT3HRcZnbtuSTMGF6axmdtqcKThUVT
LIP2SYWLy+KESW0I3UJ+02ePe6bKi8nMFHJ3sa3BJodYy05OUEcknN+dPx/FCFnK9Zn28yFdpZxH
Sa3roJ6TCt45JMbldJO3rKyPALkly38YZcm8n5OtWXRC46A7b7sY014uxoQ8CzevLR/bgcopxYQI
XKcvqow4772Ti7DtSsrnmaWoz/ryw12fekZEdrk0qNtv3axBTmt/+L3bJ9J1hlQcQIYILp8RIEEZ
VO2g1fJStv4q6SpZrcyRyA4iuLybV9I1S61rAIekwDBELhSW/GLApxecnlPHZzP4f90cVtszYG2Z
4z4xIN93ecbHKjFnAdmKHLhWy3flMBch2USmZBcLDcELH8a0dvdGxPDLGFKy5eoPDFHAN+6xUXPW
v4bUvSTLKuQuquCDOzLSw0Ppo/+Ki86UPJp/IK7W256cZoCSI2TrfZucy7rhEqg2amgCFIJ5VGXw
7CScp6YA8pIW44/CIV27YuIu44OHCvudQ4Y3Z7M2mAQI4fpYz5M+/aC+HjEkuWH8k4JqXoYO4vu8
dOs4VSZonda+q5Rlvd/j4OZHC7DNL9JYrGzXAq3nYuODxshRPyK+ASHSxXyzF4jU4k+n3bDqgd3s
7gUmmZouYwmw4mV06LsyyUWA7or1zb9JJvDAW9o14VLvl8vYDyoQe5A5m/0kGHqT2WBZUlydwffe
DXTBxLaTUncjuXnVOat89WjSkdOlQGOWf8Rfc2TbiIqFxfF5Sp0uqp6AeazlNztNGtdbnz5yGZM7
pKWdygy1elAg2YdLlvp4OBr0pS1d0xsuUwQumWCALUDFJjOhIAxMdxQI53FxyBVxHMof4sYjYwW/
KIrp/mKowesNRjOqwt7ITXzyw/YDQWM4lk5jBVCeR4IdZsluIySOvWsElWuCbjHQz9TnyDQDmCyP
2fYnuk3hxKSSGQOEu41GL0SpyYW/gFyX7VTW//+Gc2XxfGejlkJ5Ub8Ax5ufFJleEQZzt1tx2hDp
bnFov5k9t/SPYueCPdAv7tt72YfD9k1iEQ1XHJQA7QLf3p+HQargtmdFSHYK0D7YJVDB8X/rC3+u
WSNqh7MvI0JjY59sI1BSDZk2ixJ/sq18KlGki+ZGxU/wjgX0kfzWRXfQcx6oXIfdRH+OOp27/qhW
1cfgbvh8gwCb1r+vFpLuIW2B+bA+oiyO/x1+asth1WmcvK1Rx5cUve+xIxQqUfnVeTDFAv/4/EJs
EhQ0anaEJA27z3MlWWsj2QwGe4kxkSSlCvrubYkyHGziF0yLt8pTqZ1gkmT3Lykizjb3DRI57dMi
bNQcDixuXoifBgq637pLVqFXfKa5N9HjRRiEMeRLFy+NlGM1HwZorMN0V/rlHOCZBK19iCekMo7V
S/Bxd4ZYdrw2AdJtGpnhIjcEKt8yR8TXh3GAzZxfdjAr8iRy+wh/ElcLJ76G6SBbr2saZdRsPmPu
3nn7+a2pb9leIto7B3O0FPCVoPLDZA5iBxgBxOshIh4NInaJj481x7/VfhhHmYokZ2X2J/+DzlqA
MvvxhTJHv8NH9e7ur5fLG6GkkMCAeBhxfBzfJR+04leoZmmPugWe7/KRIUMGGVJtKDDbBnVBMGz4
nTLDti3mQRla+x9Xiv05rksH1/xNLw587JJsVRU1iH9R5QdCSd9wLhGGDnIOTOCVpuYg8syKWfOj
H0BT/jqsD3HskPXT8k/VW+RbQYnTGGt5/G4+IrUhFEAeqsg/FCwDhPxeYVttww/C9Pg5ucWg69gs
0PpPbMbRRmeHTNZr+CpeD40emiGX2BOX4iCmt+6m1WxSD0m9lXYBcoE9Ql5ek2Nh1+hUnxfi46eU
XuL5I253H6dAyWDAmVVUNkcbgSfBDkk8VoYHdE27570sqIT5lUR52pjUKuP04a8FtSvV56mwm0/y
nfcuSlmUWwUIj1es/w6atAD/oyJd1IqhxZGKFpLMRAhWD0i4YqqYn7y0tacbm8O3xciKkJ2z5yus
Ccru5BIuOYR6U27/MCd+8bvBOgXT6+FimYjRDLNcSK1tnC2q9SjlW5nlIaKKyIrrGcqskQ9G7Y3H
WofgLhUpvus0z1UxNcgyb7l73CCYa9ATeAZFedIhaBgX1Vuaiav6Bu3SuAGrR3Q8+CMDOjT4Mm0e
+076+FwDrnAAWwATwIQqcH5l6V8zYMynB8zzTLpgEIBSiTK3EmDPizbtfdiVQq/2I9eoXmZ2l6BU
czq30aVct5gLgNWWnqd1WnvF1PKx7b2+fKgKIjDKz0YaeHSV7mSYckg627jGIWEHy2OTHabPQBrj
qYSG9PB/sqW4pfJhHo51KYokyL+y3p+mMJSzNAGwBpxBwB5w/42VJRJ8Agz4mBCfQoVXdY4ySgCQ
HZbHkSNwf49VRR0ZDKA+8qG+oqVajb3geXpWdj9de432IwXhnMHTktFRdmzwE+vWsbcOaISDVSu+
h7VKuUzUF/lXharjQ4YJ6+t3QRVR5lNetz61GyW6Zq13Tbh6bFUuCp6xRbAsu3X7db4oWAKQGtBT
bzZfIruOxu6edRZIdmyNifS39Uo0vkIpqxISWi2CGBksY16HL0u/aecZoQhzdfRXwGAjNHkBWKPF
OsB2djhPlpJi0USDlprLbAmUg9OrvM7XTVa+Sw5uu3LC0dsHjHEhjCj9SEzaIwlVuwsqQc/Vrbnm
aqb600Ytq9CjzSLbmoOrXNQ05DyBT9w5q3Pek0X8iibsTOdm1py6vLaBL88flZG46NJbD4dkjHLM
uYh/ZhuGiNjb6JVuE4tVpPAl3COIiaIxSw2ZMNlSkPI7fuAeaMmKEsBYfywIRzn6GWLVqcshIPv7
kn9wXgCpa6fq11/H8daEqIhGIfRzSzkzGudxRMGt/Mksn0foZXGk9OAfBgO1nOsMswH3pCuSV/+0
l9PFzkBxsA2A0UCqXydrcvM6dxs6kA1ZDhbQ3Hm1up9PiBBCiJbUKETX3xKEtnh5MJP+xwWHcL2x
v8bm58BCrALLuKVKU+n+gbuQ9hGvMSfOQ5LNyPSPAlnErWE7t8//ulvD3hpn4k5kgJRTL8Wk0vq5
Lgyx07xXGMEtkarUkbgLkStTLXXrjE+2YRluPWf/kIkO0iFj8S+DZgWcNHpXV6OxE2p6GXh7YNm8
z9X2uwwjSWkJZbJwfoENvkJvfXnM8w0OtvFAZSxUMAna17AsUrKsEjyFal2ZHTvulRh3AbVq0YSf
8GjNhonw/dU+bIAuk4bCRc8TIsELsub826NXijRrMNb1sr5wpV07MHlHzS4dKFHvL+46dqAW3L/C
brODg7r+YCT3xzebSt8lQJM4WrJOnSwkMvk39dGS2rYzR/jgkjPMPByhnu16NmL6E7gf1PbEsr2A
g4z9pRflwXYpXOl/OvjXcIMrv9fC+D6c8Zb7xZfT+rm0s3swb5V08mhlrK0aKuii5jq6iMv4fcc1
TzP3Z939Xh2SujCZSckgdmjwjUt/R5JQbnAFZ1vumyH6ZhhjvS+Z45fS9Cy6iunSNRrDCO8GXagY
S5Z38EkUl24y36obQoQ1ENkiYP5HvfP4l4YroLkNnjj2GMYFChH8aWYlow3M/MB9MfMgwX25yJPk
2OUyDc2mLLh2v4IQIwtBSZp4YmB7NNRbld2Med3Y95Qy/6NmRuCn6h55lPy/EQNrRfeN1QFrufpX
di0/DG1PdFpDmYrqZtHyHFL3CDKEeFPk0RCWxoZSDoJO1mh7DxLGam48MO2tP8olI0DVwP5Bt387
+nX6gH/a/AjQ7KCXKyQHtJgQhBdz3F+OAAAvLBaZmx5HRCz1pmN0C/F2IRua7E3VqNP9h0UXVZNE
th8fq3znD1/iUbB9+mFJwnJzY3dK1JZPn8+SZWcMEoIUcgmI/2C6yYbU9LiHQoC5ThBpyMBVtvqd
idEhB5rLUQ3Us4CuneI9RoGWf2NfOQb5qXYW8FJ+jTCjpws5VBy3fXnX7Z/YwNYNjPiadd2R8Fvs
mkt/5Pef3arWJHO7c9I3u2+BzAs2KfyeZLEC8foznMovOxFuE7asUeiFkL7YRHo7VuFRPTar+RtW
RYMsnXTBeQYLDInFmwQIcuyFSOIksB0m2KMDyKNlvE+8GlSCESlOnv/KknzAK4GEuqP6BfPNBVNb
TOBFi6cJGCPWKCdtztbw2T3Hl8nPj2KGylLxwDXLkMEFQlN3l4rI0+XBilCiIXWr/iqmELjEuSD8
FN2UNenuVLufX2YknJ3hAI3kYuRlgSBpyp0OkyRNr9sQJrTJQ+Y2kJgKHn1xjc8DY7lbYT/V9cZ4
CMr8OCp1WifSHrEgqmI8m37MdihEXy1m01i52hYLYCORdjkc3gHLeZIncA9j1VUknV6zFB0q3bQE
aeJhKSDYhkklstVGDINyBy1wnZOr21JWtnr4ncnAbGz1pknRRioxFVNT8u32AMNOUR3R8eU3rHJW
slWBjTcLmpACBVwbKZXiKhBYcmqD5wBo2jUOr/DPY1Jq5F2F4yY2E8XXIfDQLQLwEaLz0LiuNbco
lP2OK/xKsGGFMdXvK6AIWNGAo9GJtLyup4HyxYDyVJTymSRnQ974d9ROddfDbLgR+WxpUxdmHV12
s4hfEbT9F9zPdnJRfxzkHuRwWtIw0miMJKkskMMN9Ab0knUxr+FY/gyH7gjaC9nSpffNntRPHYCC
jbqHs/207KPx/Ix/VjAk6U2rrn/R3gB9fX9GMkADLyfZ/V/9yBiahDcf1QoN9orM8Nu+RGvah1iz
/nVWhTwwUpGoAT3u7D+nwyTWa/WACgACqP4gWM1bFeJEpDFw522+1K+LUQxykb7jyBIYXai0WwCP
uSNiPvKVbH8uK3qPbRMSIYws4TUCJFv+H48ozZkCcfayqt/znxZTp5NSaz5WAABHhgnhdmFftQul
kvk5H/NS4QPTVdGvZ3BgA9FwY6oSazuqdB1EpEzkMKEaSHUGl5Xe6IEOLHypOfqe+i+4r72agHwY
098lxLkf7lSOn5ZbPQWnRzsJODcpYjg9AHfAOCCgrb5jrQVUtsEELWKZtBmznL6fplQLxC5jDJuV
j7mlHoKWYlQwMScnUaJRqUDuPE/SGaF+O0lDVwYJplrpj32o4OvAATDgQ0WoKynR9J6FAmHzM/Q0
tz3kHaxKKkmu0ztJziv2J5CbhwiM3lV/RWbOcuhr3LnKtBe0+XoMxdM7+UNmNdsgBRLrOtBrrgvj
HyYpo6aGywr1VDWn6fwQq8VDEatoz3Eggjk2wBwnlu1N7NRtJcELRxtIbk8HjlS1duVTe0NnzrVr
tE9r8m1admqkQby4MJfKpRfXiHZR1tvsUDapK1suKB3VpdgtDRdtZA7nhK5K34oGWpAGv+OqU5Vl
YBC8NtfHmpCCrmbysUuUTL0sIzu/2Eoyp0LopixdksMf0XIKtfJ+KMEkY+kkUQXfdQfcUwI20pFe
jkZjmqZfvTWdQpYmREbvqAbDXlE4qNJGpPuaLpFBkkRxkDTzN8d9ragqG1t9yk0SgJ2pmlC1DnP5
bvaqr9md8g2m9fpezLsD9/wTbAl0T+zd97H6oT4dZigO70nOA5g1g5kTUFMoe6Qy5ABioFHmkKg6
QqfeOWnrNDGIlEqVcst6zJcy5mbFkWHbU6NVZbcTukStEDQCPqTx31FF3S832x2KGdd1bEtaSUGa
VdW4OzUlIHMMQAUl+E24BLjm3VJWE7w96SeM05y8UJh5wd0JVotruxIxwnPNsCNKqZ+XZ3k32j9H
0bo8uNjKrZuJizCGU6290ZMAo/QmnSQTZTV8A+RWQbPh2wKiuuJdqSUZ9c3qBK4xcxfKvrdR2R+N
CZ+rwWU2bqlMw1J6xwkKUv2BEDUP3laFH13ZxedHMmS8cSnlZTgC0zRy+3KzOMvX84osOKiCeqA0
sgA7uizLDTP01GJ9YvJTsjJgl6g1kI+goeOERxpQOeFSThDrPvN3rD7c/sD0fAqT+lMRee3wpIaU
SggDBtgAZ2q5KtAwz07m0cMOCy4iAYI3kpg/fVd2iZNzXodW+r4HFPbcMIlVMEFNlgkbuai5RKRb
nKNPKz5u4kmE59dpiUha9FXEDZch8OXoYwl1Bftf8vvdOfePIl4drEOl7Rnwp7C2JZoRnhMGHpjA
uxjDIu7//8T2/PSLHYo+c1DycOXu2OuOdtPnr5V0PsQXwcLQf2Eb3iSJn1Xh2ClTn4ONWJemHf/C
Tv2NLa4lXq3dVUYHLNSg4SKyXrjDW5KMEN+MDpp1QXid2MY+xxiLrn4iC/CCQ9wC7RuhnemnRqAd
W3+auTykI+Vsj9McyrzjuKzWklckkr+T/lgeAvZlYBWfHjqShFnm6RwxkGqQl/Q4hDyvCPWQGGv1
T2YjvkGIls74X1W4i2b5dT1VYlL7GjHFh3p5nH+Jy6Nf2NhHxcQx9DejbRcGRQL8yAmZkY3g0PgL
hbJ2wbROPJH5/01CGPWUGXlU894NAA13JGKlgAPmaCUdA2awqb1ly6VdRTaOyV2A7AIOLR56zx3o
u8Pnk8eta0oft+hUrOPer7JFEG2oK4SFyu1Sd5KLmXnGFoMhDId4jmnteyuzKquuGgYnROFkqEVD
+XkK3h0JAqhHhzq7BHzu3D3QjuQE/76FU33fx9sfVCxFDqzmFVZ5/smDI0GaZ9QpJ4dUU8J6myxY
RjDT2M63dAhPuXb3Qvo/9FhXFzLgSieY6Es9b+csXXrzrx2vKASyqSRHgk8KEvMH1iyiKwxZzUc2
15FXRgKq0iv0LM79xuwe7GRkp+AeCOowQHvCxUCNJdSnlzI70BP+pwztAZSB0905om3XmiUOsK0x
NJAjTfUh3rnBngyx34t6PAS3q5A7cCsqh0HKzRrpsBuXq2fgS9aBvBrIVPdRHe31k4jprTpYWc0U
7aMhEG+8awRNrWkmzCilr/poD7WpS2Z6ivkvX432SF49kbfNbCDvm8L0yW+A7Bv8cWPVBr9p1CUU
lQO7Nt/pBngW1X78v9Pnp3hWwLgk6lR1FSkplDaOaMzQpQa0J558iq8ktMU9lXadTjbutI+Or826
DPzkv92Gxw5ZRmPhaIh5Sc6OqWH58PXhMCYBX9HXsDO4ijlGtALzloegXcKV22dTMCShkyeWRq0S
rexLmcuR038Kz9aXrSzDed55vT8m281rWkOc1KhhuAkNI/sEc2P86dbkvf2gslT3BnahtnwvYdLK
+L2Be+3nV1USjcf8dLs2UVdW14zVj9Ut6TIgkVcBjiVZYaE7cYf5v6o8nx26utC93p39QpYXz0+x
K6bUVJyQwYhXZdgkBFb4O2QC95g5fhXEfFk72R+1aNCDeio8AzIBQOFXH3OaP8Y8UDsBq3N135xQ
KD5v8WEwYR5YwICBSLp79Cw1eUXsqom4LX96YqeqlmEv3d+rOf7+4gR4hmacvDdqmEXpZGDcDc+J
PYdmqn20A+y1xPatDUta8KYIHXFbWW0TffBKyI4+bVgZdE44IQuzzu8OiXYkhKHnipqw9iVLWatS
3JNwjv30ORwighZ7Vthzsh621GuzhExf8RbARnDo4UGxVzR+cI/2hW3rM/42lM5q06vorp1oKMRB
Jl7w8YgLAhMLANLplfg0+PE4cjx93pVIAlERpsfhqxOSE/8dQTT7qsbHRZwF4blPSHpfB1MI7zPf
6XBUmTtKDoOmOfvk7joVGew9GCEx4vVoRFoDr/Po3kmB6fKlCtp2sVlqKyyvlQo7lW/Mld7FZmjB
hUSmSPEu+8jq0xe8ssggrEmXU53v3RoKZ87DgL2NsZPcs7xsfsV47kqmloSwaMsZdoYn5rVbKQov
NyTdVOrQG8h/xhTTazEd2H/Ix2KT8VqH80uCTYVCrsFZJWe8aP+6vDWMbRFonM2PglsQ4SX21HFH
9X4f/2J+U5wKebQaM//FMRwW0Q1vUKKLN42Es5+1Ot3T2kZTdZ3IOKgp72zGRsX6ApYJKf2lfMNB
/9tU9/y+3bZLXNqObuxm3HZ0UViSBTI4VeIWcfzGn1m/h0t7dKhrDSOP++daU7R69OI0DN7fZcOp
/DAO36OuP3FLMwSYVLOTNs5tnsCjRFpoPxj2Q57QhXHDpHFPJALm/1Aq2EBL6PJXzKvqDHEoxa9u
2yJiyYKJpf/HU34a84TADFRzMuXhe+/2sG56xVJefueoxCqAz5bhSoK8zCpEZ0ljhfPukeQaUkFg
pcKClUogK8QBiYDR33Ih4/juLQlwsLRFidbd928ibwoAz+j7XPyaX1brHVBcbNrrLJW9zQXohBqi
sVMZuwsU4DegyRS89rsJj/GUOg4lZLvUl7PRilAvxZiZZvSc2ERCdTy2JlDjzK4FYZKnAunbURMY
+v3Pm+m9y8MgrGhpSvxv2dZBkIAiKGSWApOmfJ4xuJVgQq0Ryhsw+aLobWvWHBrLd5S7jDZad1Nn
likufNm1hH+XZgrvDwSom4dpBHo0CLC7drOAPeROlHttgzG7Jr1FrtljeEpEuJ9KbkmKUL9NO5Lr
1hKGL9KrzJCtl2S4VJw3d9UIQ1yy88nYbg2VhCitQIZ+tqcFGYo+/ddcsYspkrFOyt5CqruL8vtT
1+tFkqmrm05kiqLMnB8Pmue8kVznSBVdWNHU3FKvK1Ie9PeKCWCvpCzpgkvj93oXPj7BeI3qQgXX
f3XWo3nnJgKjUZhTL6v76AbcIoGBIs0ug/iRyLIuuuT+qaDPfDVm6AJ9Ux1TueJS9WgntDWmrdE0
4rtemmUZqXw7AuadJlO5vuRVVbzCknri0KkKA/u/XgMUstEyP1LffvW8/jEvTfzP7wplw++d2dhC
EugrK/IxXSmDsIW5j/gTgvrMjkaAJuY4BOJv+Bq6xQmXQl2YpitwQi+n6IeC6j8O3KL1HI1bfuE5
PdD49DEMVr1UuhmUAzCT1pritCuq/Hrav4WS6jnMT1N86BLvP+RdaQzAehNoztJEu3XIjYgkp/D2
+OZ4al5htGIkL1SQRg7YtflYmQcTyBH/Pv+5TmZqliBpYWs52mL4jlUL3ArdIyt/jyAoGYIjesfl
fHuK2MoWKcdKylf43j9TCZ3J9XBiXB/7xj2Am7OoxHPxnKaVYMwHDxVTls8OojF++t4ayUyTB22c
8+d43TJhgQl1KcATeE9CgT/9kVlGOvQo7OtYxbyZP+VhiHjlB0c5+iXBxjPgaJJ/yy1QqNo2NTHU
FN6UeTYrM82ua/MJDYvzJTDfUbf/UTTXibcGdYeqlLrsRQq6dQdNH4j9deffPMgL/4lXoOiIOFJ3
SK33HPf3VBJCECyllPzuR/LLF/HKZYzlD5VKh0o/LWgixpJ6KdrJ/ocdNWv1XraYXnstfoQChXYn
KmQk03Ff5jc9hgNAXIxt24bBKAQUVNh4/TcLlhZIpk6e3c10kivDbvmomSlSZokdEoRJUcgb08P6
sVZw2NSn2PkKJ8THct7UYxjRZATbI1tet7+6H2mAWvPB/FgmyHfH7PRxKRFC/ISlPrndOkdraNnq
8jLoKVCEq6W6fTF8WSt0HByaaRX629jD3boi0J3XgG39nRiOY6SSUHadbF4B30mqgfes9A61GIEG
vaNbAwXJ7JV4k5YqOMPw4cSV2Gd0c/cua6v9nSTtu6qwe+lqohbn/Vk3eYQMpwPDjWOKEn/1BAng
JpJUAfEZwUwGGmwO3kbnZLYESZh0TSo+VHTv6r0nAvnO6/QXx9SfF+s/RWVq6xViOj6ZWqSquk1s
mGlfZKRB9s8V1E0jD5FlJISTvBl9GDQB8bYV3T8YBlOlJvOLEZWrAUOqvO2pZWRb8mB65kPxcfgJ
2La78BHdua6NIbr0WMzrBn+ICgvr/vD/2AAnmCdeJPMACXu7kuSImND6gvkLrpa8HczzKS9vlPbU
ruESNHkgR/gLINdULLB5asJ4aRrfBb5EYSQKWi/GHKB+ijqwTfdNgOLtNmanmZ4ERJXHJZ3xu0jx
C3ZzzDf8F4+QQDPlwuI4qG6L+pNM+LwmaSfM92CfmvvWAbFBaIiuPcfKEla7SwCZOKy85BA+JD8G
DOcOj2CYEMoQHXy5kMQmfLNQ79javpDSWQmXCAUE5eo5bADJPD4m8eCnER3psfqDKRoQvb1Q1bq1
QAh9mbyMkJ5ZWkEzfZBX2JmOFM9CPcnKT0AJ7PdHvnggSNbIwnPXC++au0x1tyF3dKSAkEe4Sme6
WFLye6h6iWUSKoQLrzGh9vagcFB+OfexuSarjD0OMIDA4QLtTqLqrw8BrYkkaGiq4lDhh4WXhidm
9C08b0PuosqAl3Op4yLd3q6T1ATCpQu5Q5J2pE6lxqaWw1cjo0Q5lOkOWWknAHNwT28f+2EEAfmm
geZ+jQWrcam/JMA4KjGOZzKyk4aPsqqOAUHHv6Ky+VWWCJgaBwQw47yl6prEJtepQoMCxyop7Q/l
WWSCsSO94qjwAWCL7pNW11GCCJoFl4ebkjevo2wy9Rwfhv4mKJohcOsncC57YhMvggLVzbJspKTD
mMk0puJt6QfW/UTuOS7i3Tk/IUiK3PA2L3KJ/94r4DmhoHX1UoR4JtYLFk9aKLobkPj8YxziNELT
R7nW22B1IPr2NGc3LDHLkmLUd7JBnxMduo2OOHo9SrwoR6k3C434y5MosVNHjWJF4Xhb1VzJlsnw
lpPGwEXMd+vS6kIoTPP4iRnzud9VUka+PltWjz0XMwPELoekN0duGnuetaurU8Z2Nd9KVN2HhkhT
Zozuo4w8KRK+vsbmSMXuMYfdXoi92jDj10SbmYg9PD78DYdKecJCg14M41VI3wwl83PWEZdXw623
7NZYGqgvo6B0lWdnhVQXYN4YB+KyJJXlT0H0ayjk8UM7oSnknIZ5Pmq7s0EXZ1Al80yfUi6KQQxZ
h7s8CoJHpod/RHPZ/X9lGvfFUWKTa1NX4Yg2npg4rwnGPidzxNaXkpf6x1VHQJUNdtXhYF/FVQGK
x2tCcHuAHmDz0YAqqmSmXHw06u9br73hMzXLHYVH8BMRXdNbWX7erV8OqdoPLwE5lnNRVE7MJRRa
a0I4vTq8COY6YCpGMCEB5QsqjpOZDIiqCWPACcMXQtmw+lHQWcIh13VEMuB4+jXrMiK/klHYg3fL
s4hf7nxG2HFyJgtI/jo1d1uE3QHAzOT6ASboYbYQRx66N0ilL0dgAs8Rv8JmVQyx9BsS0InXShn+
nCjkbpvWdbEUlhDuzqJzcF/Sj76uE/16fo3BbQL89qqJ85Ft4FptmryMwEGHchnRJp1NlAwPkJgk
xKvaSCf9H+Nya51b+3QHrdPmJsBOAV7VW3u7vuErk4qeEqmScFmYFAfcRB5TXtohT2P7hPLUsXWY
crdHFXB6ih//JZNR460rLlFK3nhi8584r4kxEMZev58biQWwq3tgWH/eNvVTksGgINqyZf3trufP
BsPXXCFr64JV/zLoRpOyXhkr74HOyFrARejYEl2ZvFnjHjyDY8s1mXUkV95x+DR6i9cBKpY2Q7SC
9xYHsNTmlDguW9+Tl0GeIzs8qpYmx2bB+of6EF2/Tt6uK2AVWjYcVa2EYJtlSRKyXLNCgpgm6QfZ
dVgG46dQD/k9dsYn/ZzFXVAt7jqYgdDXDXaXyytpHrK++uvA/LKz2zMQXv1AEGB9XVvb5Ivb2NB9
n1SX2hlBUUtIbSXJI+zJVwt98JmhN/uaAdEPhYXfLLlTjcwOx/k8E+ewjZsYOMwklOFm+eF7ee0M
+3n6LObFhSZy2ERujTKYOX9Q0H7dNJ+CmKVmMiYnO4SoqOKRJXpLv09PgJkaztkzPhHmHfOxjBjS
2hFz5FK8MinoNdEysFpFOrtn0VofFTvxTtDnVUR4IktOUHCBzArGNf3BbQHwT/WXtbCE7D3E0ZFa
h/H0ZIFJ2W6X5dRzIw2iH2riDLJasFgNHzV150w98PzbZbjEp79HMUHJrGBKs2IVIDNSkyulFXw+
kPfQtNDo1L0GX1rfhNytDYPZMH78iA8ztSC5/uB8/tJAG8L0tUav7WjJS6dcMFzp2xPbdZ3Ah2/y
zR2GORIbKO2QdasJvbaDX7Q36hJIZ/ykSUaAGhlYGBH6rV6R46VtCPFS9tXLugGbgCcdzi7+V3Ic
I66mX8k40kocscVwms/uaaJZvh0HAmNao+0VR5YsYNL5kOJrjIOgUQWzylwFTaFmI1XIi9i7Sy8m
WK1ys/dEEDnFKCoVVrMUs/pYEWr7zg0OMEK0A/rnO8lYA16N7H3SEAPh6mLCeoAGzD4lb1i862Vg
IN9nRUthXNJ0jqlVBl9zUI8zP3ol8c+sD/CarXRmZ1mrvPfpGekdY340hCOfmrYVyRPnc0sSW4pI
PcezNCA0V+q0n3PU+JeplHJUfP9UDKaOHfpb3Yu6zP3rgwAVr0VTIzikQjMh9aJkJKMzzXeqoIcs
D5/LSMqxHNiEZZrT/RXT85u/43oz4HnePIMlXXKoCUKBtlqzaU+SwVggT9r/kiNijtsfBASmFdoJ
LLSsZdQ3xJVbh5KT15v5/+8zrmbk11FnXwR7EnegvH6+DmZ1sit15QCC1Sv6N1j+iNbJ73Fssy7i
5A3dBGD9ImwfgYNwdiFIlR4hrIvMSVY3dtSBBoFSWG1LR0qpzWSNqWgn68PVnl3d6MnOcDxh0WS5
9BzDNHAfVSwhA8hJC7QJBPBqbzYq5BptoPez+0VLSE+Z40cJWJfSJBS4qThNmqS9MkcXiHpLoc5o
JzqhWyCoyUMZhMxfmHbU1+7qSNrEhn2DvqtCJ/ReWA0XsrW4Th2IUj2yPfaBsNf9kC9vJS7Xo7ev
7QfLS8YUFz7MDRM5VS/NrvDq1W7ZzthqIsXhpo2glGNG+cwBWAQFKO2lL/v7yXkxPCsr7n+GrZ+g
Rm3K5NETE7MnwQmHDyy+As3xT6ZWH6aClUt6t2TGJp6N2rX+Tba8orsOufOl8Y+suZzOa8MwsR2R
Hh011CKfSm2D68poMbBR8u01PhyyLeFwPWDCwG7XwO7RLL0/U2MBrVQzH1xSKNlQU/ulur3Hpu6/
vgtq7Od6Nf2/Q0v6b+i/PEdugfhxUuPdAm+fQ9+6A9Vm0SsJsNoZPNqt/Yz6qkgrDnnNpeCIHj8U
65WcQUP/SbegtiuZnancUAhxlth6cM/scJly3RzBR6UA5lMlMyyFFKLard5Df5nxgZgHra7Sprle
ldK5/5UgVotot+iKosyrui+sh3xO5RcO3LUxQpwewWIzYO7g96a+7ZsxqPNNzJMu15LDwVihtIjK
CLGohFOVC5GznIXtjX55+TSYApr4Rf5YdS29LhLSfFXjkpKgaJA/LqzKjFSYs7VyJFV+JmZ1a19b
24K2tNh20osQia06PrroYdDnEkLgyUVMPFES5shVwUk0OHeqMkuSqVIdzTvlPm40c0+gX3zF4Nkp
/wYd6xtC7krx+1k2FbkQQ1xWUUPxLurGyCoD9RsUFvHzDVi3BWmU9iKucDxKGcwN2Bc2GkSeTaRv
ldj7hIjC+cMIc0JFf08klgizHDpVwmPD7fxzNUs10sCdl75Y5udf2ueoy4tOtCX1pVG/kgr3T7ED
6zyy7xP4ExhYynxKjqkU19AdhotqZvnPC4Lo4crZQ8INUBCm87972uXNPrgHwLtDbNcocbIh5xul
vFecIWSORE2dWRjkKLvwJA7Re+VtdmUT0n1pCaPqKKc0R/hWdZE1EEojyMY0KTGaJ9bLfDxtB11B
3H3Hmwrct42ThUonGebwlu4FVkTzblMZq3L0+i1BJLzUjWdZz10BLohPKooocKdqoDauPNqpmbAE
88+HsZ6yGr7iP5v4vkdd2+SFeQD3o3/om0l0GhoVGRl0p9z+CgV1Xezd/mml7sW18we526D80brZ
s8BP9k/bWfsvSCJA2MESAF1syq85uFASAScLUVpkJYHtPSSwxPWBZZEJIljtQ2e9pTcQAEKUbga5
7FML59gezMt32MmhBcNwrW/Ri7t0eQ0uXu2qQarGTCIFCsaoW2ifMMVvFCMgGFxeDAd9bVMOTdPn
0KpiNm4q10lyABuiGJWIV80LOqtI9MG4js7Lu4JhNxiODHYlJT98ZAdNqryE2CrZ6YSdqIbHjPFg
PIUPobhKCY2YUqECgd5V4iEzXXrmwZTqD1fDsdQrTOsivWn5bs75NWE9TCVA/lKV9CPQWAFwkF67
Wt41kWIBToO7ZFyXMmb1+sH0HfOtLhw521X8X+gbMr8IGz2hpYpPu0qH5B8UUE/tUwT0vV6IzlHg
fV2PgmQ8XMcJF2wsjUf3FA0Uive484eZC18iaKWx0L9gaw2sKcP09Dj31r3DC8sgOlP5iAwOm3r0
yNFc7YV7m2i4Y/sXTGMQHAw5D3CqSo93xv0v1sA+4MK7bR1ugw6GaZF6M7lahcaNbkOfh8J/Xyod
1Wcs9qwq+jP3EFI80E8jkAE2l/ujYfm5PcazOL9ICy/dOn4kRT3ZF4dT3hSoxYbtaMVZnuSdfCpl
CvcX91hBPTOxG2VCXP3xjkPgbZip6qns1fLVI9tVjoINIaA8yDYeA68fTTHzmVct24RgLUZ4a2RW
//ap9wESKBkrFPV8Pf5gpk6zHwPyBb8P/+8BVT4GIzJGvlxfFyWtbzVigrrGEdUmGPhjsiNgwWBA
axYak+JOYCJvFeecfUN7hJPF9ff2mbSoo6csTqwaVaQIWXH9WzAgYe0+zB9PwJF3yaNA40lLaeuV
mevxxxk/FCGPro5g/uTAgMt+lHfoj6t20bZVNdnsd7A4usGAWsdDhi0xN0zHVLWy5LSej/BA0lJl
UiOvLNwgnQXKfJ3WNv5sxkmjcHCUp8V2dUtz4/ddsBE21mwnHI/FNvylihh4M2FdnSShNS+sasPD
rDIx6Edhr03QeCLSYJgQLIK5c4DDxF863G8S4W3rB/hhIicTcZc+29FWAzszuZF4NLGPjdnU1VqY
rLGz37+SktwgwzInxeorWE+E6DvIR/LT1/jicD0qLI6BQm7/XKq4uAqjkmLVHFZ3kPfqm8doGF5v
mtFwaJSXr8bhPs6J6a4A5og5D2v6IXmeG9UTVu+jUM1+jAJVB4AFaduu04qL41rn8u1IvZzrGrQq
y6AWmdbaJAcnydYqr4zLUOVeYsZ3iqs6UG2A4CamAYQsQwXU3dGYeTBy4cFV5+Q920DVS8iCtKJN
vaDaya7lmqjPQMNp0LKSw6V4H3n5BOJCNWwqffFIBTET3Alv/OaYgVjoUHPE7KX4Q0ELozQkD1+p
Kozt7ETPnCoG37zRL25Jsg8XaoVXH+DvMs7Wi5atUxdcfGsXOMszwlpHFtRRs96K//P4gSmWjrQ7
JSZewJv2i75Fwgth+U4nw5I3Pg2YXw+T6J9gmzNQTY9jFmwQjvZpqQ11YCmbPVzcrn6Wg8xc3YOr
DHa37DQRHaFB5b7qBTd6KxanN4y0YrX3lUK/4DIZXN3wOnkqwVtlHtjSIk6MykVJH1aynTBch/se
WQnoyPtP0ZFg84r90lIqdxjP/ZBEsiHl5SWpv+AGnbSAqwUD+lpWObT3jalWZfhQI//uVIQ2cP20
tpFq6EOEJraBNXicTIdlRkM0rdPIcuWulkql9Muw3r7JzNJtEgM32oAUmR1x/7ioExdGM+kqIeWA
Gyur8qqQ1PcaAMjq9aKvzEotk9FbDPjA/QsXaBZSByhOfZwW+DWHvcvTNTSyfemToC8lpsu+WBAS
/YPt7KKamfYPFfPKMB8IBhGdCnW6NNyTBbTp0y+IGHeMXUN6MLe/snOOrjyOg+jeZgfOh8bWIEsB
GNh2cQH54Rv8CgCqiovMYevpGg09JIpVjP4OmR406UDeOwjGisU1Z3o/UIFWtF0l4uehQ13Oi/Vt
+qRZ8Tzg6QZ5nbGW5uYzUB1VGJXxpBpSFgYkvKeoxlmPyl1KpG+XnENaXOfl5nR8kpqT9kU+LY3L
eGfPNmCv/ohE+rKQ7fYoa6SgzxOxLEiU7+isCfMCbsYYxcEiD1LwzPByBV++7xBEeXAfbG9OJT6L
hwSZYhT697Uwis2GPiOtCHD4LW2FoPepLDAf2bj0ftalBxrjKa+8U2O2oE2uzwCvX/A5mHuGS+A2
y0nxn3PRN4Se2Jrsf95X1OSE62n6rVK6ozL5O05vIiYe5jM6tfpFtAiXmpjLGEI5/8Pev0QLsCgu
lGq9W64tXQIBOnxencNf2uiWe62OGZw3wUyFIWWcQmOFREqlYHU5pyZw05xJpZwseCVLn4IF+frh
DqkEsXXmOE81acwUSu050u+NNiCi2F53dmhPYZgd+A0Is4InqqGxoRo+vEIEhzQj7XD7S4Foid36
ihsa3Asm1dMdtdOKpOycMXU0FVKpo6zWyXdQREUpdYtueblexjkdMi7lkvrk1V/ZmIU2kKUj50rx
T5cBs691Mju/UJ79sipXK3L67QMIE7K/X7iW50Rs0v8YRitumk4/LbJ+cXw1YESQXplHxw71KvjH
mexKK0pu3U1xPmGqvyCYL/enR1Pkx+xowwxfALTf6VPBAFA02vljGhBwWUJ1ZdVXia92rkHBTHla
itCupyZxnfY7qZRZkpfMomdITMwqChnoWLkGwawbrSgAfzVwXGuUEX4J0I5CvqS3QIP+D/6SVrxi
sAij0QJIOwloc6lmmjto/+o5G8r2zY7p9WpXlPC/tQftmGYKmXdUKn99vhyPJdm4XVCzQXRPMYgp
LHy53UpuxS/NCj/oyirtqORz0jkJ8Igg8dNT5v6yaVQD9tDQduUAdDgG4RtjFvYx61TcEyD+sCNv
mKTpUC38awtNgTmwwIIBpfk2etGpw2vmx8g3nR/+BjPlhPFF5IqWmIf76EQHmQbln8PsiFSZgPsg
GNbU+pZUD35nBRnJ3HivozjzpoBqPMQlAf45Yy8HaJYZwbd+HUMCeBpLv2Jazsooq9zt0tzWMUfK
bLMftdJUCeGU124eg1k5z2UXJK2nRa6N217FIB0RPSNOcAIJ9HmR7CtspoQVqKLa/KaB7SisNXOK
JeucGCopZuQpuEBPZGo94fnjnlxMd2QNpAr9Fjxqo/MZicPdACgFI9YujpqTK9jVllDhPNex4feM
R7hlJbiayFDKqHGsjMZgkV4pavO/fX50xR5d/ezTgYabDTPGfJx34JU6jp8Nk3itK+7fdyVhccsy
ulB4dBYK/aZoWYh1z5QAAD9XXz7uNSqSX/8heI35/F6s4si2val+XDfkgkXveElbtoo86wMdTZ67
MV6/+zXX4eYFZ+BIKcdQJhmcB3nqryYP9bK1DJaHLZUzKOiBwt7hvjpj+LitAx2bTJDDns868Akt
vRFOU8XHxhk9ZAZy40yT0PW8aXwasVdAn2P9CD+RZLh+MN5/g0ocSlTGpHNBLlrhEMCY9jGQ1N0U
W6aP1Ty+vmOYm3km0LXvS8W5ETkclHfbkDEKiZ/I53QTyvQVK0YIxmQ6bB2fmJ/iAR7SFVRya86L
1eXFTDpkA3XW8y7Ul7cZBMzBshMa2Qc7APAHB+uhRBznDr+LdHGOe5yWxm1gorrrbN/xKwLMBynC
qVGsmoJ0MKCGZujkLXFMiExSOST4YJpvu+BYvWTCFOcGzagZ5IBRK4hD80PD46zYbcYUcJIlLc5F
o5vQKhFMnEEromWDdrct8oINSHAeVK8CBt/vWfZ1y9nAnVjZD/W2dkGb7pw7MioikoZkiWXmy7Xz
MWI65Dsb7pEkPhcBIy10ur3zqqxV3oFJ2z6+Zqbe0cvku+aSITNo6yssb7xKA2jk4c36uEJaS46k
qoE+UJWgXlVSSVELoXWR0XIKzozvglKe9s/SNgHnWI0Fye3UUHsmzErJaL+2EFK0bxE8EDC3p/4W
Zdib2MuTSTf3gKLLBqMDLcQmThlATGJ05RYPuqV4Gx4voSc+DvnSwaPWxzSvYSOVm8jeE5qQjnNB
oWOy+EggjTIXf/il4aT3hWi/ZVJlO8SnYWWyGCVZQpUDy3ljjZQFOJVYQnTxPAAZWEWc84meO24h
FT4HykDzJMGeyuYCt7SRBtzHFvFl8xL5JTEkbxavisB3MTnk5gAPA6mVgbYBGCzUbt3sn9nspQpm
PrgNvm0zcDtMadBg182X0DcZILA/po8Bo42OLxqiTGr0m4WblJbTPkoVHQCVVAfoixQiD+ye6iBD
5G+4QejceO/GagPfr4QMc5PIqXlAHkW8K4yUp/epwCIH673asVdDh+amxJ17NPCBiEm19AVLs/B9
LETmxUxvLIrnKwg33U99aTkzlYe/obOx6zcr1iidCxuVrzBohsMIF+o2GM6SFZggF1CRfdYfAO6A
cXH6yV/NjzJmug+xA5Ji9FZXBXOjN3Kz8G5pBsGapeTfEum8/oFPYEmRNJOWcKi5TFXpPJvZojEp
qj+X35H/R/8ki3Hel7znBgP5o38rxLm0ChfJ73nQ0NaP2AcjOXDRSRpltVIk7VHSJXJY9/Mp8YjV
whd3/d3EqXW+yeyNXjTjgbNrYNtqEX/nWm/kqy6DiJLIiuMgmL7H1yhm/lHn9b9eEfwN8iK/JxU5
kuIymIQXRbds+v3aSgof7FddRckN3WztQfVomDx6oHdhHLrkhIMYhuu/a9xZ3CDu4xvJa19R9D/p
Gx6CNr7NGnVJGAMLF00q1B9tVb7eYrTygwBjFImxKGTvt7bXuz7pUJ1gsPOwIwpyvGIViodAW02T
d/OcuHK01miOodE0NQdxDGzR7anYX25yxEv+9Pl9FjKLiJ7R2VryDxT7n1VKhYBAnR4yXBIpO+X/
/ctQcPPuLnmaafYfGZzTscaYPJMJF5St0lEBneHG5mzcG06aCxBEoNBVzJgqShwqCS8ZHFTJMy2/
7iAigck7s5L2QOyX1quTJ7DsyQOHaLt2K3PZqNiE7AHyPgZO6nUkvURV543f/gjIOKIZA/QeWzsh
UTue50bRx+CjSyQZI8ENEEJdXnzryrYxnmsI/mOydz539SHf2xEi+QiBWDfdCw18VP4QGqMZav7H
dJEmBjAD5cBHgeTkrH0Mf5mVJi5EelzwfagtqYS4qkpCQk6lFj5n2dvR2mvobMeRtR/KsZ4T9v83
3gJ42GFP+5tKsyYbXQx6KHgaMXAcMMLwQ3qKUAT4fHasejyZOBL3HJUXl3D6RFlGKN3x3Lck3eOd
/FGIL3WUN3kQw4BAN7B/4OweL4MxBzeLUnfnDMYCUPwj1cz4opFEucDcO0A292nliORdF58j8YNM
IThuBVO2rCeK2cLBtPVtGVSlInWzjprtt5V+gvDPd9yv0eAwtnyPzrWdZe5VH3iR5GecMOABI4JH
/F3rfZfg8B9pthblEYP+0ja+k1FnrvWbZF9OAIfl9nk8A4yjjePyzdY5qL8JVjU3yu9u+Oi0D0ng
Vy6n/Dwgj+CYcr9fKLAbEy70FhQGr9kyDdeBCY+WYB15fbktKZwiY1cqZJqUbMs9VA67bKCDYNiR
/hhU9v6PG18jZYwM2sst9uzFzjUksUI9n8MFNYL86BjZrHgSrU5MT1U+YE1aUL8fTND2dPElVY/u
977zFWWNvwyZc4/VSl0J2G9Wl9Zr5yl5OCpgyZJ5RdPqm24aAUeKSlVyALy2k7V7PfxKhyVSmkMw
rrgGH2JNPsvCVLGGnEgt9OcC+liF7b67gQbRYAkLuZOzfrvvJvBBc0O2q1YxiTOCz2lFXB1V0tAd
VvRiF24tri8aiMfQwz4FbCn3CC2R8LD1IaDFKlnCb7YUMN4IeEDeW0kv5kRh3G7Al6LU7N7fiHiW
qyRSzfSqkf26xvp6G4mdx3LGCgMjg4vETR7ypEL80rkNxZFifV8WO/GrBuBLHZUGgw8fFGnnHZFN
9HeQmmGdtzKCq9ideKHllDuIGV94pr0zay9dq3CSP02eMo+eCLN0lxvfB0Shra6q6T29W1EA2GBa
IJp+5TiAf6zD/ydjITMwECWtZF3OUa8uLBgGyi7g3MT40gsDMTqCLUhVnC7FAVztoizuszN6Bixe
baq+d2bfHD2ZvemQtHwOKJZC/7Td/JxURuggQLctBE2onki0hUWKXB6ZlPSSzmKPar5V1+55bRMJ
LaymfcwfNBG8igEiY1xGwGH+20VUP/cKhIWlT1X/ita5Y5Te4Qvm6wHysS63AVgA0dvHqVETDQc5
8Ms1eB6P41wpptVKFgFu1mdKQTIyBdapQatE7f58UnhMTrBfk8J6MjaRUq+0u8NJmKINytGTyPo7
GS5vrvusIB/3OnPGDNRPg2v0LWdmF2rklpM3LoYPdntmOfP6P+fz798Rj9xvXmo6xHkpx76HM9v/
XO6uNCIbzMYBVCsl7S3XJejTzbKXehjeSGxv7El5mEn62UzdVJZm9PGF3u2WHhex341PkZs20X/i
GhoeLqo2hVc6p0YfOR7vQgdelCqLQMmoScwfswUmOEqDEfwU/2YyiQNX+GQy8KmxexdyBRJFKjKv
giytIl6qerQ/GOOLH/gm4bhqdicM5Z1kEhrkb16R0QcC8hE+jX4rJCOaAmeiMT8g1fS+2hkTp0xo
zaThO5kJ109l6xj/XAM9h39Owb+EQZDa4D/RyWRe8NjHGR/VmjWS9q41PnFoqv3fEs0ZGKFvm+dP
5m6+u0hG4VuQIMV/RHuwG7yrmomAjH9E7YvkrAgqzIA4BS+/gh/BCHLNfyciSQS6Igq6Foauf0EW
rdpWStoveyXdLzeRN5UlUZSbps7JSLJz0sEMv25aadcqusx4U6I5qjrSXx0ASnmDqi4nMXy/aa6b
7G9J75DRzMN8giAfQJo6jwaSH6XtHPD1vI6TTTFLr8Cz8N2QbU1DuXN91SW9Ucmejh1kA2jBacQX
ev216gYgPIZtsFBx1SaLNZCKLu4WHr+Kd4qGP2Khw3MmYiYff0ksH+AFhiWU1yKH3vT+pP2BDgmx
+LgONZEpLSk1GHqjaa5xsm4A6JXx1cCyLE6nBK6p2pZg2uQbiGNUDWyTuDxK8eswvxF5vJnCuHka
PySXAmzZIncwtjwQtBKxpN57J7vDdtptkL+xvBeDgJYeS5KRlesFbD+TK4goXxU4xcToj/ZlSIFY
xpiZbsBxWEinnDnaElQVFwRGqhHAyEEaDU0XpNKbPNYXFKABHtM4e+i/3VOxLXDtwzZsVthYCslK
O7WJqbAtZNoB6Op6GWHxHJHCxLYTEZHvaBDCoI0ljRolRZVrNFt2cOeTN5bB3OKBjFgiplrQQHyU
Ec5cXvR7pCPZDNF3bfnWWyNoxubl2FP4Ws/zlIMRZZNx3i0vLjhwXyw4KHH//Kizl1J9qfojk4Jq
3Ay6LNicuLQ/VrRTTLIv1XlxOyXmGS8TWRO+LMgVU97zo4ZA6q7AxkQmti2/KsJ+IarHMgE24j5E
n5vBRVxfXVOVB9moXMRt4/n2D3BpGpyLf8wVfXUjPsItDS4UkuOjjLj0HnJfFRsvKjhtMRIXhZn2
hGqSqmfyYXOoZS3hHmIkqaBtmOyMt9mduFaD+NuvZydTYkIdC5suea0YbOJB0M5PKSqF9wRpuQ6H
DMugJ3IAYICuTgXr1glHJFNdKgKmSQuov5jWyfFX4z12QjZw2wGCyffgq47QqFDkUsPndOacenEZ
vZ3rupXW8RHlOWELv3Eej9ME9V+0/2fpMRPZBbOeLex4UTgGEqt30QEQ6ddrPolb0ZXd2EKwckYd
yFF0NU6DFWOEz+OX8b4W2i2S4d0FN0RxVAET5Gd4puJi/tZsOnjIsKxEAraae1a86uw/9HanF97s
AnBFy1thU6KHSLe6z8B7ihBWydCDDHz5QB++PrSHhfcHVJka0Ehx6vajH4nE9166tKqDSTus/w4H
hzglVTyhjr1RNl5mnqTBBh33qLtBX59Ud5FzqN4AQcqse2P/Up8WZnzS2b+nneH0PP7LItr0GryI
VPB5rY04EEu2tMCCwuPL8P1LRKDRIpnG7LdYlSk1d5/cVZdY3fBpOfNRFRYwpR1HbO6eYk5ta7Ve
F/xHAbm5bmRtG8UAH7JkLTiNTtAtWRXi08FsSw15XvsDqPbwuXLkC7GhzcRkbV5OTjW6LGakaA/r
Bw1A/ZJEolRlM6lV5ORHund4weZnm3KrUu1NKAno04mJplQvJ6DAJewp4I5+4fNkds6Le2KNGdBd
K1loVgBV1fCgYiIRiVX9oYpfawzAQHE5+22o4TSebr6s3+AQl7etr9Pjku72DDGfTtFs4SPncKzu
sgMzE9Etiy0TqhmA/tQPG9xFl2mDDttbtM+J3gK7a3RTQvUEKVryfO1HxMDq+pG7PfcGwbzIU8Vu
GsLIdcS3/qb+BOlAqRFk0KdFJVlg/pLbl3zlcQuQXJNiTKrJI/zdxaqQmzNBdJpt+D7vAV/knYhF
CSd3r5PrOsWviL/SOB3MpBIylbr63JFvvFb8qBBWCEVAz8exF4Rd8lgQnkzegHJb+tCoHIGn+BXe
HliPt/eDXA736aE9qqbJl+PcKqh+puBY84gD0lRP5EJlwilKUh77IyCvdoyx3oziaW7aywMG6Tiy
CFY95J0ssYkDs3lygRLEVcML1XOQ8+6yxH3U7IxyxQqPXLT2jkW7R29cSfKQey9CByIoJhPJypEm
prY2xGUBxH/oD9joOPDDEEcUemlo4RHEsuP7joTFM0M3tJ0NxPD90/GtEFYba90ahBQJi1D6g8qG
QqQUd7HqsT/iorw6T7I6m2vfklkWCYXjOcmEVPUH3X0576++/P7zr5FxjeZlawH3zNdpZ/RYgBQx
llbaZrUQTo4P+4ubdbALPLK7nbKjIqXu/vIj5rINvlHyKJ4tu0wPoJR08WkorGW8DQJmm0WggnW/
C1UG8pAgH0n0atjlo83jB40WR0Fntv1mX5BrZqeYlDxCxTFMHtQzQUnNiHOszS9chCsleQbOWavX
OjSA2rnRYvB4+lwzZqzwDaYd+8vLYv35Mc7+NFHOpIO5p6GYN2vhQc8XrkyDrSrWcxuCyKOkFu8K
IrnjpM6ob6/MqQBhVOFyb0n9Wx9JiYI5eZKeeq4L+tpki9rJpLYlstlkF/DZIpuQHCojy67Fp3bX
X6TpwO/Qugs6iU8W6/VmObZzqge+Wt3hzPebh+3IBWHqXa21T3NXLvSDwRrGwz0u6K61Qk6OfEPK
riESDud5SwmLlmlUxlr3+tQCrqN2CLHEKkVnFGywoZsR+EvgmkEPdX168c+WZ2WhDg4762E8/Qs9
5ECDBFjstfxtkbwCz+jFWUp35i2/qSNr+CAxzjPifS7UpLQ1L9YwEDjc/a7ZTrQnXfPAsZRkfjqx
yi6YQt2gYRAgPK9fPsnotiKn2QKkxnSKbKC8dXd6ZF3kKkf0jmcgfepvb92/uSLsMP6RSYls0r/p
y3ZZ4rxMY5PS6Gt0RwRZLNUAoRpHaSoyGzhbNBHzNHsn38o22ROPV7oBWMzHT8wbzpYYV7OhWzxK
qkGpvIm7kT03KBW4h8uomgcfDl79Mxa/UmFReOcr09yyYLr6+F6AaoNZHsK/s49RiY/MrSw9+oDM
DX/PNeOjqqXMv+zsR7qYE0TxKgoeo5m8btgox666Dm2zcFyffCvzPNKy5WvcZgst4Oaet43X2DwH
HL3feES+UGaqIWzoN7rSb0qn/wDF+fVuIK4cOcA6Ovf00WEoiAmJRAV2L+pjg4prl9/UAn0B7hOr
Vd74io7k7HXXjLDrCOibHuDInVjFwonmVB7GWDR0KjXZWJJsM0Tle9EeozcJxU4gYyM7iXvgEbsX
3ZU2uy0BFUmOOcmYAQWAq0lsWWKJPoTF/ixByC/nS/94r1NmWArUACE4fZF0AhhgaBDXjbYSq4ZE
nhFoAlgKFWrmDIYONB/044vAlFiEER4hGx9Oe0UtGJPMxBzibZyKC5hrjODicyOlN+ABFPZEXMqu
1vzAJJkWRbHzp6wNhWv2zywSg6U38oykDa8WYyflY/en9hSFQ2zkTyYWgST4OowQ6UAStkj0615S
R/glvNmjwNWSmkakgAMJYbfai1e9UAs3aeUnQ4OYdPWHgVnVVJ2drzSgVdjJILiePs2avLxmmO2b
ElDnvdGk2nr2MpYWZKl0WJsBJoXQwEzR2QiXa7ztTDVFqKVWmhdUlv+USA/1G0PAJwpC+t+rX21T
9/NVN68vVZfuPvJdNXFW1+utW7f0zZTcRSwVbISaTaaoalCrJ51JI2QYEsE9p5P1ZK1CA1qFUFGB
WLkp86XBku+7wFA2qQBZGKokKSgE8qPWhqU2JRN+L6ru3AJVZAUNPx0BJi7xtrNQ+KKQpI5DFBCc
qy6ZOAtEX6nU/fGkACPiTxL+tqPGz6iPwL52wn3xJejjEV7QE4Uqm7UaK5e22cH7KMrM2QqVoXJw
svmve0kAeojeDTHENv4VeFZboz0WVydS2RQxkrzxpSVIa4wyP7b5FvXuJCQY5xLQtAfqH82zUw4a
qKGGJH/QzGTILY9DDQVne44nqJBtSwF/kEQ2KxJbPhJ3ge8FqSIJ2quGdGrOp2aK9now4vJC9tTx
zHzGImZXdTF9bM2zAo1P2dY4KfcMCdQInTOd9qSr9t9CtMsBmKLOwG5/kyJkNxfww5wbNoZtGsXo
0NbyPB5gGpvLfQ1XXaeGgzYtBtA1qQGhOpxG6Hy6jmCWHobfOcJLE3HJ+xIq6BP7mioG55SmAxT3
3K58eOW/PYISKs+hllYIib7gUA9C01kGldHumg1cguVXbWdiMI+yVw6rwoxKpMErYPyBldO5cZhB
tIUCTt/xC5Cvk/YQIr7JzanK5yt9zO/wUAoBBsIfEwpIQDB2m2SHlD6rvAs/3D3oMPGPari7OzGR
ay0moQNJ1pEph4rwd5dVEKVMt3xjm9bpdN+S5h425PkLuvoUb+XNLZUWaRvIbEqwcLpB5FzO+CPH
4A082LrxxHg9inn0C8fnAwxu04xOXVNqUmGBWxzHdMxFWeJrvQkBwYduqpMHXQ3oMWHQswRxNPzG
JquQUOfQNfqU9j/tEVndSzvxCgkneG1okAmlu60mXnljsLl6hm+bzd9A1/fpS8uBKZ9wfGfYOG0C
RDX8t5z8fM4hdS7T3hyVK0x7Wv2Bh8Z0MMIMeSWwORlN2P7wxO+O0c6SG2fb2CDnZ73mzvd5XYgz
3oTE7HSlHYnp6r2oYuWpboHa85Hs8c/iubcZLKcLRJJn6CteOPBHMDSxh+6q659+ar33ekxEOU9A
domA8/CSTp0MD9LXm6CooDWsp+V7z0nVzXlJc6KXeWVc+0UGWFScCfgA4HiatCovFDxdHH87Oqi2
C4Go6218RRRDV5f5aH9U/oMqG+DoWNzh1BwUPkoWxdjYotmQjPno+v0aF8IUfhr7c/eV/F7lH40U
ijl/ptGUs36vhnW/UWR5y7QX5ybc9jRotack+0RqBxmGKNgtb/y3h0I0Hxt6vCgmJfoDdmaoFtzK
u8BCTbEuBlW3Xsgrw2GEyJGRKOHdLLnzUzhErd4N3RaILL+eQKnuPvLlo55P0Luty5onaYRJuUoG
r66hVtlCyHS2Bv3eOtu7CL8xS+/t3xQPs7HVBOvPpFxghicVdHuVYaVU2c/pZP7BBRN75M9Oih49
GbMLLvtY9tw7PmlCUfh9YmgO/nlANkx5SgVlWwJ742QX9/78Ter/VcZ8VGLmzQbZpCKchZEf2W0b
6/++N12bTaAzPakF/vnz0jwSTcOLmGODDj9t1Iw0RHdEFDNX0aUjPFfMMgTSn2C/pxfmb75in+Gr
NleyszuAWBGICYXM1mCmQF/RIq5bepS+uRjAULxdq0n8LBZybB3yGb9YnM+Q377JQ9tHNPmHnAvo
lYeh7gIwqM1nI+iCJ9RtHg7VE510jNxZPpFhcHwxffwTRiB8nMLlAA73WKnnOMJxvy8LoDohNRcw
SQnVneBzJ7fFZCEpNtX1UGsuw2+BiZhmnLUZjb1/sl5+GfHZpVs/XLKryyZiyg08NaPR5suD+Fxn
RisS0U9G/eoeBjayPoMv1PZws2Fdm/NIZ6oxsggkad1oYXCluz8CUdYcRDhVthEd/eflSY6Xcekt
jC0FhNUG0SREPE0Wq1fD+iE0RzxicChcTqwoNrceL8IypWHw5RgvQM8vj/qst7LpPykm4b6kImfK
wEgdpGD5aIJS4XhsyWTkwSYfU/zUxYoXdrXmdjMuVPm17Jt+ADjH0F2pwfXkmNCV4mZAJyveU63H
hcYfgDfvWazXNcRQuqv6ghNc20bw86NF1N2Q6XRC3ntYlpnJXgKmmTpfK+zK9T1GyRpzmWa40OBk
FrCKD2/uZeX5b8kL0AftGQqNNtBySVUo0PniCXmJGgMs1j+G8HxmxaSAjLHEP+1hydF0ZcU0nUST
wsTSVaZyu/14nNOpwV9rg3H5U2SrfiA3q1MPCTFf6TFlUphDl5qNagNLyO17G7HY2BaEjqQPtHaf
vGPF+4azvvaU9P+EC6HQNCvxvZ2Va13juH6X0k3jGTczuxdeCWQLieIG1B9GEe9LDkObSlTi6ZE5
L0OwMFjEeRVYRDlnpSE2S/+F9+e3S+rezFg7yREiSP2h2SNU77oazXrHauAB67YQRlzhITmP3vWc
8QrRv7g3S+WCQEBvk7JbGL5XZiXeJJl89y9+PTBjZwPeifOB8YwaB3a0yMamvf4n3jt64Wt9nqZA
9EaSiFoHN3ZptkPWR9TR2mR9h0oLgL9CjXfZbnCZ5ytt2ZhkiWuyqumfLzvS3YxJNgACsMtyO5kt
wFBTGrnSPz07GyC+T5KcAjgBRwZmS6cWGYWw07TN21+K9lSUot8jXt9262bmWrrbzNTyZwSUjyN3
+2ObcJmgZ5lFIXGrNga+sx/hwzBBQAwPt43u7lelh4sMk7l28apmqV17a2ap49d957/KMQJPaT0U
zzB3CUZa8yUGof8j+v/WztxnLHRFl1JDwj2PzqjF1x6aw3ZEK9Ws4J+lYSIo+U/51H47AA9tD/dk
dcfNqbHc4z+/2FaWuuX/Ct89sq4yidgEdsdanRtwks+niIYurq/mPdA5cHivv8oIa4YoX9DcjMxj
oe8YEKbdW8kgrMc70UXDuLZt0jgu8GqMWcwUssddgdHH70nO2p1XP00jyR6wv+1vKXnVG+lAO3GL
bhDUyjCI5A125+hhfvhsob21tArAv5XOWGlC4m7b1Fd2SWIK/iYXOqYi+IDuBzq0CNUcKM3Svd91
ISnKobMq+eB0rGQTsvNTtmtVk3xTHXurPaBoeg2Iakf0sdmIg9JmjEicMljo57CgrlT7z59qyIFu
l4xZsvGS+sVj9I6d+pB0EtfQoLWjZOEFYcObbMWIUF4G8/ixzcobwVKCOzrQ9dRNfDuUkDg3Pdjn
5ELpfeAFmsWRi2KSjoqKoUnr0ihYVeDFcs+jlBVrzXhk/b2/OwR79/jVQkZJnIxfVk3os3L5zTBE
ne4FwYeiaxJjvkW3hA/ffoH4W8MQ21vUki0vepN4odesZyOsEivzKaVpf4YFO4io2e+soMWl6HKQ
cNfEQ+64rk/8oWR6VYec0S3TwezDfTiIz1wcGuNz3zH1g0rWS0C+2VKJdx6qN9dSo4KI5NMuusMA
0ipidZ7HOhkI0YUI631dBmh9F5n43dgNtJi/kosIqKW2HtFlKvsKcLdQdEZ3ILGCb+4oQVGHBPEV
PAxmNDYj6MbeHJyTPYTGuBkWRQc/qkcZ32Vsoclbh23MZRdyrQCLPCTkoAKY2oRJyp5x8KQBU2wD
lzXKNqavUv0zzyy1UzRy0cCqYJ4EwHnrNnOlE9Zx7kUaQGJDAGugFXPmJmq1Qz6U3jScT1OKMdBC
0AnWqlOgUMSdxXo0RnvysPaT9sFOMjfABGJaFiQoVZ6+N9Hm7+NGU7V9mMVMhGStyPb1PU7pyi2N
NunyJHlCBauMuRNW8uzj7hWU6Tr3YCbpJp5L67RAkGX4T4/I8GjWArL1CEmQPZXztKQPTVfJ6JBk
ICCCfpnmRzh8dJIvhqFbGmVq4XJK+zi2xSZyRMAs1mrWczC+x9Nm467R8NSuk3spb+f1Djp37hUE
F8u4gjZQT3ZcXDY0uu9Lvw5zPktoZAo/BYXhfcWUMQtHuunxXDU3Vu28HCXr1DxAktLM+dCQZg2C
JzC1Rd3y/nyiJF9wBKEJ5Z6VuJMVebvzy+xfYY8+gXRn7XlaL4PYA0tQtu64rPyt8+rLNuhDpOTh
jCkAYXDznb8cCWBEWJsHLz9njlFe+X6IjMCpm6HrRDi6XHQXv7ASxEvqy5rVnI/5H7LZrj/dr6sV
cMah5tqPUU7bI7z3umndmvoNoC8YYJhHXVRziwNCK0aTbSFitJJqS0U3SKpqZthK7/vHVxRHOUpl
L8TiQiT41OJEbyrV17hYqSvpFlH8Nw1RB1ZHHium4cDKYjrF1M1gA9upB9zAEkkru7gySZGwGWYW
Onj4h1y4lMDqpM2LlXtmH5IV15BVIOaZ9Ytbbg/Rw8ow8CFwphpgLveaWaEtI1Q9vCQCcqgtuZSY
VrynGKXW/VXPsWxAeoLU7iC5gCy/gLzkvKwUTFidaDGe27PRF7a0XHpD3sATkyW4XuIfEfYZ4GsV
kG4PZ35Iwy3fUXTu0Bw9VGH5u0DulIX/ZG7zVYCGuJ3NW1EZvf7UVgKGKrg2zmaWXbk+kJdaRTpp
U8zpHZKoEBqWVEGQSGF0fKUzBjBGpE4Eh6aOTJu8bK7rDBZRMzUoxqp/zPImjGq/FkG5nnboPQG8
o+a95MExn9phKqg8hbZ4yM2FjZWikHeBTNVcrhCXWmsq49kH6F8J4ophClmbSKOjJtdaICtPhCCq
2FlB+c7eD65opjsaFrsonHHtPc4nN03TXJ5G+VUzjq/TDCG6388mauygwjGYmfd0LMqMm4l6K6uB
nY2mnp79UliEi2MR1jpX75Q9/y3/P+/hNCxhxwGX6rxaCLnymPRlFbwODDLkhQZIbjneAwUqQ4n/
EGpEwUSFH4VDMWaLt3k9FGeFQF418xsHZHiH9p774K3tv27uOc94FZqYM7mICdBNdpVvwPfma3bB
WxyvkCqPPeAQhO8vCZ8yHdqmfN2Hy/FRa4RrQtRIcXlEr8Wr1sk8NTuJoM5HRBgPV40MI2efAFso
aMsD/PJtSt8lYeqO3hY3BEvuJ2OQQGiqVdBfMVQ3er/jUJCzdIZKsmSFR5ninvn4wxb7daAUHA7/
HJbtL/yzgusQvOrfY8mnm2Btpc9JmlXAN+TDxPCUxGxgwBJocikdJ7i/DPUT+A9k/sWxlE5otnBs
IQnVqJ9xQQnVZ3jUZvcM0ep4tQKxwCIg9+1KQglK8N7bqcmLK9+vbYOPRmWfJqf9HI3lQPTTa2Ez
fwF1n+hKr1Y4dszLgnPk0QV4ZZl0D7XIAzzP6TWiszXIT30pNovSIhND/HX/VMN/4g/dMVzFzdrs
Ed0/IF4irs5sqhqZf598RF5uardqOh8DuOyK4sKBhcMoyPBGpRITorVySS5WqjUU7YooMKWHYwm/
Dnr+udrlq0/xBc8rAhlCn6rlcSUIm9oHqaywl/d53kfMPtKIT7YL70FxAPorqkWNQluxcMV4T3Ss
IlGlpPbXlQn+fi55DpITWy0sPX18i1l6LkF62QR3iOVVUozzAFZlLdqguvWUSY2dcvDXXkma2Khi
qvbT90YBrVuDjg9GyNbBIvmDYb3lghHmpn4/E6rXioRzbseB1o6gvtevmR5bBidvvr/gTI2RnwRY
aRkbzE9kb2zuv2dtFFJ3uGPQDcPrt4lYNyKwHPEnauMsewMgTIkakAE49IHOptc8nIL1f42xYenK
77E1OuzgpWlbuJLi8iz4nN6ghhydfhWFWVvZSAF5yP+k0UaPn4nggstF3JYSawdoU3rfdduol3s/
4bfCslIBxB/xeesKgH4Y8NfLfyyozbZIMsUxY5evG6Q3IoWcjo+/9hh2shq/QVqDDVeSAtLoJD1i
//bjlR9B8tQuVMQWsKUhu4wpV7hhQ/L2AIGeRZRmUS9jK7/aBT+TpexvRmbXJijfjuif0g9omBZ9
U50ienHHuQnKAqUzRZ0VIhnjegFQnlj94KTGv35RBUmMu7oOomBazWCJmJk2HNdhYr+Ggw5f7fOm
k+veAo8zxDp+x6m0XvQH5EhVp8yVlai57ZQ2s6yTkGbn5CxKI8OlnCA4ktixOIucthouHYneO9o7
xljSsDvHWZW8/30GW/2oXZpKOxKIAdooz862Dy2ixuhs1l+4WK2BATwX13QG0e8Suynn8DvMKAgu
bVlcsBMKhYU8ifKB0oNkhSMdkIgZ6INP7MvHCWjVIkmAhChYjlSLWCzrIXEH1GhpOru5rP3+9Csz
3OuIrDrG9vdiuPsIMJpBSQJqtdzt52k5TsOh5PTe6gxAwpUT92KaykKFx+L7XSInIIGS/sZd/9dN
HdFtJ/Q51Vc2d73OPkBCr82M0Qi6xpDe7Ndk0Wwkrxo+DFexHKFeKxKs8Bhczpp0Bhfqep5dWVRJ
DV6EWXvuwx8IaO4i+/il3QyS4a9JEHfU698VIkKEDbj3cGLkaDi20BZORbVEht8jc/ZZS487e1xy
nBznFmNthab4f+Mk7AJVTF7IvJT6WOUwDD803BEB0EyjS/5ZCi8zaX6iph0ko41RPZ42OZkdQemu
61kkJFkZb640i//S1QR38mOCWok8FiwnxaOFF4CX4HOGg7gut6q58BjqOtezcEBLprdnyaVrrdvT
D+ywoTh9nZIwmxf+LzPVYTuNAxHqjSCS8XWi2qSCLF3RItR0BaorUd73YBGKBlo163X08GbNsCFD
ycAiwG5kYlBeJm4nQETH1FIJSpO122KkmvEDpuyQfethmMURS0WSJi5CnPzGIv30xS+1uH5xRN+Q
u+ELZ91mfdf/1hkfi1izJGD5y9jPmKn/qZS8vXbC2kmBiv8jivfxQ/Jq+l8XRImzMMvD2g3JT1iM
42/N4YWS+mgdm+J6tfyTtf4XP0/61js2zr4GzCkEnKI6AOXXy6gCFnRtKLggIDgjdFtMaBeumr5c
ug0H53yrO0O8/n42DBn5InvtzKYScOprzS0OEmxNtudNuZHrt8TSzLz8yp6+vMIscK5Nvn6Wlz/i
M5/li7dXhxYXVXYtg429Ampv7VenAza50BKO1nQJOiv37aYIEg/55NOaBVk3lKDuGtfWUuyrN18A
Yf293jR7timiC9ExPmCQpPdNlr5ammLsd0LzdOO4a0OxeZXCUbKBPiMUosIRPe2pRSMmhg1ocv6H
WRxKPqP2bRijdIHyj/xU5uajWVsJqK62HscEkVeRa4CqMDVtAX2NeIR7Fbu2jGwLSqTT81KPOzkn
zMmcGXSMrHPkNLLHYt9iwe2kBM5u1mVtvVcZ9wagiL/yEiWshD/8t0wP+FxiceVKWFahjVwmu4Se
X4louwYZ98lvpC46fTTHyADuAo0d3SwdqXhBYACnrya98/V6ixRF3Kg8dlYaTs2wPko53eNRC1jD
Xf7NbV/IXcerzW5zPwE7f09neZVmW3lIMZkN89Vm7Iv7ffbRP5h6BLmOBzyjsuqJJKvuohOY4ZoR
L4jz1m9p0uJI9IiDlIvtva68EUub14FIFX4Xn/LDiz5c19aH9rq8clqN91ZAFXtsHr67U0kEHJpi
a4Cxrlv8nGsKfzWlVbnocFC08NJqz1AHyGUsN7OmtvNfYSHGe/3+QiAD14HYUvbeNRWMGmZlClvS
m7Ct7VL+0dFCcOMDH6Bjj0zwWKcbwUQexOKzW46hTfPRUWwTf4Ru6C7EnQDf1nJGxj7EA7f54NZF
SnfmORgaqwX1sk2PE7k2Uy8sn73dG4vK1G5dvUbsdOUWFkEx4Cw15ML4VsoemzK+rxCm3hP2QDOo
pOeILMNtl/SrwSGvFG0GqxAo+sFPeihuNOAPMI/PF/d2tcB0RUBie29QdWzRcCdXsx0EvyMmAMY2
bTMZCCBZrPr1Qid3aXMswT16qZnZIKrzG5WUvSedO8WFDGJulj2BQuBu8E57E3uNviBLm1OzsD8q
RyI2Y7YEn78nofqzcpf5vYHSg2z9Xu7VR5sVxYlVX2r0XeWN0NyG1b7U8ZJfXodJjCbaGm5A+eiv
FuGGkVI5H38BRsRw2ZA7eHI+s7CZD5oTY/5TwDW/e7lky3wbXungTTGqP8Qfh9o9EuB6SMwwM6fd
zOy8cg1ABR0qhfi6baTLn1Jy2oPxrd0Mi5EbytaEXYz+1JfyShlK/D3MRurs7fg2PK/AtBUVLHpl
mQj+Ctzz9FcgGBhsYwZcGt+JLkS3u2mpIhKQZbbTISJE76a8o7gADN70qCaBmz32i+Z8rwiR6n0u
tz9j4vVxEy5fJ6gq9o/zjLz5aE1duQ8mUHvlobuvVDAiYvN4ylE6ewtZE0BSneAjKy0bNVLhNyrD
NckQsf2wft+uroq0rL9PIph3O+3ldYtwy2ijXMwVRhpmb5ioPsSv9SvNz3DvNnsDZgqT7sO/5HeR
GHH990cYSmgjKuwxJDo6Oi/AKXHsQ0ip7qptAxw2u0ohaDtIT06l8AMRVV0O3Ldi+jmiUgdTOElv
s0iOhbfE0nXG6BXCVoLR8ehLEDsAoGnFdYO7wyzZmmYKy64RC+kljL6GCaNso0t4tSPbMfWHg5fQ
d3W1ZjSd6LqFrekni5guOqdAjAtPnfB1U0FU1xagK3iqGa82papbvkgWEEhR9NCmzH6cKxsC/gFf
EY5QDftoBHOqfrN3oBmozGM3LZJbhy531eGBZtU3scZ7mCIR1IcWLPd7ZZVClRkoPenOB2wozled
1JRfkceTOO+AoOZ7Ua51iLFJ3bHzpAQMezpJfdS1HdkGUBrVwUp/+by5RooXb/DiK5hAh3B1+rHF
ovK1ey1koIKCeQ/+5l/r1Y+aA0SCAe0m3SJTfrnhpDZJIIt6wmbmuJcSicoEGrArJgmb/JzzlCUE
anbjQ2CcrgLEIQNM1D3MNlnDXHE4PW5QXl0pRmN9ixq+cwNj6nIQDe3oVVSSayIiL4sv7cKTRv8Y
/23nyAo0K1fAY6St95+uPZimnl98em+f59etSEytPvJXwU2DFxWiTVtwhR8MIu4jDx0BIwppw638
9260cE7dxosVGCcDPoY0tEWDEBkztKz9ACLPpMGAZ1QcberT0od6cRnkByUO8FXofLQQtNwyDxzl
tG0vjlIay94Z+2OZmhKINMe1YrQ6Bul2xxMjUrNNSFdRzsK70T/JVvl6KSTSzOcfYeQZHYd0FR9y
g9eSwHOaaHEvcQre5fuA/HZHg8QAXW1owLsKH3qHMyItM5YbpCd/HZhUfq0e0Cg6AWozmislA9AS
m518y9F5IduxxAwCHdtv52bXnn8b6y7lPAwno/tR5vCN0AjvSUouxVdnsq2TLsmL7awlTau+7n/W
Jq/gON7RP5CWZyGWj4GaV09qeQ8F9Vf5yyZnji22tj6Oq17qVbctDCND6TLZFszAJCX892Id1+AC
IOGZCr98tT4QD2ZQ8u569uQ7l2eUH1uijA4EnaN5m3vMX8b3MmIL2Kg+C8sN3XMrTw2W5qNZ8SMg
al7mxAExCzNaynF84r513J5+Kekzq6inFBoqpincutnGUccpnMHU5hwB1XDOdtCC1SNI6TERksh5
HBQc1EKdzBHzyLX3/2oCLaheL8XJ7esyU6v+ZkNmfvL6v8850+Ko5033/vjo+VkikqlNnv/XKcFL
mhP8WK+9CHw+Ffc/BpjRy7THulV0XNYQKmxqIuVIf6CabO+YAFp8XvpY47peop/zpK6lGSdwCWGa
/MVxrZRBeXWLVYiaL9SLLL1jPe0lQmRr6HY1mxlCkluVc9nWTakYMeZZgIEjIeujE+XhQGAUfjpA
fE9u7ddC6q+L5VdVWP58bXblPca2RTFjv/EWR4CgksfZ29u/gwk6/ox6fkugRG/gfbshN9Zt4xNW
ofLjTMASA2RkFWz+i8Xz4PnX17gFgtdm7J7AWmarbyI/q2WWPC9kJh9PxX0osaXttRyZ2UL+L42w
YNt2/MsbWCGKBuhNva8GtuY/godl3mO+vSedNqGRjfWbFiTt0HV9edNp9MQn7+uA2AmW8ZQPf8O8
tg6uRXnYy6AlNmzCg7pUhxQrVia0gP6A6ptp8wfnCS3Cv8+gQKGhB030NlgsPiNSvfOu9QLpPI5p
VbhBMsLN4SCTWdPIRdrTlDXAjiA2s8NQRxoy6HolzEeWaPPSFJWqmYoAi6J//sioYv6zIt22GzE5
8tqpU0OXgf0tnf/NLaX+yW/kmRgk63JqGpw5GXS1W+hx+Ox6kNzB8PmHjgvtnkU3rswbfQslGGAY
2bzbIeyyxEhD/NpFaXfJQbHKv64SqEZ317jGrgsu4aBVNwK1GaGW3l31V0A7YaA3GZNf06sNfpFh
9SCxgptIf1ZNptdKLNHSC6guNqSblLQUIR54oDOuXIQ1hCDka/c1EtTklPSr1edXR7Bb9xzt4RoY
+qn1m+AUmMObvYeYjnse/S7DSCWr6uoR0TjlAm1q0X69tnSOqyNdDx/9v9tKEJMXB/UElGtJi1aq
DD1XjIt+mWwQFq9WWcKMAYae2RAolwdqIFHxqUMo4wYRt8O9qDY2Fftfh5ppSXcGZJm+z2Z0S5YR
0twC+MYjeq360ctY7Ha3p7/OUV79ew8dMZ73YxIVVmgR5STG406YvxqkDYic7JOOOfR5PF35pCGm
xKwZh1S/PUdEFqQ+jcIU5QKD+Zp9q02+lPH/34WpGcVthrQd1uXcqyFP0TKgp5bIrhoAsI+tcl5X
SJ+1PuL5jVsOl5ofSNIkvWd+M/V6IDRWS0JRFJDxuDNo/mmwktXsle0UTakRU3sabQ85v5Nn34mq
8yv5yRdkPIuVgOAk9x6CPnKxQUZQ8W/3/pSo7SfYDE3mo6FLcNIuJxNdVOSMaAJg6zx9jB3ZZWyB
BilnbSRrKh99639k3lnYwL+MebQ/snR9FwHTeyI/7XrhQfuq5wze74YRJjhlvOMrdRo0cc/MWvic
3QZouQVnx4vAkxgATtHaAyYaHUI973VMRP6kGrmHUlOty/aXhEqPtvdix/b8fHERXNVSlVP9TEQK
z7Y43VFNL27A46T+MoNhJmREtgSs5kw8P3bT7nDTLFvJo78gaRvLZPYJDbl4rAk3Qjt6BNB5xNX4
go5cMhc5vf4yiudSFAERhsz+qvLQ40lI/EBx/H6OHXDmvSVB9I0h4pZPXWHZ51eYgaxmt3bDTEXj
BiToG2EN9aNiEDW7a0mAy9ft2fHI0VAUzZUviHKZMp2YdY5F4XhdzqzN/BLYUfWfIND3Sh1JHGEk
EzXneMiLAOM0usoXoYTPaDmO7sTbcAH4nlE5gu9n31V4akAZXAKLZTGAiaWtvzITssTlXYiGJYqT
qrSUe8J2q5spIMyv8ys5egy1TEGLGEccVv9S27X5PYvv+mjQNnbK5x5l5o9rcljupE5eYEUtiEiX
z9cjwIYIU51R+4Auz4WdYO/FtCmV/Etcrg0Q96k4OcWSBvSR9SoJr3sDtA0+EB/HQnIVQ03g9A7o
ojshHe9bupyCzA7IRZ4C6rYxnoWJ9Eg8pexDjCOAk8hW44cSQXqTLgrUOZSHECa7cCK6cLOU+I7d
XxV7rXIy48wihHFVmrggygLvb5BL8AvX5pDSwOtLjJAq2FcstRQfffFjg9Q6UlCcYicrXF+K9Y/O
g7oF47qf76vAjt3RAx48J8ps9Xv/AQN54xcD6hVdHNlOOGDWHyKD09F2pvws6ww/NepRDEqlkZX+
sbaMqwqzKBLWl1BkuHXYeXieMFNeZ2kelxfHq7+1XOCRd8WrXBFXiORraOqldlxd0U++jbhFg7gs
IQy/Z7i//h0KedmNpNo4igPD6djBBG96wmdybvLT7DaoCHIIo34oSADHFw0C2yHFqG2LizcZz+tL
PM6flq+nO8KxDos7y310RVbWfPb5sJBm4YVPnIfTmyvY+jQ8Kp6yyNs5kIhmXs+kmohWghmjXiJs
zjq07ZquoIaOZt6QnJq5caGpybwrAluMMMItehhRUAzELD4031qFnPOHmxlDWFBw7ydDi0SA6ln+
5LrL31g6qDr93a72d35fVQ7NGLRDF0S/THWR45dt/q/u4mxakcbSMlF7seUhDZ6x9x1lyBmOwr+f
dq5i7/TZ+LPwZFtDfofndPuuIlIrZ88JAehBMTdii+OmZdUh3UcK2hAnbPijx+ThS3siDOJNO0DL
cLqtk6O1yInVRV5RNM9Wz44rdQ58hhcCqU/c9DnQL/V+7sQXTdOQM3hDFjmJfpZb2zLjTbBJfmH8
jYpaiFaZ4osD+Xf4fIGRJrjA/NOQp2zRvekg7oABdPqYDCsY7NohW/LZfyIHXHj89CgFUH10zmbp
MUWuGRbf44t76UDoY2ndEGYW1ohRrsAwh30/pFhEhUZwKzPZuU/6k5jQ/0cDStwxX+d0JzYDGP+L
OHYIzPt4mS0RdIOyzrNn5eLnx8oKY2LDm2b3LZkfu2uPm7CuEnEzZTB7z/CK0jGuGKOJ6dpsidKw
KQKebICfVk3yFDNMbeXV7lXP9crPvU5Bl7f5E2eKoRwN/IAy6D9ANYUC/t4YRQRt8Z5TcrgixDdG
VuKiLDL3C6q70+cB9dR5WybA8nadill983p+r5lz9IVQGdvQG2GqOB+RWnnT6Q39LcUkiK5tDh/d
EObZsWw6ESoniKVw11u7ZCb0jXXyCtPcf6Y6rCTHNEXfqWU70CaNufx68g2JIxw02RtyfpySO4bO
ZhkjkqKbxrBrC+2rBrLpmkYURzXikN1sDGTEIIDiHlGpJ11eGazSGUAAq7h7DJEmGBaDZnVm4T5G
vj1PmCINvJ+1yBRuV9OrOGR1D6pLoZT+4l3GG1c3KVpSN0srDBCJdhAhAI0nj3xVSx+WHRPeGYNE
8SQWNZsWzTU9cGQuCjWcRQFLm+YKG2ZsTumkaqc4+x1BPQ3ct0g0PSm6znDMelJUkCgWIxSQCvik
+Zw+o3mIESoHW+sx5jmY6W8F7wad+Ix2kSp+DrwuUzFpHirH/etrrLUe3omDyqKKMVxElZ+z0jVH
68hbIdACLO4WzcRFiTZDf7D0MGdnx8dpZqBB/3M1vQcIJweXVIbN9D/OGTEd2ZCg8tPiMYV0Me8Z
ggIRe5kWKvE+hIBsDQ6TiwZCNbtxBj9DsxIMgpcsaDEZk1o0OYbIIheHUGFmxuA6lV5jd7I9skBW
nQ0iUfiz/5ukfS5HoExaYw1mCWN6ghtZ/4pTpb4ue+KXeHT2RY8wUUhyagHkPG602XL+qk4oshG0
egFHCtQcY5tVdtXRUH3TRf7kCnchgM7oylf3FffgnaHcnyw0x3/6EsPXczV5pMfAJzJwEH6zac9Z
WKCAfoEsby1DGnq0ZE2QQ2mm0GnAalF0+4bb8OGRc5AxVwzqr3px91L9ns3iaeY8jOolLz7U+ZuG
i1oa8v8fjloUs4NwjqoIg6LAcgKtv/twgn/5FJ7jp0JTbvM5R03+07Z6e0mHMmHnKHM3zKrBzAK9
U7WGNYujVOZekM7y8CGIV892Qyg8Yim4Dk4OW/5dujpP6NaNp4ewTq0a5iFmQtVKEVcW1JWrhpPR
WgwAnHMFbG1Pa/tE7imevtAsyTwlhrkeraRgdJxyWPZkamOHFdypQ8+GqAnX3XXEJmXClrx1RVHg
ogg9kSwRKDKgxDtAAdkGFdip92mMU4oYtVS0jCbhx+jboYMZEkoUdzXqQjFAChMsAwsbjXhnq4Mh
yNTq/SBC0LFrmX3DLzReOpR5z8unBd9XJvKg7wqPXARyCpiPJ2bfNWKuZ0+XaV11JbiVZ+73QBqm
+4e12DvkYBkpWPVKVIPCEMRRpqpMOPDEzrGGP+/Dzxh17+opDHUxo6HvK/MrazOZ4aD1KwenQh5U
ePAChF0e/tU7qmaCM+FPuvZUAea/ov/Fiu0WMMgaaQKeWOosmdeRexHvGKOFeiS8eLsVEx6IMS4G
gScdz3uSioMKbWZTPDmLfFwVmnGJcmubFjG9pshgB3IiBq887ufiJpzTnYpDnvCFVq3gBfAAOaR2
GWOWAR52xJyXaUcbE84feJHANUQ5EkJCyWzF0EBxwI3rfkPPbkT83x6NUfUf07ILzBOAiyMjdDfX
s4BsOdDY82QGbgidJ5LBYbmgo7+gtgRa5/XRIhu6XQTBkXEDvs3Vi7sdhbHKfPIsUalle6KSfvSu
U/g29eezn1L7sOMqdyLG+7eoLCrB5WfB/7NZtk+03+kpSAFq5V0JT0LgrdTexkXXKw+NC/nxkolI
dSEyNnrN2ARf9FQU83SZ6MhWsBPlboylzRAU8kCbwrsnkU9P2GPdKZ2lryWhSi6QkytKZxuF700B
QnECBLrRbmWQPsBQ8Gg1KAH6IiM8DoLgABtVvd25NS4eM18e8VIw2giG2xLzRtYkg2U1zi68Iq4E
smA1FyGEJ7so0mvW8CgvJPK/x0lVpiN0FuOqPmlVLjJ8Pn03C9TgBzx4N96Qq3lgWEUoLz4/vpRZ
2HG9+J8LLk6PPhxT/QeMMESw7Qnar0OpILdHYcF5ylZFh+6xPi5nQXHO8LCHF6nHzOQzUCa0ExCQ
FVXo7ll1Z4X5aQlrJ49c3hybkGffZ3iTHe4dSFx1CMXzrfY3knckV52qRR+pJ9iEIohAaFsZg0cp
+m/oDAHti8eLNqlYqdoM9++kMrDU+gneC0k1hOWzBMK6Wb0dIbRl8YXULgXcNXKKv2+okC7o9AVH
NNS4iiLleqQLuyXsAyWizgaxbJFnd8mYZ2sYol14o96bHOE7a9bzYx1uzoygmWll6FAatlF3iFTp
ba98O6c2EfbHPMJKVYH4kTEKxrLpgn8JezfxlPT6lKifD7I+myF8NzuWqDQHlSNRJjnIJPR1UsSD
UmaFZr9mfYuISDUHOMy50Nflzf5x37aTSvzfrV5zDBOflojmxBnWsGbZRqu0BzN5M8A/fHLo4R2A
2GPkkLprnP5Sl3C/ZgeYVVbpE94r49ZVhEom7RKjzsl3PK1vg0hei++WvmbnTSd2Bj5Rdak+qMom
DaZrshTppHrOk56wFS2pbgTNmJ8yvhUZHrzDY4haRbX0Yl07+9XBKIwAJHpv02bg/Rzwgrrd7xyP
izpqBfFfpAjQKjUtgssqbQ8ArlwG+5aGejbSz/bcG8/sAHbnBRRwnjBcAcq0YebO4FSNex4tuyer
1q4ziEe1oyvauRfPfI0kz0teivMgX0yeOxlC8uDUM85m+sY1H2Kc2cGjzpVbNfyC+fzpSZxRSVoG
t6wFKYevAwmg/U6WEVs1TpYA1tNNK5xjExWf6KO71MdoTbE7TVVG0XxDy7SmVv8nFAHUOiCCZ/Uy
JNcxIxlMAapZw4535t56aa0KyiNXIlf/eI1yJqNQyMq5d1j4YFrtXpSj87aVO6OUYcprz3lJt97/
3IlVgeUwos4OLAN55MiZ7zDSxQL1Z8XDJrXr+edKqILJKEwP8n6YU0t16JP+pTFcpTy3CA3pVB+7
/EF7gvOy5t5F0UqglpiXv/9cFiVNNE5XhSyz6lgUUvhiqa9uMZvX1ntnUq05idFRL+4pW/S8P+Jd
GP4gldzlUkLMHGt5RMZrJr/2Dgm2wYd3+Tn4Eq+hgH2nI2O5GL7QfUREmwrIK5Ukm4p6iGp6AjPS
3PmZqZEcuQK9ZkcKsGP/2EjeVdavCvD5+FaDeS0mxqkqsqzg3wJmxkmKPmMPmLvscXDlSoSY2xY+
MXoWsu6mBU36BcF/xoEAYZ7AnlFOhYGt8nxiMbRPdopJoEHqyGBsIrv6ur3M+ZZUULWSRsh5iyP4
9zyVVrIvxllFp2Vh12gkon4O13neNphsKo58CrV8cerp4nj90Wl1CbI8zaq9G20Z1vXCfJ4rs18f
G9wIF6+sQFcLbEq8RLPm7bR5/LWZbpZw1XE5cNT+ogZWoIJnI3wn6Uru1w8yrOk6zCz5FsAKzG9F
97aszBU5aVapVVBpwEs/9VnMJLDi/dwNe+FhgYBJfUw3IL4JjdFUuDhl74Nd5J/HUCHZwauGPGiL
eYTfywUf4UzLaV8b1Qb+bnWTXyRzMJthTpHsnQ9MFkOYqfXjiV6bYzipfbPrIPn0n1ADS4lVk+P3
6mAiuiR5NCkPca8h7r9qb+fGHm2ivdlLjLhXPii8AOR13oy/5J1XOu0qhY4ean8ByyV3Mu8YboXr
qNByovA9MPk7WN3umPzaVuu/8tvru3bNs+1ySToDM6XjFsiiuuCrkOMm0z1w3Ix0riybpXphRhss
Bnc7SG9S9evApm522u0fV4zRhpOtqZ/yJ52lThBtf+XDpOBOjCF6JnmEIEplmSsED8uDovfd5bwX
28jyb4ztcbzDLgpc8EwNi3EI6Q+ygDqyEzDwW0KgtZ7ce+OSkFfEcRJDAVnIIXgd+EFlMOuMFSLL
mtthL9kKd+0/w4eiNPa8kMqe0cmUJu1tsVnuTwJXJU6enbLqDSwVAuOxpjJo4lWD1lw5AtoJrm4g
Qpm/+uoNouzMM1tQs5aO+yXl87Gz+UNFsAPnLUaks/aj984U6InwdBEmeTjWiDvHfsuDyAV7U+6f
CJiCZOUhD0+J7O1NnzXne2neA1hArXsaW4RBHLF1B/4af+oMG1ovSrjzbp/XTKDbi6TchGy13nHr
diMZDUlyj0+hMmlA7UjwIGsjRuBoXmgtargkMFU7lgFNQRO4XsT7q+7o0OYG2ciY8s6xONJ74JRQ
76iHqdi4la1mtQqqefZ204zJcqOlELHRAP4Ub20YGQVQQ6KkxwYTQ5XdhN9VYjOT8d6w45zjZW+B
K5hnKGe1CG12JyegGi2U4+rFHq6BjjiKcZjfNaP1/9e1WeqgqSwH6s/rb1vqu2rB34qRBWnOt2nS
th+JAk04WMN9os79zE5M/r303ZlUjhsVj0RDuJsMjOv+zBVQr2F5Le5QkFDoSwu9nItoBt5aJe+y
UOK0C/1ZUqsI98FK1B1Z4TJz+DZIPewATNC09SptKZ0fdugs7+y/Mwm9cHHrfQCEIRKhIm9k+HTj
9I8du8Ky5a6ZVj/cmAw5SNd57FivHA2aJc7mg32esOQucH39ug6/ws+TYPVWWrV1xMl60SLJYvVu
aoNWrwOG+4Ee4PCsQGS/awyrYsM9RrznNb+fSLtUKmOOe7RerEvohaN+0dlcrAWDvweWBlStMFi+
rbYOKVwGVpJ0FwsT5HnzHLa82mU+d70fr8KXSrebXfKgukNyGGxJ5e2tc2d40C/MvuMJiYI6vkT8
MU5sarmhHz2rDsZgE4pncP5NlofwHwHT2chyjRTQC0gmTJ9fJ/Zf8NQ2V3OHTdOi9Ricqm1a/RYg
+6+4O17VVWVP9vfPBWyoXHK81I9Lq6MvnLuWlltZW2xSgAoC6Nnm6VewWktpzZtsjf0bLj32Xub6
SalTa0tnL5P8u7jY1LHWbuYN6TGEAwKsijNsY5HeLMGhwQ8LWQARVWcq97KgXL5uOcykIA8HB9XV
S78sHNLJa2++mCDCB6Bdj4D7nPfB6mumYwZ3Js40Tfi1HelnLD37a4VsI8nt24uECGlqdFEuX/gg
kXYsAGmUS6A9MPzu1hu0sjWuLHubOgewOoFx20LU9hcLrH/tzLof3gxQ8fe6YY1yYi4degRD3VdB
WTmAiBdklG+NODgiTxo6hdK4O4Kp+47hNTEriKc7vQen+1daPq110BO/OPrj4ezGU7IGU0+qWziK
NssSEY9KpV3j5CS0yeljXRYSUpmvi/P3ltyhCyEg2/ZYNU+WiALMtKXKE0a743exnv4XoN/G4PfA
NluXcqUvlhndsvF3MGUzDnRGemCa7qs8QOhnRoNbOrgh1HZyntExdI9sfhWekXyQa4CW91abFJm6
c/2SHjhmlq7epa4qXG625UNDoWiknZS5aZUEKFVlUyk9UsiO2jqinBGZrI2fBZ9+W1bcWXysXIac
ZuXQFRYLMQrKw9kYl5ypvsOhDJ277l3Z83BX25K3ZEx84gechr6pE3okl8z6qVX93RL4KO83/XHn
fcRQJqbpFNAhnsI330Y0sYjOlfMqICvMNS+Yim/y+yCI+8CduZInlxtn/Xg5sLR1keg7gDhduNO3
WmRRtbJgTQYzcp8xQHP3f7umgENaOjIH66Dy8kOHmjMCn17p06BVh/OXpYACrF5KPejbFwnnlMEK
rSlby/8Omig7HyGutcWaZkaht9UCKzPwWj01b93v6zksHMwjeeAX4Jj+d8nUMLKc5H1UFYzzL1Sq
+Oiz8Xl2KTvFe+z3MLP7LSxhKQtdg3rzSaU5rv2CA7oBgLkqPhrOaMQIVg9ss+EdfF2z6RwNz4CA
mqONmL4eUD81s+Pto3ULNkUFNxaTqJrYVOtLU1N4bDierFRTtRSGbqz7gxlaTCceYwt2dVB1Ib6a
nWleijUM4jKEhLB6tBnhrRWMD7+RAI9l0z+jpaUyVG7NB0wWLNX63o/3G66ULvkaEIyx7GTqpez4
no0+lMrY3z9owdT4wdlpKsjFdGrvWPxkiUfn9uNJoW7TdhEP4LIG2pcI6hES65bAP5sHZiHaRWSo
qh3VGvKjIGrvrJIZcC60MCad8iYTAAY25ZsPyw0qLdSqNkzUAd1V2cspHiw+Kt8rDKwK2RFN+i/P
UJiI913hpHjObvmvb9DREJ9t3sA/P+i0NPR4uHPlb4FibK81Gj9lFJU6h8maDfOBfgHyGkYBvt4L
uRshXo6fRrBvYoi+sOmlPDing0D376W5LEL0eqYUC/nxZs2qzUv5cwYIYgzge8d6AB+eJgUHfYSE
WLnw+cuOFGMtWUXERwgVP1BcQDPoS7OoWr1rnUiq7nD54ez35dWGOiuy+a5lsPOGHoxbJbYOgL8k
Y1g8RDcoNDgLZkuIWcafMjt6NCMNNglcT2hnP++dkbdkZaZIZyXj0JLZfyuEXLjbAhMSB/i9MW9o
Qv4HEzA4K1Y5O/itFIBvfXbxkgTwlAYQRTIFtw4kxjD6ajZAg7ZDlix48QVyaboO+GaKHFqpusUo
ZkAspi1RzTqkuNqOE9Xc/YasHqgbCu9btiibkx2PH20P/hsWrR5hqQTR9UkHfJh6TC7cbbEUgdIo
FUJ4Q8scvKA9bO9H4rGULRAK/Oq60E9Q3af6y8zVMrCOVr6AKCXffrvpqtTn5DmoiBbLgi7xsmTq
EGJB0GPSTgVuE1r6JbSaFHn4DLawJAGBjFtmZfaXiB6wqcbgDqaU2hzW6zPC+c3Q0xysr7pR1NyY
4ETpaSUDfzE0BYx40NP7OXMjY9CKymYEgPNMragz+OaqVH/PbD9c9xuGoVH/mQRzcBosUPAkEi2n
yf02C2JVmF0BqB4WvG+Gt60bLjvc6I8F81VAAvSasXsJx9ND6yh/Ukt39vX5ndSSspfJ1Hsf14JI
OTAtK9rRuQRIRPnApIYalwGJLYCFt6uMnKVNJr5+nxeEJlzF7Bkqy7dFf4eRWXDwVbjSLn4aMSLP
ZzdtLhvD8F3hQKcvFifQEwDiPz7dYw2f55SLLqwWJHgvCgT/i6gIutCYpy/OIbnd70M0Ad/3fnba
kNGQfd9rwGq/c+Q7B6Tp/Q09qLUSPamdmj+6QZzHz2ZaileqGPwQ/rqjyd8MlcmwFpUUkei8H8wl
2u1ceW2UqBfLAExRyoZuhbrgpGffhd6YiHI/gxBzZA3AIH3Z/o+ZtJVDkup+n8lBiMNwUVK9v45a
WQXAgBi4MwiHeSalp73hpYLeqZZVfUDoL01cOBUJSa3whLRdM5NaBcAERXBteY84/juc7s2i0sx6
ID7kPDnw0IQhE+Un4/D+oKMJFbcvEemqmHEvouDzGGswfONyRIaiiUxNOqjWTL6v93giAqMGuW60
snSEiRLCUbOOYI5d9j8GNrpnvGPe6SHUjpGERL9ibadzvcC5hD5vZm4TgmWlWqpArrqomvD9ubrw
5Ru3sEQjFFpxB+reeL9xuxeUnNvVcY2F2g8ZlvOS36la3kfldPtUs4kH/yKM5HkEHhQgowbbm1T/
3EJBCmZDKhlnKtRzWI9zy7oldAnNM/q8Dpc8BfMelkc8Ze8wqZEFlVd9uFKpQQaxZisAXBZdg6tF
YtsvrxKfgV0BI+7XolZp2QZ1J2+vzzYQznmwymwahWMZTk3NeGpMm4A4tsHvm0W8cknwvkZdc5hS
R8QK7nQaLztLFtTpwyV0CfaEhKAZGhFqM+b11wy4qJL77eh85y1mcTwLwpdx9QPGLUoZgZ3VS+2e
BHACmHH6KJR3+ZXbT8wQXdYwFapCV4AmKivGhFrctXBui8ZrDhcfhKquFbfwfwysZ14riG3BRueL
L1HFMb1w/Q4vxiIwOHK+25KzHU1M2jfFWBKIEG8TN+pyYT5qbXNM5A7lr9nfOKBYyJ9DNkQJxW5K
wrHdPA+pzrr6lH+VjqS9BZxRCWVgBnS+EUUdTx9AtYrPuJB+pe+tbR9ws17e6aLKHjtWKhGhYUzO
wUKRUL2zsiRdmKxmj4lQqLKn7m+mvkyhpWK9PEeSmYCzfSkM7Dk4GI9x8jBkLWWDK8zqIBuF6g81
+MjjidX3JAaf+RTWa//ZrF6pPgKiIqinE92ELzJXkue10c6k08J/2zWMYNlE0wa04M9CBZwrRb6d
5HkLD2e9EdV8H+yMdoygwVsOSiJvhEeBJAFqy05kkZ+apb/VNtxjjaQJDB75Y/QKhHbOb8CNrqU4
oFQj3gPF/TncNKpTlz6QEMYkSRYgDJvdArIfzICLLM8URgrVTEF8KfZ6Y555z4eUSyElqCfOj9cj
Z6C8gcDfHxP2R/hCwrNcaAV0sRUIt5DeBjKkkm0m3FqLblgpxUMDku2mCCdoiqRSNDejf4HUqDsC
kJa9zBDMbMEYDvUBipepgkTDfKRT5Z0Y+XqQ2lccH75J3Z0iEGwU3NwD74TB15L+UoA/FMv7lFZA
Ad3aid7Fm5XPtJ+90mFRytwbeRcjK9jqhDOvjK77X/JRA0HY/3I4nl9OwpARdHnGzzyteye8bbAD
spNebkikIVFygmThIcHX2kNt/oDpBC798Y2BvLv3PRlfK/adyh/HP0uW2K1Qv/hs9uXra90BsEJh
nybUcpFbDx1lF0bWvWg4y5XtNmgG5B70EAYOSkpIcjdiX3KqLQ1wElYDAOVdmNq45Af7m06pkkHo
1Eu3zL9Zy4KUW9iyG/dySXsroNo64bem3bprZHZGNjJD29Ds270IGcbzoWZT/AOg/wvPR1uHusLN
wIIvR5YrgAP/vHXC2BluKeGG33zU/3m+jt5SS++wbLuoThPqczQKIWmhPJrspDMJtPJTi3ihDiba
WNJum97oBe16jlizriZVpEI6ck4qzf1JHoQR9SisQ5PBp5UzKTVQlKdYUlk9Cx47FPu5Pbtq53tO
66faZDkub4/VKI95JT7Rj1gkmbWNVso6v+0tfHfw/0vj942VT3r8YIqYmeOtgHF6rDI1ZV1OFonq
0HK2OW8u3ldbvB9ZxPoUDqIL7JeJVQ/CS+ScUwjwD9eV/9go5E41yiroL32Y5x9JRmwlrPYNm2yd
AcAEYTjk8+Ns2422ar+SThpGne5yUoVfOOkDxySgFTN8WNuKjGTk4L9V5njpkM69iQipEwlHGh/D
sqYMoLQVTqqxUNL6NhvCK1wYHrgWVzHgO0WOIML/ztLa/ktBIFDOc3X6xenAJcY6E074njjf+yTx
KUFSEpIAVYZUgYIUYAXbw6Ty+QEhan6gthXYprzADn6m9Q+P1sKU8f6KAyC0WEwrNjiDApK0LO1e
Ae8bYtr3prTupA5i10nn9CqVVdSpMIm991VbiLX0Ja0mvAJZ1GZl7MyKAR9Rbv0YfhhIJhLmY5pY
57yz+fz0WGk84gwDRrcD2wDXoUTp58nzd6/1UnrEBm0+s76XRBwsDgYPl4G/BSv/JGZEgYDqKTn3
3SIqTnj0xfK/xuTBo7kfh/1sTk0c3cNWhquy35FkGxLdznTC/GwH+yfYlQoJQN15wBciSNgdIrSC
j6pOVASa41Ffah+NqdXXaxMFkLrWT3wjhqKG+BbNvwFNjHtAYliv7Jg4zKqmpo/xdRah4x+c3yiR
BR9vVguxl38iBp6+vynG8pj+sKXCxoSglzIe8AftADPtGHz+thuLssxknHHZlkoMEtWYmRGc9vaN
kFKrCixueBer1CK26CT4owrTW37lYovx9E/OQ3gk2/IgTM/2XsUOkNa9Q/FqZIJ8MfDbH5xbQlCc
lQkn2pA+9EqBeIduFiOFYMu2gj8groKfHXiQ1iB4fHPSrmMa0qRXWXcBXUnq5mAtWKEJV6IWXa8S
r1ubgU547CPrVFGW8cr6SP7R2T7WElsBCiZNV+C6v2eSWomK+eD8VWoJ60EfWaqto7F0epr3Ay1L
5Gy6iLj+exnwtPGxxk22LpN5895pnWzzcJNjuTXUwP5u/HdOldPTdhZ74sr9YZMglvFIbGYOa1NO
0lb/QKlURJ1ZpDUrpk/qc+uCMvlzH5nhBa/Uf8LiGWLKk9V/poZkf+CYzshmCR8RcLq/fuMHkWbI
YO5d2SOmdU+uU4qnhUgK46eDcrAlYfqrm8LFwzm9UYAcIrNPo6QQzkd0fuTKXP2DqKMfgG5s59qH
o4vsh3XFNIGG4KUalxe6Dlq2RfPof2RXX/hImSdk85KaCbadUc3K1xiASmhrjy+77akXlAiKy4iQ
T7+NJgy0FbAC4iXSadtRp+iYVNKJP2QjcjPsGzsR9XfWS6v5uo1ANwgPDHdL2JEPinuRotfDlhiA
ZKMAfSt7D/iCy8zGRKmPsKkDdTTHHPg1o4jOJTddo3mdutZrNIwxqTzQAdSzZLC8TG+7cFJ+99f6
IQoPxM/uSJnEhMcAlX0YoGrKsntV8F5FjjX3B7AG52ahOgnGYv7SiAMNkzEFjbSUZ59/Ml+dVSiw
6tXpyY9/r+5LFySO+iH9miif40akPGempdGo4oP4OYPEp25Js0/CWoGfauttz5cAH5uVi/HQxbfV
PbP64X0DZsyMAQ6dtfdh7oojh+OomNlhDHtp2bbIbNhHUhsI0dDB0vHAmvcTNZqB/t6KMtqbVe8u
5aIiW4/HnnlaeXduyY9HFERG5eLRvYkC7dTvgd6lRNsx6QvLmfi6lUJrWyzN+b+pfrQA84hHwUHS
swb+eIFp2JwjthfUy+U9491JkJ3PEWGELDVJuQ/MfeROCDzFckXmfY0wBkKDoiGGrnoDLSmiQkSk
CNsj7sdXX8gKkVBrrsULrGXqhcp1MQCnUQF/oTxieaxyEWxWDfbwRh0yeanwkSfy5DDmtc1YrkpM
gZhtSqm9v1VacErnvJ6Y5EK3n9WwgaiNRpYYQOdUKBrNx3IrnUOfFfo0Dfq3eS2YXCLgyHHZIBu3
EOMjluoPVj9II5MsVPcDQ6P+Gv/dvznNqvogeeNdZgWsqFj4HBYb/7g6l7RZoN24tQsCbaW//YVi
2VqEa8EWr3reVp17unqdGG6/JPvg1WRetaFcsp7wKcXgzdRDgOsxN7LhgjU4VkjrNQe/KDe9Qc/w
Sg7C12iyikS4l2rjfYCy4LfRA1n1TXpEYhNNhtnFog1LG2rFQ/rr6K5xkEMpWRycwwtgPC7ZhC2K
79wZ5BMn1EhII/ugUnNAnM7nZ30fQNwawzMZZF8+hSyOrk6UrcfwvjEj9B/0MEVqRAG3O+pJ/ynm
GRrUqGbH/5ItJuvEmQZcqW4aAMEXQI+Amz2QbmNiPqTkRVjsQek69Roq/bny2nKlf4t7AdQfej/4
7bLXuUBRKqL7bOZtpR3XlZi1Jmoy/rH8h8p5p5zrA+u9W/4W2VwfPj1J5plPt0JU5h2mTuQ7dpSr
1NjqSP+1s1mwizltYsB4OVxOJBRzjl+18Y75BdHdaFMb1dvQf5aEfhbp1I4tCkL20eWXLs0Lie8L
Jt8+8i9VHCeX11ry4zkNcWeabfqGUPhMZ5E4eS+KOkIfU1xCOIUM+8NJrlKGq0y4Cv9ew0ncP55+
cqh5khDGVl65hYSwgOeLAuHfxDcIqePjt24+I20zKqyKugnLc1ix24/fRX2WywItVnhT0W6iHtyk
u4fy5fuPZwPHpox5fgeb/8JwaaN4oYNfv4H3buTi3XhvrGXpsnGm04uXqXoQDf0RmH3yu8Wnvxz8
Qw54nwr+KoegcUUzvqIKQCK3pUP80mF/YHJxcEpGmRkDEdeWULS9QbPUsUmKC7ftO/ppHDqXRv5M
JB4TohRkGRVvNI7aKOisSDlMDS7k/AQFn+fH9w2pnKmI5v6PiAF1wFIk9j4sMuwlDqGSXPj1zf0B
3fsvksJRnAxX3D9aEh4s0zi+Xh3N25YFSo140RC2n+fEaHh8JZ/kmtlZw7HKOBnCx92jEh0qJoej
4vbSsY99ato+R8Zw6v8Y3/oJWD73Qh6gY+OdWLRtLg12SNPWJU8lvq965H/HdxJL0/J4/11BZTVQ
vjvkjel/r2HSkFPSk6PQ1xjyFklDTOPN/0tCEPORuiRphSUniTCAXO+W6/zDfJvxbyNIA6ogO7WK
VT0g6e4x++46m8WBprhfIQuYGCoNwhhgz35P4gl0Ol/VaAGVXP/AI3SxCQGb8U2VADxs/0HOvJpf
hDeCdZmuBTf6TwLzypYbUphvtsYighW2wV4cdAv0gpze8Qphr+5mowfnEZZ4uUN+VDXCkFQpDftK
7f8Smogugbni22MYA0e4N/4/kI5KW0vHBgZgHD+Ih+UbA9haUp/hdXvxEO6xqRHuN3ZPKCrbOCjW
eynN149Zpx0d6NNQRBBzIRuL3ShqIZpEnSVU5eJkPAmVNK7yAi/oLSY2fsRDo9esqfIaBSvItLpy
YbnbtPXH6Z6fZ0hwIZGuISmTjWzhKNJswqfvZMX+l6hVt2JZE57tbQXMrSiRHxtMnpcXkikoV9U1
qENUpFYIMH/Ew4PeR8/itFNj19dRdP1rt1Gv/PL2zZf9q4jiHAGSJgtUmhR5jKA2dGuz3d7cvNon
N/WJqgSPPVhzrnKpH/LMCEyvbE3Nl3maJNNlNzG/cq7QEBTjkL3Slp1I1Qdnh4SwzWWqhuM+rVkk
ms813NibUlNkUh9w0WUSI4/g4EFcB0AbyemzoKuEQW/P4pX8FsGNPO6zp4bnTp6BgCCLhiOpbJ7r
P/8OW9+Y6R9RGbDYOe35DflnHa4YgsCJ4n7su28oXtJ8wfcOrcvtI5fxLW59ctPC34lVTzB9x/jL
alEkx0dkgNDxQyZl3dC5Aizc5RrrD0qRCJJmduYMzao2SIpkKR7qgfQ+P4i1Jj96UbnHfv4RmCmd
Ii557ZF50loaSXm4JGLXF/nyCcZhMIC4sg4qJAxKICf4bWUCL90na7TWwcXLRJZ/E9zB6K/CKVxK
20LcoB0Wy61jGcCI3SptpR2PjIQPedUI5cEPF/py13mteYSjdquJKTV5Uo3eZFBoZa90CrCV4Tuv
Mz/E+oFeUcMpab/EjvLgEeyoDRWLrq3yjpYspDvTV3urfgw7W57+v6PGRzpdALnJhtRuDzowMFgm
ibeJSSZQPs1Dm0B34VGe+DpFxtSTiON/GwCvj8aPZocJyaOkRAV+93mvS8h5ZlcLwUs9gu368gSt
MzzyhawBaBhvOgTcWMWxZYXNLSttT7m9YKHz+TBXsbQ58EG86fuwGY65OWOXxTZFT+Ky+bEz75nk
b224gskcyjDKE0eJ0/ukzVFmTURh1lgslc0hg041/cwUACxG5+pSkczAkrjjv/1LF+K3kdspuWwD
+NHX5dUWeSpPA19+Yk/EtSEEJTKAdCjn9vJuQlf09lBWTgVB1bVsOCNa0BgoHzGK3OTpkj19hv5l
3ybG/FrC3/dEW+xXE6D7ujhGofEBfTmg9YBnKYTDZwa77HdLTGCsZXyvNI8NbKtCs2DWHPqWDs8U
PL64kICEgv2lwYlSDXef+wi+CrEHHqt2PbcAfLRAr58M/ltu+xcDbbDqVSVvsr46eiFhktJt7MES
l13QRKBflrbmgM+0bl2BF9tLR4IB+6lz5iIPS4qzLneJ0nAVe474S06IoKuTUnlUMyWijf9nqx2X
mSxWepzy7xieWZ0Hw/Z6EQtioVHemJnkQw2XOFozcj1LFVsdxzjoP/MQGLKNydik6xqGEtsxEsD1
UUMP3oW53HAUZvz6ot6nKZo5w2f+xrKB+4jMjbglRg63OallWmClOsmvEVDMQMvO75nTH3yX0KXY
X8h+kZshrJwi92VEAriHkbSNJXPQUCQ9Be6f5EOadpzA4uruZvAC2LMcvXGYSAhHttDdznDAEcyG
Lym5xVb11zZWzNlMt9bClEn0vza8VZHv58tcjM6/Q2/mMfrpszGBl+aZgLfQZsCD1ZcRY6QuZTTP
Oc+AnlSaOxBLvaleWoT19jvjTFU0XHesIpGyJ916qdSiexOsmK8Kh4ENDuEYPcZ72JyCqqclUZV/
Q0q3lcYrQK6E6abbsiK5CiGKLakeQr9CTId3zTXxd2EDLDt9c845ecSyO3OJkG/r2gX9VySLpTay
o13hw2VeGRKz/WgYTYkYt5l8bWud2okUHyd4C0KZWbIVxB8Dn6pWEcZQfVZkEKDr4R+kEpJZpbhj
qNugdVBYz4+9ab/iJD46NuYtcsoTnauvt7Vcym/GSr1HRqEom+f62id5XL65YHfaGwNPiSJihXOT
5/Ey3VMakQLwmUiFfI4unh8YE0CYm14uDTqXQyoKktADXVm6Vc3bUprb/fTu8WSJoPsKmZamA0Bv
3hQk7Tzmr3HvRB8uK9/+aEHQu8mwuZCkHRSxoioYn7wZwyNyIEGi3mZCUF82GZjUwQn6mNRErDbF
zsrUlM4WfjaAhMOJOeW8eeCrSdKliC9zQNoKfX0AmyGuyTuO6mtoxAmhYX19RXXTi9Q0F7BABUq7
kxwRG6g40lbAYxmQ2kBpYsXWvV7v4SDvDYQPC4AEWN1UUeZoCWHFlorv0XjKj3/CYgYi3O93AH3+
LbAUzzfZa+x567ZAzHyLAwqPZZIY+sh+3T8OtUyg7/l+GNcLTjboOlACEq24MAb0HIGHc541Q78H
0F1B95LyeMn7NDPq0pIqrmve5q0WdjY4ytl/7L3fmItjLO8zu0aGyE1oeeZ+nkZP+pHpbeQeYJE6
v0tQW00BwswSxUjXVOgl2yZxyQZwbiiVfvYhvHtFqa0vOwXpj3IUiYG1oG557gsb75UohB3Zn551
9eWDZ2AK5dXXd5szBZNVwn/tjj3TxrD8Otyal+qRY7CDaKr0AsJJsjkO7L2Oh4gm73wU1wSwfrSW
JjrrqfpjXj1u7cGKOvEnMnQUvTch8YP0TT/HcBWkWMnjQKrme57PZaQ96/ezRWz3pjknTGHBALc+
DlaJO497w0W7kB5lZ/OOS21JA4VWgAgTD2Q1gf10930pM6sFTPHHP9tE/QOtxOne3nsDRfVDXBba
FeNVWbQx9dX+HIG+iko3/4Wn/RwYDBIZCbRJURCmxwRFaCIK+iS9j9uiFLmdSvCkOAJR7MnubF5D
itasnF6I3vo//bIg++knALus0X+KzvSSU8wS2COHNuqJUFr7EQ5n6kczdM6z+X5l2z3OOauK6eHZ
jbH2TOwt/vyyoyP80f0cWuGD2jsFfymw54b/wdWF5V2FXPsKthzhM2vjWxmTO5LLP+f1ES+pKIFZ
zNMq/oFs+hVrXSZtrHQLczx9PVqTqsf5TQ1Z+y4ssdHr2CCANSwkOj6da5BAAj55qQCKnjBeBQmu
bGZEb8OLJBb/FTx5BqQytvZiI4oDROl7kUYCf0PI1FXyneQzlNi/gOvMGWyAxUiYSFqmv1rgTQvy
/WMxmiPH8sZikAJJGrhySn+8AtVmY3+OOjpbQ1B7bdcchSMi/38/0k1AzhwA5zIX0m9V7DRAeQ8R
wESvH6dUcajiGdW0ucokE1ImB/AjusYzD9ozKAkKHe4X/tVguLOMWpqRvfLHZ41C7bn83Bgc5gfM
+/VSNGx/yO1zGBTJB7jCXHp9lFjn9WRj3ZX+CHOuwO0y0jgk9YQLfx+5cl5S4Y5nX+awMWR8egOQ
3BLFt5JL6zKrKhEsEBeHz1UG8ldc80+g61VWy47fPGiN+FqjrXEAKg05K9SB8/zMG3ARhF6igXFE
RW7fZ4UnsEfNQLeM8k4d7keVL+uf/kipGpXZG0oRge9AecGCiMiNBufos6mWZ3S367zX0IhNBI5z
S6v7wqVAFhI1Xhysoj98OmhAG2jN6O9DUfrCpVT85ISEHhBdLdL6RRgamgLPdTARip+fFNtRhkHG
HmcUn15bxYeToAa76/GA1gDUEYLvdx0fCwtLMWtihkrCoZrFw3yy8Fnw/YcPdRpi8MrBrADK2TUE
ZFbyVmBxl6RhSXlT9UjzAMbRQawqa/39sf+wmdeV8e0uiqffJV4mTPKnVsB6yRV7L4V5dDSZ1aTP
AZ8rMeAKZM53YUKHKcrJsAdmvLHIMyfVdwlueKmh5PRuKGvcDmbEV+3+YIyN6xu8zOVS+MJBySJD
a1U/5yqMjzRwcg6/ODtZoo3tCLu1bXIFaa/ZycKQCVHTsXEYv0hK5U2HzUfnhgnyI+K3h9Z/KOJ4
aP0mYcoXNyTOn1m3cV43S8JcRw9sjOA2ErpQhqWx6IQ3sNWfRcRCHogFMeD7Jx0mpkMN/oKnlo0z
URWQsSrzWAUO34XX1eK25mxQea1EevKJYQ2H/9U7qKGikG/ghk0u0t8gBZVmuS6bUGK6DfwE1NHA
iouQ0NwqMwQ7PWat6Y01lD842Fk5oIKZq/skPkNjgSMEef7DvoE9sTxBXMHdae2hDWuP8FewNdpc
Ohfc+B7nQJxJld0m/fK+Ff6+Ptext+dDKwZRqxSLq5sVYdk8rss9y5mPSLFijhwKDKcLkRFAJ19A
ootyRnMKGooLTiCkbOshaErBIQWEXm+KezCIKn4X+xrAfoh6GccJbDJP5Ys4gxDpWM+3RpF4c7wq
2ZPFtXjrKO3ZBPP4pkEjSXQLaES27061YjUhIOCkBke2hvIdTAoGVKkIOiGnPNtZIYrtJjyklPG9
7whM2ExcyoWPA7aLZ65AysNQqFBOKuCm4iI8UpHp2qW7nHgBZqaLVj3K9iIX0ppxBCuwCxB9A5bX
HWz61/0Wz0YqZrTUzJ+0VN/gT4GcydDK6j6nhIzd1WTlf6s6sjP7mW4VxKlqWXiMykFoF+gTNGKc
QItPKVdxWd50w+eQomOZ3BjT7D8zpeO+WmBEHfx9EU3ZMW6Nihyk61E8/ZraIKAm5PNvhc9AkSm6
KJyjCZRHa6Hld051Ix/na65PKW84atv3wClpdSwUPgcNcWB9swC8UEQuCQuJzgUMTEMw816pFjSN
N0oRhl8t/O106IzTElvhVZ/byAHcPIV+85Pmy1ogX3c+bWa1NKFGYkgwEIGwhSZLkvsTZq0Jrfma
ZzhICo/1YuRLL92pp/nHDIP8ieBVEKGkg05zfqFeQHFVfPZA9aPRHqOV0xW1043UxamIKdydctg9
KBv94ue/OwFKhKxLWYrg4s5KUfezPg3sbnWtUsnzzr7lN+zW3tzSL9c0kksLdbcSs81qSIGTeuAt
LvzjeMDxd01v62CzTYnmdaLGIj9ilmW2Vx1rj/4ZRickzXwZvfXAceIT5UKHPki95W/Pf1ZzOn6L
Ck+rhqYRxUIxSJA7mpjndZk6/eg7rv/TVNep/qT5s4BcxhoaZGocX5WY00LlhQ1Pw2jn9R2Sj3Js
RryhJD7RcivtgLs9q0D8VmCc+gCaegNfs3TFcWJfW7dXVny681j9pC8oXDGTQ6IRl7KOWfzACHkn
f01JcQv8q0INyLNb90pkcYSu7VCQrm/4+5PYVuNFiSaC1vBel2cv/wgcqcH085BHNrohlUJGxqyN
30gEEMX7IuvSIeOTDFL1ysDl01i4I5s7RBDyuWuLE0x9bm29hWBaOKHFBU2tX/JWFUN3x+kUQkHN
XJV8nkmIUqlzXJCpXxm1es5TvWSvxLqMafEPapAgEsFieZS2Dk5oTg87F7PsNHT2oFZn913KV29O
NCRJWxMLyykqEtQfZBqoDGl7SweA4bAojd7OKFECcVxaSr6sg7WyU58LrZ8pVosE56HtbkRLex0j
gA77geO8sf+ivFZRQ1x2wZqM04x6Wcnk1j3rmmH/CJgv6xTBsp4D12G/e2YN0BO3ZYmOVQ+z9vOc
/4+g9OA4287CsFg/TDrmVe29vcybwcQUjSs7YVsHRUUi2p/cKXeJAkJ++NVOVaj2aObtFtccRfYS
MZelA1pPKHD9WK8ENN7UlmOapHbibvZBsZnZq6+zZSQeU2B2pt+Lqwis29h/8WYpG2moesZjGj38
aVzRhLhTK6EXSt9Yf9gadHdCoSncYvnl3meL+cas2bQO6EhoUsf/4/eYDhHgnGRR8EItW8kXiMXz
ukBqN6PLU/m0Ka4XrlDrOBpdirZI27ze1zdrCQVWOfmVyZer8Ms2+j9uw8XmuVdyb1OcfpXmoxvG
UtHKQyCp9v7g+gYrUGMiIlYsoTixYf/QnLEcqJDTOmjGuKfXNOFJAzLJ6INbAeWL/PfSvCkT0zp6
AOyukEqlbypjSXQNdfEkW1neY/JvoKMTAem98IamBr0iaPoGVFBiwWFLHcotmMN+dH9r06SzSpt5
j/JEns6EaG4OwstW/6FvUmr0PygqUsMLCZh0ke1wN4SN6hSQzm9UDJCtDDrU0jC2z8rKn7znkU+e
0daQyD1p0g4KI7iDKK3nBQoTRNjJ9QR06l8C880ZoHK6RioBjdR2w+L6I8pVYTuq56MqZTjlflKO
Z7l8Pm6PzVeeWAnmBMYbaDr/AE+PARK7gIGWwCmUKofdtdHRKJ5M99lJNgmhUMjNLfqL8fsM8VdA
NDIzF5tx5Hw9/F+N0tWH17gvWMi5FV4D0SIbP6brBRTONE4x2gcDKs2sBMQWvNiOGqW73CWYdG8R
llWyn4VNFZ8Hj2ctemxav4d4UuWnrojCptAy47b/xqgdxn1aQ4i9HGrwywQPFlWdm7i37kl14fwn
QJskILvYbPiOqzpdRWOvdWDyT88AwVk2gZjHU52E+B0T+ohyCpGdkXVE5mXxhb7TpjpBfLTISzYK
kxX+/WYwIEzMPujm1Comax3o2juV+kNIoS4FFEQmCD4sycpsLK8tk2r9gkHlSGiqW+afVj/DZDO/
c3iIjN5sOfj7165iEmqfbaKxwPCErJsThIkIHaRq8Gnk6VtX5jdgc0q7BYHgJc3havyI7sGTX54r
clxg8uioQozWttXbAF7uD+i7SRJjrIcmgECsh8tx07lSyb700lGqmcjzKHTWGRDZ18PKP8JpraSv
L/5TNQmXDQCli97fj4iftKSHTJ1KUYCLE8auhFwBIM5bsngn3i4HXl115S2tr2qLaF47llOEdCH+
lDW0/jdp8/RmsRqSJpj+UeA+T8ZgM6SMe4to4pJoaEDmkXSoIYllZCxbLid7j9iF+stUifZQRdTr
etWVWDpRzjpPDbvtMvFf1VaSajJleTFd9PyKn44wE5roL92IrQ7btcKSLSr+emKhx5VSlbFnkbA7
zMamdqumT2wyZckZjgsocKVl5EhBeVnRJ1VXSYNGu6shdY81BAagSbrR8KkcTj2CcfkaRdYYL00A
4hTzQAs5isObaGdgjqjc/dcZfNMKjesT092RvvmRR1Bi1ix8dyeAMCgF/4jNXQFq7OXh2hesReUK
2rqp8ekiiXLBogi2zAvHHE/uCx69EkBb2V0HZo6prO/0790PTNOKmACzUJLxUYsk+DsNU6d+Nw/D
BLMcuaFcotfdTNcCVJ08dKpVu7r58RRcKcujxUTgsKT+MlRSXm1jV+N6RQqJrTmsgOQHaOt4d6PB
R8Akdc+AuP6dhemnLk+0M2lR0+iaA7wL0dLpj+HMIpX7pSQFZ6G2jhJoumrhx6KWvkCyj+Haba1l
YG74K/mhI0iVi+eov7LxZl7NNA/0kx7Zy9xo+Kt+DVjO3A6J6sGTvkUTKczpLjLi60T2i4fe1jtz
WP7tjPJzXojy85uk8mrdjKGzsRqf9AyQIM+u752C0CDxRl2Ntnd4eSJT1ZyOUhcFyU8YXUZvAQAh
QPFUyQu3397IbIiaC0fgYHuIErVaczWaZzZRGH80lKD1aIhRUldmGsdpWlNOCJfJv6cHL2hkAL/y
IWRpeEIOFpkwntRl2Hno8sndAoZDuS9WvQM0xocjOaPPEadRp8ZLdJEoWbvDDp5Hb9+ivWZ/gf0r
xjL0G80XlDBKd7ds77yE4/nNBQbd649CyYIl/fRv/JjSPXXFvZTFjUMGID+bWwrED9xN73N5IpQL
TAq4kDwXV3yOYifdblq7T424KXPo1a1s0KLf2TDBrwkGAR8OmXTM/1sF7k//kYpjPJx/ThwuKSPl
iIwDewPeZWq3yT5wmWScOpCxZExA6EpExmAkDVRhcc2t22DpD41MmgjBHff8Axgp5zYITmqS6PPm
IfRXUti5Sz2EC82G23Kq0n5zxrKqiCnvi5WMSeyn3NBCsW20KM7/2rCd0/En4LlNS/ljlAuPJzA9
Rn+cPeWTTAvWoDekFcPzz+zl6BfDdQvPZbnGdZ01U81y9KMeGq3OYrLlw/rl1lNP6Eg2Hk+ZIlMd
+BYZqlbUY8LMoqydyoiT3aWRULlAWE7DZeXnWwWYwMg7MmGmDFqIU1Q1vPtyqHxNCBRT91XzA+p4
yYYPy65KJ/KBsgVgNDoCMJM1fLoVnVZCLmm+M3rWYantnKSjYOhOwPXUV245zkObRYAgbFx5UcLR
c6KWKb15OynyIosYZCgDuN7SrvwwM4aMXYyLePCdJdj4mzxIPR9e3G4BeIeuzTo7hCEMIvCVlAn3
EMPvrx+ghzrNxuD7i9LN3dl+Qi4tBd8xWnz39krLcFxZwmcnyAl4Ut2jk2RRv0aT3XulzE/c6GZo
ugXCmnSXexwcYSvw57RU0CbkRgkQ2po1IRsZ78No+kk5BFoSB7+llCNy1UqWn37kEHR/XPn1fwLW
tHoVM7LP5uwnu4eoi47j8tvCb44buy/598LTy6sTntd72PXxXsxXgA+KnttMm0yY5UgoyhKY8Dct
3lmQAXo/VzKsPA31ebYXag59X8VUGlZ+n3NT6eLPdLP1J14p2s+OXA9WsOvBEaYZXuyEtO6/HhXD
RrDHuu4AMWnk6aV6EdsU2GqUnAPFDieQ2YcRcCuYPYDgYETMEm7eqLI8zELyElf2A9TrUU5kNBcu
p/NbfYgqH3/UY70Eh0Hv8Fnr87VBguN5viSet50fr55SM3VpaEdhPxODPYK9i2kKeN7jK6m9Dryg
UplX4ZTG20xl9dLf6TgsL+BkE73S+UEUAJ7w56KtYW5Ofb/WY4aOxHrkOOTa3/20IzMd9oUZzD7G
x1FwyMxFmxVIPfcUVcfga8iIVNSXHOnDthxmIl4SI0AGXP03CdCMhnQy2bxx4b4ErDE0vhNLBdjW
Vcogxi9gL00IHuL+C0zIGC7ibK5OL7o2mwNa3bYF2dIkEQT1w0hAR/ECXAvmeQnh7rFzAhKFuMZx
xstG+EnvWxheXR45Be+406b5IhxGHW2hXW4Im4OHXVc4AIEtOHroCkENsYrK7/n4X7X2G+Z9G218
+QRmCveK61K2UOnLme1eru1nUqbBoV2jOzSm5FCZZXX1ZtryG7B8jt9F+iapKeN9UG9Fzdi0UGHG
fEnefqhC9uxsuuErkhhd3oBSVw+7tlUoHk7TauSOrRJaXsunF09fNAEJDcqNSzd6QT3xvK7LxwPz
jA7hVipbraam2LZiu2bJIH8hVmApP7BDs9azqWgnTLFo/XeAOfte+e+THZTZWFwmfuugdiudeWGd
65QCBDuXobBy8SnRIeiTm2/X50XN6UQ5eN6/1NwEWvh8JpxTM9zVQPAc2S+fBORMdh7ewy84+1pw
BcyT9DgRl72q70pMRxLD43X6XjZPFqEymi6WMvPYLvoxqVfWAVaZ8Utx2xXFCcvdFbPLVn8tDT+s
DToU5UQvTNc2yNz70ySZyEQXq4unI3TRYj9k6WaGvO3iaTJWz8eo1zc2782f0cz2MpOBzHBiIhnH
AyVwt2LQBgc5tSmGaHSfCI9lQl0xALp6hrMOp2ijlJ6sfnogQjCFhuH8OL8XOchROBpa3xH9vLJz
QRePA8IvH5j8ZhqyR1g8+bEgNfrctjkhW1N8HHDw389WePuT97ttlU35cjyKaFyFZGUxLep4nZch
WCAx+7rZCLTBO1I3CzSsLVquNA5Awo7wiOdEKcVljrGDUSZpJ+y4UTkZP2hKow/benL+th31Hjf9
0856/+9PfRtexdiX7I2D/SeUfKUnwkbU9+HTYQcPJXfjdfq2gAYGL3E/gsTfdQ5x8E0TE10R1rx5
q2ssuNW0N4pugHteWPI+eM1IZEBWIXctlihFeQh37uhcbMQPE9tPCk6xt67A1SvQsEJ/+EXyykdd
xj9Nh9aM/kAgca1vlq3IC8LWVTBBn28/cnNG92i2+GhDh0wgRwMTwzUG/WonuTklmDCt5KcqI+93
c+md8Pt3NeD8b5xLlGSOTbOOHyjK9aZ5uA+h2PCSrVIJdOfyenwBdmw000/jt3WzMb5m9gPKrDDG
hWY28cIhXiqeqXs/GA6SPrcxiq5zz3x1muSp5tRkKUAseaCXb7XdMqyFzQGbvLjn9bE5trjb0jYX
RXcgGzs2KN7T02/Hpyy1mLsOzv0gDdQkUzdIKGv4M33DAgscOnvf2rD7VrL99QmrvEKqUaftoAN/
4zs3GCOi3ojU1FCZUAdr/NJ7sBSo7PlQDXjn9wCePwA4H64C28wvkVHAJm91fpgklLe7QvNAjwPL
SHQouFZgmYvqvpXX9HVOb3s3RUMpjukHE6fU4s1Q2x+N2haR+helAX6yxcrNQa7ODMP27RfN4460
GCASohTqdFZDMC2t/mDuAtdJHMfJtTsK3IiL+2DnpCOjsowRqtXnY7qhooFphNuLtReE2bqU6n+t
Y60V54cjG7I93gXIgHM01CAXUsXXogqRwHF8GUcQ6rW768qhqwSRdaxi13XQciI6UcrXzfuLiQRH
CZho5EK6wypn+/oRmbKa5fcDx5jCIag8W2X0Zj1fJ79XdIKllyOcUmj9AUkwkRvTXde24rUAV0sR
10YGL5gjA2NAV0VfO9HwnvJknBmi1l4pVwo4bEzCCkHIAXb3CksmCUqh45g2Rcwh54jRYrXThHPy
g7WFHaNqUTePi3gt/l+XpVyrPeSwrcTWmSWcvybq1vGR3mOLjvpqdtMfj+6JWXCqhVQx7Ak5T3Oj
eoDmQ+OitQ7Ugp4oeGrgTpbLIo64NX/hwyIMgvJHQtqr+BXSdlzb4siQzm5pgd3NEsZjorJOMFWG
0PHTOp2MXZr66kOa40X4V37+agpmF43bSbjF3P5BKaSvI3ks0m4Q4JLKSEwZ3jQL90cNlMeaCcrr
d2mB9QtoRUh6UTmlPDyzQUoObdnxHvyUUlw/fg6iQJIbMdEmwaF/UWqKmH8B7iZasHrJhTDBWVlb
tT/1qYfWAWvBOsdCXBIVbhCX+AjZVxQZhutYrL9CT2ytVanMh7ZaQX2po4I7aK5gZHqcDixH6eNg
qNL6vfBbNi9/wvLdhcFarv1ULSVvCOUenLErxarY4rG1+GdnKmk+vPZl9QR6x66tVPeBlDpYDF0I
FSjODVr9DV4jTIyWHtDJ/u1xPpGhpWlJCNSk7NJZVM2LgTPQ3khZsd9nWMypE9wcEoUvZY8AXXnJ
/UnfS5LfJdhrxIcAMI59tOuhGYIBey7Do552r5DKwHK4oNAchpsyyPd0z6cxHOl5V3IRAYngr9zo
fevMbkWsGEDEjkuCcfwlSzV1a/5Tboy5cXmm4zhHMy4jeDLZx3Ap6bzmtjv4jWdRo5nBLli3d90N
m3SVDc0uEeWpD10NrcTjVOkcmg4aiWe0zVAqBqHMmOg0Pj/4g5cCyfWlnsCEv403c22Ub49AnpQn
R3SzvECng70L+vwckaSyD7bBGl4J/LC65xCmG+1z5OiBP4QAMe3GSZBGoMSPS2hQooZVviLjf4CM
VE+2zHyqgg0Sh9bcNVWv8r42q2Ipmy+6Ag3ctFdN1SwEXvyQ3tdYYpJKZ5JPbk2IKpUJ9K8+SGS4
WOBIsQkSX850xo49KD1R5lVFTDaxMpmA5LpdoYxWNWuz8KLi+Y3qQTfo6Ez9N2Ep8pj1SLw+RmK+
XYC9XKw+Zd96qMgw8EEk8mDIG809p9K32NtXJr3s2grN12DYQtihbrZIP4WmtICN4/LYoWKHkAv/
25obkm6L3uFtuSg7gSry3G290tSFevBUpT/4OnryuE7aMEBjOiXuJwbmW9bsiCZBLe5IQbGjItAC
Hf/RV7vRSxWvLOp5d4WQNCWv/NIZdxMj0yF87m0wN2rgmbvb5FSeAZGqGqeEjU2o1gp2Fl5d3z7x
29qQtLjD5PjjbhvjkpzGLt1C7wC37TcKabi3P2n2dGZvAabWaTQgzEmEaioaA8wsMvHGoacJv00z
h69etzzGHpZiK5NiHrZe4aCizTCUuVGTKDtT64iw4BmC1ifTPfzIDxLs0aWfnDL2DjSYsnUxNfPh
+bzp7fmF7ROkYNZ+WIW2pIorDbArU58JXmnJhMNhctFk9OzGnNCW8JTdE1R91zUz/504+2qoams7
ccKErcW5W4IgsUyPOPXr6LR05mnaPTftMS2vVfwVNEp/VlIPjFQehSydOnaZSx4WCq94l05jlEYs
0uWnbfKf/lDvq+8x0booIgqvXNZvT8sPVvv3+qtlC6+aO/BvcHTJIMTfYVIHgirE1xhmBs3yCtdy
SWbH0dKZNm3yCi5pjwqjLhc3kxhJhfUhALUw6sDDqEtdQsIoasX7WeMLOXmwB23e94OXiSNb2OTB
6hAgn/G1N1ArFstUnidkkc2nSKx0heSBwaar7lt6SaX/yWW+XxavetUTgX4yrJKcFJeElkrMe0/x
evmVCuDMJe+Al86/xmJA8XSO0zuN3Vj4jBFc0G5IsZ/lZUYCqmwNg2pvUPt/V1BJ88eaCOX6vX4J
KZGsgpKvs5keSh0gLP253pI6lV9AJHnqyt8Jhjp+Ng465vY4W2lyWJW7LWbEBBBCPLnC/2DLWLZd
TGLAUqMkqm9l2XPUt3bEHaIx86NeC+1dpu2hT/8hSs6HjqtbvkaXt4kK+FA0zP+8heCH8njoybZt
rpxrRiSd8xrb8wHvPPmm+JVuT+9sFy8eHfnvMvtyLEzlaRcrEjHDDIdGfFD3j2S2wEpU4dN1uaOw
Mp32SZOPsOcDBt3xP2ei+zknlD7C+w1cmlQyzYC9DAplBkBvt6dRCitSllC5d2CILFGbR2O9yNZz
SKgwluoQouVsglZDwr1h5jtFRspN8Y+Orr6QFEJvDBVUqLAtbNIHc1LoOzjG6loK4jdySo3Ooi0C
8zg/apLxJGz/yAyAV5j6kZO7BAKiNUzbIxcoem2BlOpJLdXbPC7BeGutshwEG8rh+sKTyyyJuXnv
VPNn4JRnhL0zkFdCOTCkziYJZ0JmwnygbvkeKVfumLyJqBY1g7O0dyES0olVp9rYbzjD4BogkbiT
rG4uF2FgM5Py5Sb07ewK3TEnDkYkVNx1t3bqDc6lgaCzKFqS/7ZrpR0TLYbbasRo7mxwkRI+S6Wh
4zL0w/I2A7wHJnjBkfqVOeva/reVXgQ7jzCi6lN6sZYLzmgWfPH2D7g4c1EPn2Yjbx4xVhengfAG
b+TYBrlEi/mPhI72avmzqrGWxyvajhbTI1RIv+bDwdUA3UB2H7MyfdXIA5HEK8bqmfOjC5dszqlG
kBuB1rXKvEYCPsv/SODe0oW7DaQwk5i84D/GCqRsrepeL6t1DSO/Kg8GwGp1XSQaBw7rti0KQ6Yp
XETIivtiFq1h3ROuRLcI/brYI8QEXNZXlArJSbolVheMEljdNwA42GLgeerfgkHgdjuuAVPAtRyR
1qYssPbbm68zcK3DrtrckIzYj/sduGT1GSvDSm5btx/mK+IORLZN39cxxuOS0puR8l3slq6MP+fZ
H7Pha69VqJ+6PZl/ra7tpIde9Nwncxslts6aMu08snuTbtetn9VHGqxfHQUw3XoEyufO7pkAyFV+
xAXSQdg01me8zPIOjUqN/d/A9w0W8POxKWaM8VH2wzKgn33fo0RfE5ah1J4E7mrNzqXp9BQFToHv
fSYRI9gG5X7aigqQATeAnQQkafEh4o1KTPoZQMZ+RvNp0MHcx8i98gjIocrhenKHvWHmFYtimgtT
PB/HsJVEyKanoMjrfDsVfzRUUMhMRPmometbfCa+ZWHsmTqDF3Wn+2UmHC5GjePTd+VhaaoHKr+w
9GTDETDMy/InC3WrrtLdADFZ+D0xqzsVoNCx9Xqn+KRQUz7PvMo8DpOsrD78gxmn0BYrw4ac4dzU
OLrT9HlvtzKDEvFFhbBwUOs07YBOU4O6sAKCe6RYDcmqboEQIUSKV4vu3oDtPb9UF8RdeqR1lv1f
lzOGVlFcCBy91qeD1ej+1/AyFHDlx+9Ccw+jumKuL8/OLq4z3wlJ+OmVQXifkPkzh5CQcqWoY1Md
pmBKGq/1kDAI9+N5U4pIACxXfJSk3mJFItr9NOZzf4QQIrl5FZE69VpbmTxhuMkffTYhDJVkGPVg
RxyJpFWLiM7AOk25Is77/CqZrr1/BvmDeXlvHeMlQj0viU8sUbLX6TvidSElqn/aKJFzWnnmvfey
//pHaCymY8b/zzDfu1K9TuFZeGWCja6Qe/TrhdY+RQBGQGNu2YtIiWBwwGw0I5yGSVMx19ShtyrJ
4zxK2VhgfJxt5oeuERiRT68KA0CiHEbTKjBGdrzMnCq11qiNJTKrw49edHwPjGBsXai98SsZCcH0
swjBbBdzAXZ88MP9ZQFmEfEWrv/yA+ySIrXweSiCmlWcWVbffMRCDE6UuTaZx8U083hxmp/2YdrC
lcEgb+PcLkzMgxd7vpWOteTbcnIA53JgvfK736ecqO7xlsbdx1bN82nhKNm72ZLqx1OWvC+dFBH/
nLXAsNM+Um4i5j4lWrjXN3jnZCCYzwnv76lGNYgsoMoPuUILP1xdy00q+SxqhvEgFLx8dY8WWSBF
9L9TM1wmtY5XnjGlxkewHXjIh3swfr7RESCAlocyHXLScsqXw7Ao93IsIsdjzBivp09K4NVNpod6
g7g+2u4Rw9KZpVzdQ/aFAEQ7k8ihCey8KrlJLn/TrM0z/KGSMBudKYLdghBEOQd0Ah9JJH/8SpCR
j9tsdiPIqB8soRnk72NWtc4QlxqaA5/QDZxOlEZE6FgLkYcyhM+kTTUkoOCFnAY6BG4IwGflFKsg
yqXu8bIoZFEGGikFr1wMMwAeXk62RpkBiK8B39qEzIvM/F1KYn3+6smqOEK8DqBrHJSfyZxHGpAx
GBjcqFWLba/cHIL7KurNiH+b3yEIK8unGUig13gl2T38we7sgzowmvci5uZwfDo8iS/Sc8HRUnK3
5npmNQYAu2yKPlDp30cHbO86jX+kChLYit2Sq0Y947+/8T99IhDhRi8FCr770z+ks/7Fp0CSUhD2
NN+sJZVrodPgw0HKs53Xeg3i2Attr+WwAaRQZIsJ0EJ0GFKkxLffhgCnsamAE1T6aMu2asUKwTgt
nyDQMQx5fuEQ7ATD28xJq+ChLavvSCP8Iok7GiL5+bkjx6cO43pyYVk0RAPP5b3ff2jOtg698SuZ
rG/nvA8/abM1d35XnuwECeGrGKchPNmhaxw91M7sE5gYfcJhcwa9JlNC71SpBIbIbS+TXrD4MaWT
XbfHWGsSNxL+zsbG2/MCRazld3ikon7uFDUzo3Dv2tfiFuiFLkcD3pnfEuGvWQPoqO7ZPSDQXoF6
gPITRwzgj+7AJ4cnqDDnOSneTm92wcnb9JFLIh0UVixDFFqQHvzQPTiHL5ALjylDrzthTbkrbRNX
BGr/C5787QkJOym1zgimnXv5CL7nYgOUoe+ETjEB3CGgGXpQcsSPnM7ZnZVBTkGiqqrYJAbCpY7M
5z9q0Ah4i0gaZOB74MJgUcMtqBf8zUTcYFkJgAL84Vge7GjSDLu7oZTkhAe9DP/XDLmXN8+EV98C
3UnCbccZWZOxJEwhV4NyqSZ0g3Blvt04BfqIUw5NYTSDnOk+DCf9EnDEOKvU7wvZ6OmHxKN0FBle
QSQymbWjXmIK3NPz/6FrmRYBts28Wa55+wUCxwJUBjkq6QDp78NPmuk574t53S3c79CoAZU0O877
gBj5ht4I4IoocwwQ6wrXoVnB61RF4eMJwV6zkzw4GYuLyQASZJ/MwMiXRM7OBdl+dkqKGQzot89B
Mo6jzfuL7It+xkI1+a5nITgWSTiZPNf2wibw8dLYt3GjVXJmoyzef1djbRw2u96NATf/gacciMck
3GGoVPHap2HwmzGf338lpbciqxdFfYPMk51M1EpFDWHVVR0B5Ln/nyJ6Sq0GtlwSoBrx17o6wgQA
mcyQnpG6Bx1QGlXTCzmp+fjYf8o0NEuZNLr7LKNFqB/YIbbvJbC0csGhM0Q1g9RSHdeA82CUMhB7
npE9PYHlnGiqJ7yCKyuSIRaTwQKryvuoZfnoWjAH+vPKNKYdRc+gAOLgZzOuw8NfGoZR1mxYAWWc
AGJDfVsb99g2nHuZM6bVi2P3ad+xXs3ZtM69YCmTIGOSifsmYK5PwlzoD0kZau1dovps4aPTzGL8
LScjfD3enrQerpD/UP7X08K0/xeAkuC0GysJ/OHs5/M74miCKNrQU//Q1wBgE9pm0e2LAWGRi0We
d50e5t1T6YKgduwjvCbzGmkfvomlesmORyU85Z67O8d1KA4aOxQBrU3xf99FP9piwK5q9ZdfLKsJ
dTA+TCRPyiTNuZeDjiIP2zxgSmy8axkYTTUakXngGQqbLU583yQulSMqsRPwT1ATbcGfqcEBG4HL
fTb9yglZzw1yYOWktuh8U0kjcI6tC+cNQthuIT/m37xgMSEYX+D1821UQq92yZj9+o3xZZZU0Oq0
tjXW4CpwqMpE4qxobwoJG7ITswO9FDLopOSvw1A4pJppjH54KnTCslg4cZL665G7vOcSl/Sa5IT5
ZNxD2DyHtiCQ6sey2TVg8acRNbNrSgBWb4HEIHNtD8/wOILmWPsYCM9d1Uoqg9YIllrXNWjiO6CZ
7iP+Ai+RoqITyCR+bW+92vS98McclyU6KESVg7SQWZE2CM/Byf3e5kpkMQcuGk+my91CitfnoXEh
xYhKtEjrLq3bfWM8w8vUhPbnzcHFG7uTKzXBe4RBuW+l6PzE64f+ZRQ6o09FzkaIbQOmYOGQkNkF
jHfIgK72gfILF2Ns8TN8A8hROgXZ1DHzQBDxhG3Ig/Mh9meWe5GuJkoL9OsMDdRJ82tBow+59dSe
xZWP4+cp9OEXx/NbljdVKSwwjGToRYaoTuzvcbqsl90HBlApNJW+wUBRbEbgj802nIbJY8I6o/ZK
j3tWKw9yJYCczYB2GrFKJtvdgUrZJ7+Vpw6ZagvLaGFDwIefqhxVRYPovVaNMTo/4mpycIKtfCRu
BCa2OCsI0sojDhGvs3hG80sc60H+sntPwTWE2Wu/3wLSV8617iAWk7h4kT664KJuUB/m/drwecha
QdJkgvde7wt8U27I96KFzjf3ATAs628q3uxBiSASFrbhsxJ6aqZBBl92XW0llY8reUmpeziSct6c
P1g+lr9Chet7AVBJxxP8hBfBF6xutbjdRCeWJAmh2J2+9YGc5PT/pwG4N0CYAltIAa4yAlVMR2yd
BwqZBi6b/UwF1+pO6ODoLXbJ/GXASJKZG95nz4BCZ06qk5OZYPqxj4kZHu8VF/CTk9ag+I53Lyww
9My+w55yiijLg+iYyeHbNggAG7rPp9nyzNMBOqvXA/CockOOwsH8tTGVrG6YLQJgx4hMZ6EtazA4
6a8pcBJO9B+UANmULljLpjsFE338XvSTDopTnXRW5N81nHl8elG81BUv3iEOOSJaCoVvhwP3tmB4
z1vLNh+8uka8UwCGYm01eYATAlTYRGmD/8PAuKz5My8IGHV4lAvCi2V30lr2kkTSZExn2FgKxFOE
McFBFHpr0nJWlTLkmX3xNcMCy0qEQh9QBLDo4CSj71/L0oszrNLMhEP1qn6wFU9+keE3IEKZO49D
b6i3zvORVyLx4UYf2N93zn8yvx4dRvFEO5w6cWcDUqVyB5v1GovUWz6w1pnX8crPZ2SEdmlbiXRE
rw39CmCV9/cO4dMNoX/waQxqw8hhjduh2AvtIUuVsoMoqdYUxlBZkOSSzz1T1S8dksK3GZZc/ine
WTB8zaB0km8YyQXJWMPwN7VfJDV/JJgy/BpGO3FI7UMQNLQYL85bAaxloxeB8O4ddyxozDwNgY8S
0rd0HFAo8211TayOk2g4YQ42oa7qxsF1GEql522u+4AZ+DR6dIDV4RsCbB4sePt7Ga8xr4A59WDP
XEPcCmpYlcjt4K1gmepaPQnHSnyjoLn5wpxZOSZ032lf4G7A4/qYd+yDkwCROrtX6h1SiIRsP6vI
6vt29fCrtlE4KiFZe3Vu+tEI8junwEYC/CgNfnd7yAeMpqTFqnsz8j4hLsasAd6pgUMxoVuQkxP8
ospernDdT/tfB0+9SEXtLvf8+xDQHGNky3qjacqh2lpL2lcbF86KFXppyOf4iFLffaBrfXNNpn5B
cL25YIxo5IQJPZhTqmuYymeEKHQiLiIzEW0zY/kRJePJ1d51TkT84VxULt5HXPmgYmM2m+/J5xp8
is0+aqVVcY/dFGYhiuq6L39yHTE21MPNaPV3xtjeK+MMZBoBaPgkEW4iP3MiyiVuXuI2f1fgCSRi
4pf8d43fSoKOFWZe0907RSO9BPNnsy1LTjBi+ukTccfPeLJxjxcLMNCl+6y8dpjyUcFPSOKWv26G
p7G/d3hy9X0zyZMQ4WRUYunRnmWAjrhXV3xviT2NaGO5P8JH2KYFKS0ax310een66/uhAKLoZE1s
BwG4y/Vx2cdTafmDBuCZbr8TW1ztGmoE+cECx4H43oUArQA685vBw30X+Yk7X31ZOzHiCoLkEew8
aqE1Pe5IRJmlCrCaSUhXd/QNoJGRzm7tnnpDhBfW2BQZYM0tY+aWyAnn+xpIEFG0gSiI6Vf4py4B
Y4sXrE8YrN+z/tjaL8MV0JFMTDbsnHH25lENESbnWHaymqTrqbu4L7IPIYTmKkuOUaDr1owhdg31
6IMf+bsaduA7dqUyEzdB7z/RWRkzGFzxBQKc460RUd0HBobHP+FejKqdOsNzrkzQ2ppmB9G/5x+d
spHPYkYh9vR9GUs0/NYSsZ5jWAw3bdqUjeAFawxTuwZLaG7nAVV2+zTaeH8oQ6O9HaU0hT4Wvqr/
Ml6SAXR3fMrObrVhR75bqROSueBszJOikvR/7WrM7p/ruhHILvdZXp5ERKK+/F7CyG/bFTsYCoDu
brprXMFx/luMvPUaIrpgspJb41IhqGKjaxOdqb2Fd6VvUsz6fdPOsE+0y+g9UoFVirhp5eOu4gtg
d20qQHjwSrS+ccAHK/3hNUQRRY4m7E3s3xxpSQ9eb19vrcmjlHTSVSXZnPBSxwERcZDeeVAR7PGq
kNZiLfRgX0YvB9hZZOP42DE+mG6uuFS3s0sCcdiCLvRlXvFK6N23NiruDyW04IenA3sqoWdCGolB
T3TgwPCL0NagyoUyStxrH0vbn0AGkK18POH7AFubdzDzI7E63zKGs/LqYwhwioh3zBUO1j4b9bio
NwJPQsRznuz9ig4GTew3DDA1jaMrBJ5ZupMwCXLtXlejQK87hIL5VmqB1suQSR1BbVDAILHLRKSc
sklo4CUUIoeRxkYRWtYpEeJhyU3fOw4w7dnR2R/49rjsfeBtce0yly5sY5O9wC5BR4yrNidh1eKf
xO6Snront8WS5eHI8ecYpEIKEqlnDr58NcTNDgfDWqTBmrFwsTJUA+QjBMiKAYmoyrU1h15nlEoz
qmL6nwTAW3c7IxUju08Muc1G4lr3+v5ajdBwq3qouj5Udqzk3xWxOeWOaLOl59yHDZkAE3iaowsO
FoeCo9dALCM6H1KNp5JTXvAjyRW86tFd53OiwpxGyuBGVkbVuA74Kr7PnahUK4aa2HvDizmww48y
eqyhyeK4h3dv9+yqsBMMNhISkYvtQR4JoFc73stsDwPoYE3m61nwyZKilQx4NiddDCqdQGOwBWbw
B1zT3dlalWa9GE0FJ/9KMSYglFlyoo5TRytwKemKvNfncaGsnVkpUmKydDziiiqODM6UUvDrB4qL
NkqvMd7tY8Dpf8n1dHmcdxvmFlqv7xl5O6vCr4pPMCvWoRrFm95eBa97cIWVqxXS1g7h7E8Lg3O0
WB81kWOsaVpAEq80ohTtKoVo0MTytR+WFzOU4wscHC15bnmAs7TUstxm96AT0TNGiGlJkWU2DNX7
vCsZMvdkQPntKifZkYyNSKSYc+SfHz77NhAkYCi5yZ+f/Og8wpUEOm4gITZO+KEDamNeLRCh5nNE
UECFTY2YVK7fP7lAmT+E17KU9puS4mlE0g7HNAneVu0eoHX8Xc01Lo+zPM9pIDmrCl6vLZFg+yyY
R43DbxRbOYT0oDwtnZLGHTVO/J+r8+jsrEqXFxG3kMc6QiKRcJnup/61SB5B9mmHRA7QUm9r1QZZ
PdrU9GcaVkRAs3k9eVpaM0YA3C4cQiboWU33vZtNRZm0px+5sQgO8R6T4eFE851CJ3X/Ztr6+eVj
oVD8DVqpDAny8VFo8ySRtwbfzb1uUMR0DCFnJqqpCV7FTb1HuspWXLcjL52keyHeLP2cGfJN+D/i
rX3QXsUGZsp2gNKL1oAZjB9ROG48fQffUcSnVPX3G8Jyc8M58i4BSC7BlTcVWAFpOQlIEJgfBHeQ
PqzWxmvVcBj+qtN5e0aXJ1qn9Tq0t3Lz5XzI85A4+7C14M5J9CnRfC1S2d5SZgIxAkMzPtaVbUZF
jwCIzl23H8D6Wmdll7nvSVp89BBnfap4G/inx1CFSP4kv4edhEu+BFIFdLeWPVV/yaS9uMogQ1pT
rya30Qi9x+ugZ3ARQsG949Khf90GeKQcnChHlKpg0prCr+HlhZ80Aj8yV7Y1kLT/zN6aGehAG6Sc
dPo8EnpQZdibwSs6iOSs54dHIz/TnbXIew/mvMDOg6taHWShnAxsNv8fUobkdBL9RXk/Tys05gVY
S39Y0C03H++tzJHf6NXlihI7RCbVy843MJcXtaU6tIakqpbS0ibbI/XmkoxvtXNDMlmqpuA+pg0A
jWwYnX9SN0xTU/VKpaduzGORetR7djKU+1fdRzRlY4SkXENkd5VmLAUQvqGP0I+4qTh74HoSxpBG
syuWAjoqD3oiTVQsOpnIGicMBsnTQsYylhGLtj9rs1XwD/emurSB2LRk3ku5LjGoWzlOHDkBCTGK
0F7/PnazNw54Ul7TO5D/X1ZxYaTgXTWSQmBWTcYUM3BJ9Ttk+OdqOo6wFMlnAc6n2uBkeIvDf0f7
h9LPmefGIGQWJ/OW1ZSTIOUb+YPoPkwUDFFYUOHu8Y7ZClnAF/+Bq71i2Msuc0v1NF6qofpnMe/t
rT9sx+KjXj6tBZ6/iF0WoOqPeEu/MX4NmHLUkfhcTtl498UbJNpb5JdSXxPIZnGmfhRxEdCjWOD+
kUaCPNyHusUNaVy6OZ55iRb2eqrlPxrcze1dmqWrRiWp+xFP8rYwTr77SDad6cp6wkqWLLW/SV6K
KLtCVkMx5FlEMS8zST/Mg3LCKE+b9d4cQIPiD7nlGrije1kFbZVFi8uI/wXOrYSY+5m2nO0g+mZG
OP4zy6UBYNtDWzeQETSClShDEDf/q5a8Dr9GQ0M5XEguLq2ZYmTaFP/wWFA7xAu3TYSXWNT8oUQG
kC794nBaoL0ifW8CeEDpf20Wa0ouqdxVibbhhvxj7LmcdRcfK3AeY4N+W1Q3SyvNmvtSI6K8Ahzw
z82mOCXXR42h3jFgtCU28SAw7LjqGP6MlZ+JH6jt1PKZgiklm4dfFKUUlZy01fIyEb5PsqzPw0iV
S6uzdKy6S2etE2JlPGI4+jjUu0t+a3srM/ZX2EcdSfd24BkJC8+dMSWqxiUWf0P3bj6E8DQWs6NK
fGK3LoC+hiedZn5RMIYTGmLc7Tl1mZt9+T8xuyilKo3pYoYevqHjkSPUJpMTtMc1leAceocWlgq0
JFvWPkzsCbyurNO4JrZlsA3Tjt8G1eG9e/TAHdH6N02igW40brYg5l1XP1g7YbKAZc682XRDwY/L
iLtZJ/359ohwK6yAgM7MqoMWT3FTLcpuZ2LoIs9DQMhNe/g7hYTgG+lzPlXoAidioOn3SPo9LKTu
e3tmzGDVDNMPPBuPJm+Chkxw9wkD1bueLyHwAP+dYlstu3r/ieySKFxq3dQzemqe+uere9u/OHFw
sbubLhSDr/YKmpo/wATTuhGmSZr8SLJULPOzznbQSoVcPTo/08nMR3Xduoev0aNT9zB3AtpP8pXQ
V8QzfkkE0/XRJyIlGkp71jRarT+/lZYgjV7u2/Wv3n5N5yLRwZX3KxzhNDwbpzfDnGUZoRmlmCjO
9UdGjkvvp1pLILD0Ej0jgR50tkT+mVBKMbc2XAOpIQTD58LmCBJPk6x5M87ZGJx0GaP9h492co3/
hC+NugkCCZ+//DWNCkqRuDXYV2NXgFkuvJS3nMTbh4G+5cIwfuy92S0JDgDd4v0sZzxkH7WMw6QZ
wjqxpmWhERsIVt3LggA8I6G2mJ5ssbD+c9qF3UgcmKVIhIG0YPqmNu0TROTWgWlB6RIwmxkTtvCl
URcIRWFXge0MQUeRo9UwbciAoKVlpr8FDz6S2n/aLc/CiJuCB82+mEH1NAImIx+DCs1BBxk/Qolg
jSZ+aqUVTmpWmpFOqbIM7Kq/9UfjAidnDBu9BM6AO44zEvxM0dF3CtV10e05nTrIT6eaaZnx1kyL
SNpjjeV7Fs1nMyzltCNTIeU7fUOiBox94VCc8nrJjzaWA7Q55ddq+ds2krPaR+gnRriY0nf1pm73
zZ2+kF4cnF2qohN423buXzC/oQYZnczFZGadJV6yEt9SQonGj3cWGHbomndKX2GXPRoU3qLEDGXW
RS72aPHzSxhmeHN1mz6MjeanXqlKUYnzOjPkNvp4otT7AUPcqHtNmMjekws9bsp0lDirRjURqWFQ
WmNksan18kWO8TcOhKQIXwr9vVBm8diIi+5g8PDt7g4zaaJsOo1X8fkcxn9O4Wsi7vfQYPnk2uBw
/C+Zs0UxopUYGzSiI3agsEbGeQPFuqW3EQNA7C83eHr7w+2aBd61EbvDCYZdALVobiXZeehBK5qS
MQC9tUSEtnKUdf+Utr+/gPOTa4zJGEOK1ByOA7ByOeQNGY+5k2jO3ISYYptGdKVTj5xVs9VjXjrV
+bwCLpWONExQxejSGNVl/JzIJmBHGAqMAKbTHgOZ16Z1N29NcNyHsBuTQcojC8HnN641zoIb+cCR
TSEK8tgbBaTyLwUqSNfZCiLRoBT21akmCWq0w/iGbCNn002C9bw4nP7KzVUA+3K0Z3eHV37a3Xk2
Nv6vfUTGE836aUFoMQ45iGiupUlAGh0yECSu0Yph2S4ZXX/y5YqByT1ODK3CVR93fE7Yf4LkRcN/
lqbVhzGj82SY4RAwJWartkQu6sSSBCWFZfWsYz1O0U6T/pq7ndeeuV7MHaTiFTPIQv9Mtd+OhcDY
wc0CWfNxBYEXq+/EWGQm2QClbL2tsYOnBi5PZU9Xj/SXkZMShRG1lx7Z24md8Co8rD6hgfAf5jKw
Y4WQCX2809JgBoUV3yyFnJ2ogO/1WtLUWojNncIZcL58Eke3uJLDvDkikuIIjzOIbyC8ZTuf7Rdv
0W3JyYhNy8SVvrw7voxhAaqPIOBQ7kye4kUs0jDwkfUun7dt6OiTSoKplrPasbYp+CM8tcBY/OVr
ps46YgHMafi+qpELYKurTyK9oBlM3oax5moTSdR1J29requbSETMo7bfmfHYl4ACETDWTpCoa4dw
todfNrmIm7gc4q02TVKZLJv8bsIvZtIlTG9Z9ObXYi0z4F6m1n4qVRyiawb5cgu2LJPSXpqrO2fF
eT9vixT4CHsLbJr2nqX7r2IO6v0mxHbu4etkcngZ0rswRiQ5yvB5MJQqiPLBl5o1pps03+VcrrDd
0w0f0CkrtBlsj8WYrxH7GlgpPrlOAtrwNXP3CGO6KLvHiDdASg2VI08/njp9QwmQgt6/Az5UGTiH
x4NvXTaY9/F54W0cdqO0PvLU6dyqZwu4UQK6btldNUFlV834eXxolvNVRm9+F+/Gkcgk2/J2inXS
8NwR4FbLD8mp7gwnrKnbY/+R1bWqKB8T7xWfR0RHH6dElhGtB1VCyVrMoDhAw2xvqon/HEjNUo4l
dYOh93DhrXEX4jyTGnzhhHh40fzCpFuKOR31FuBQSS7n5Si6mHM8+P2iSDmDASOShgnLYL+q2g9+
LoakdDqxxLgAUUNzXXa31dHFs3MhYK2N+oR6Afyte5DixIYe/lNmWGngJwJdTQk+FXG1SmwKs8fQ
hAFVySvBux+xgouVtqyo9O6IIfOPj3sVdFqD2FCRmF+39TM8RO2N5crmR5p07g3k5BtUEfkdcdq+
oD7nAN23jUAK/bE1p02iOHZ5q3VrImREsCNUuqFFs3Lu8r2hFlgiPgQzITui5esQLDv/fr6cs0gZ
9IUZM0Ro+FyAeLR1p/37aCBZWgk/Oq89WIqSv+ccTl0jUbsXFWtQx9POOJCaQrLJ3A6TflwZDQnR
37+xNSWxpSADsDSkCv8Kz1Tfn46VOjA8kmXRQIJXe+jeZJFDih0vHx9bwZ395/Xdu3EnwctMjGtN
saWKswc0CNx851XCrJkyMxGMwAjLvy51hwTRsSQ7C7iEWOu7iX67Jy3lVv9QQQhUTJG89/tkhnoj
xG9AJ7lyiI1OHSfKAyo+lxRHMkv3ZZA/nuckaD0Bth9rXnTLoDMCZHrTV2Bi/JhMb015DRXCjJUk
xzCly7iwwWuNWr6Yf8GxSnQd1EbzPy2S/aeMRPAW3iN/fjkfR8mSnF3ufg8XSfy/yJiGPrtAEY8/
5yXjp39Gs61bHOtjrkvmCoWt7/TMNKfJEfnsTyLOGFGGaxSf/HsgtmHveIcR3f8gRKi5N0Dg30JI
oDXoWsYuCBnmC0pIk3NEHp4GbhnHhOylGSYzRsj6WUNkyq6/NtmhA0UQRd85xIzscR1+KKU9591f
JkZEiGVL0oESovNNenGm4IBurzwgkFPyRZo6ByWxdPYFFuVQ/Y/ccraivxox4DxMvLn2/8yutybl
dgNvT4JKA/+Wu/W3oxVSXn7HW+16bpFg47/S2yfwcsskfY8vicORZ87JlQ1FXK1Nf/MVCST06Rn8
aO64RqZ/kmDFY8BVh8iynWiHRuSN+Kr/lY6GVAr9lnQenLs6ixLfA8Uql+LQ9Mfu8fwI+OJ5kaGc
CW5j+2uJJTACADzG/xI3N9fIDPh0Za62LpP2LBn1OodejlSr4YHoAUaVeRoUkGSyKO55AdMkXHGc
3uhlm6/6tsMZM9oPF1t3loYBl5UXdBNS35EuK36dtgTNpdu9noquY5X0ZEOgDGCWpvzguncpMnqv
0qyTLikdNxTlWq2+/x3e2G0i+Zooc5qMJ5ij6jvvdwpSo+QFLBPlg3ECR6r9TjkJOaFRyDbS2GL5
WZGsnskU+bOsZeFPtXHuoq/ahs7ysGGEyCFt5ect4FBLW7zfnK3sl4jYP5h+QAqPl5Y7znVUZHC/
Fp0lmlsSPfnSJQeB6P05TI5ALPcdSpcv10Ipyd7QyiyPVC3WTky7kOhkXe1xKNRMoJkLxQUAmpd0
P6+DJbrt698d+SJLI+NR6ffve9PIIQGctw8xz4P46upwxn0v8IjcF13qKhYW48WBng3eQbXL2NcW
8p3wUjT365JsnMo4moZnL+UN7XRbVXxMFF+imXII9xpQI6PxXMCOOK6ySQUZR12Y+qXd/G9QySYC
BwsZtXXxqBQgUMP4mMoSSHwpbOPMFvprSppoWdBxiAVpqK3XEviCm1wLTRgiclJm3wUDtr5PClee
zFTDdcBbCqyTKrhBY+9q66IzDsrUDJxzl8N7TF1/h/V1WKVRK4Kpwm2ScOxX4BFQwG56+kLjX7Uw
OxjwP+gZD7hrt4WB4hEl0yhn/tKjV8zSPAGriH6PMfqmcbenkxxx7+6gjhQ6T8IAxOirs2ccdjHX
veyr5IMIm0fWFXJux3OVnWZYbj0lLuYKQrpyY9tjs+nc4T7CJqaignPTQ/UPYlFKmFadZ0N6ZZpS
Ttf1g/dssa1EwIRRi8dXNXT2IwlJgOLaYJeBo1G/t18XeWytcpvVNG9L3JAvpRA2k7qOrh3Kdrps
GNxZL2vCjy71QuSzNhPCZm7HiVv98+AfhxUnvG4R/wgpHVc2+4i95pWpRlm8HiFrNdRvXsVjZ9Yn
i6GQ+0UpTdyMq8pn4BwqPyMMDIuUaYFovr1FMzvTi/Xn10SpzPN9oXttp4mfyZKGvEjQnn2yImOK
fMzKItN9l4xgmixu56tpSgU1c9gWU/PeLtJgijfG/rqnBOw3gejdlnSmsSqqMK3ecEB9UTMTQQ9t
STghvBInQawLGMKazTr4XzPc+AjjXMK8frYX6fpwbhgEiEfhbDT4xu2PChn5szxL/asM5GkbnKeJ
WqrEvPv4OwNZJnSdPnuycL+wUkGwlVOjWqKbMX6ntvwcp9VrJFrSkca83IQODP2z3B3kq13XdUoR
cvYP5lsGCEFKxH9pEapQoTi3i5W44Comlt++dUVEoNLb0jUbwmclV8GPiMhHwhym4EFJnonzhCXW
4zg39Kb2sHXx5MtKAdpeVdgWrX1m3kONva3nsYrtNY55+iO8SuVi7k1RbebvGbwZ//ZCzyj6cppp
cufVB65kO8TQBoTcZOy9e3Uu3IZW880qyV8uRoknNNzaSM4DdQR7u9czVXllDdBd+p13ZF5+Uc5n
M41nuAV7QBUJ6arXEGkREDKoY2za2WTpXacygs3i3rSfJxukn2R40jcPJAxysMgawrd/AClUNJgu
rvBN++gR7boDtjnIKQB3Fwv/mPiDz1TM6ttWqFV0BzoaXQ05MSaTqIl2ec9WYWX9d0oHBs06zJAP
Lli2AhXQ7UHBCkwEOdoMBI49QXejVbeUvUyop+mb1+uHxOyOhpJ7G2DPDeR3V6fVpP8AJEfsshz6
DImY7Sb7wdJOkz8rYPaha0/xbUO4Wo3cTpWBVLtlduT17xuYubshSh9szBmywuc8SaF40I/dpxn/
94H0zTl8PvuTU2wQkFEn495CPAliTAjqn9yxcOOzDyS7VzGRq/kJTomRZBcQQp3ZEg/3a+AsENyy
Vo7HuwSzVN21dbwdqqcUuJAJfGydvA1oh6JyuakPNJuHWGdM5AS+cmxdUYdsC1J8jVkw4Ps7jOjW
9gvhB4Px0KsVCs0ptiQKqrH6vKcqfPDE8owFaJoGnfdz8otjB4azCjjKgTKouLOpDhhK4ybSQi4N
rWVo8L8AHTciuQSEXljGhYh49gXHKNA40AIIpPtImyxKo/a38mX5R2JBVO/Rih/pU7KaHySBc4E6
d4ug3DaKnFwqZjn5w/GhidjwyGA22Dl6Ctd3HXDKNRK1ZvPCT/1bqarDxg12t7MHCAn86jfnwW0j
tf5vM3xFU9hzn6LF4dr6wrXS6+D9Yga3IXZpaDx0LCokQg8OiD8AbBTXx0TTSiQU31eYbG7hSIM1
Z7NsrrdrjAgKBYEL1uteJnv18vEgFywQ2vBXbpo4QJQ7FbH5FkS6PYWRl+Mzf1aUwcNAMGSpIbAA
4A833zsb+/DC1mCmIcpKq/L9vxiOpVbwnSW1siAW9rinHTnMTwSBFtFA8hrQOEdfb9TFmDCM38IG
FBrNgy6mLWpBT9ZCmSElNzWe+UeLntSWKG2Lp90VLqaGzU6vTZFCapmbJI2gZ0Y/6YpebKdLpygC
2YQHJgHFW7GL08HrqkIpvj7L9Q+of3phAL+n5M5I5kitjpnlaQtMXUF1pz1huPnlSkrGTntCT33H
oG5dv97LkOCxPfouxvvTelSKUmt9Rr35DUZFcxkPhc2LTb19qip6k9m24L5daGU36AHCmTRh2wPR
2lVveXtDZFvUAMAb/CduXQDVTkbwBWV7o29hCW+RZ/7aD/CcQ5A7EFs6V8n/i+ax2ZPN2/yYK0GH
lJXK7ZnQfbE4TBPShKXMYoTAxoKZj2y7u982XQ7C29laYExN+tcG8VUQ0ph58kWyOo5cSTwI8mJp
hCTbKcEOx82EqT8i0RTv6VPLaYMwrZsS7KBeslQrTkvVp90h0wBoR10jWNEzQHFnof0gqFLbeKu+
BIRgEYRrdk1xy3SOnS3YXWkN0YDkqIquUSWuOwCQSzQ2x7ke691sZR6rzhVq5kDUxIKwEXIBXRUR
fQK9AxwphpMoJl2T/s+5EFHOIUAwATIWGlS+xO2tIfGX/RAhAMfNRArAHZFokcQI4BNgnngTuKeX
9nFJCJKbfTNyWZKnA9oZaKo1TmAC1HcPcIfYF0syRAwBOiZiu/CS/HSSFfHHgqIdZaaBf0tUxMB/
+WfJ3TPT78L7foezJrzO6erMFpMK6f9d8bDVqzmQGfm0wSEt8qEBk/MtjICWnFjrSjyRrK1OCTAe
fBuli2pOhaIRjJfUqkdCHb6s8BQaBrJhZ9JoNzU4Yq4QSkpF1WhvZFBLdQ4iAWw15SqiFhOFdATM
OX3anRn0lAmmtNuHyo537FFGbOANnljb27ziJgBsb3D9Cko6omuoxoeU0CC1EEqMOCMeEy7tDK6r
nUDsl3l+sGxwsQwMe+C7hrsZKWjf3mtJnVX/omfQgUC6kUXxWg9F2C9eZVJ5+Uj/abomrQd1ie90
6yznS//waTSF2uDf0FXiam8eXigmwGtqBETBLTcoNCMHdfE2c4+S3EF6RtabFLRlkv1IQTy8ZqFu
pnFjzmOpabX5J98HXjougYWk7UQb8S+xk4sHDYbzD5HEPV0+0r03e9Hen4Aje9wW6eXiSZKjK7Iy
kypQFAkvvM6GDKuLopr/BeO0PWyMESFbvM0ZsOtDC14HRkOkiUqc7C/rXBn46huX/pBH4xmsrCr5
T1DqvNZr7y3KX0ziQX7GhYL8cvwAQN7XPbyOhb+II3OEgoFutk0N3IyZmCFAi3McvmDxzpQCzcPu
bayuh34GQeSjH66g3ZqmFomKmEkAIk0MIYAgPkpHmAkhengrynnoBjVLDx3tZR1EZKF82MrZmxtL
wO2NWcAVXd/UdWuZCmsJN48J6eLT8+rctBC98PQszA3ehAgzdfr1ihAiQy73cY1gAnJqJnMCUW/a
K6MGzWFfEx76A3zJKAOBfyOGpH+so/ANajYtSAfoaCvJEqbtRjh3IkruNI7v9hQ4Jmhvn4lnWIKs
ZVlfjq6iWTwonXXwZ3b5LuRp1u/fu4BI1M5CUS3MofAkjSLulULUxCo3DyugL5GRnZCnYM20R1TS
OyyQBb/TI/4XpQEnJsIZlkKTCvv0/4uLPtcPdxoXnQaYyfqXIbSqjAVc6qsIOMAYrq12t+WsN2sf
FfepUL/ZyLBNDxFLjtQtZqgKlOU7nQoqLfGc7pg0GVU9PEawxxs0/bSsVjwTuSpxsHAWGzaqOkkm
spn9LhsE/eASXGIzcL93uW+V2qIcLohR7TyTfF4eEg7ti0VxdLoAxVwvbX4ewWYPSPhkHRoA7UUV
sTukBP746g9NtfjcfTn0yPPE96T8PLVw/3zsJNpt3Vf7/Sef/LH5u7gvzRcHS+ipjNvW4/gVXNPc
nBnlZ+MPYEWslawPsY0aegQHnIkaB9arnYGiB0JEebz6rG+5BY8NAf6KXo7+zI1179/Vtn00XQD8
CD2Qt+EO81cJcHiWzNfRRBm/HAnVUQUgQ7NU7rZTWjzAVpqSWIqXpa6xEF8GwifTBdY51OWIhve2
EkNw5Of9RknGX8l76Hbv3W7UIwy9yheRtzPfB+S3CMDDJkQLF+a4oOfpJIn5uczq2LBDqmWtPxSR
ZGMz4SV8V5AlSgdjPBUuDMf4G6JIAFrG7WhqphUZ4VQx5KB12bERPCnIr1mos+xbTLhygbN3KPxM
yVSf61yHQW23SHByEvtAdNK0xIRWECj+lXGvEYe4PaIRLxf1WZVzTYBhDH1fweiSZGtX3eOnKCnF
MZd7cbO9lIgyzkLNHgDvItNwAvHjtEEETF/OHlU4xQLPVBfD9crUeLBr2CZC4OvbB5vyES7AmMoE
dLIyHOUAdotlV3/InUXThBqKRC1U6Am1iMapfM78Tlptdg3u8fOXQ3R3kdmb9HEifhYM5bcjraC/
Tmqp6x9E7NLI5ThHOUFMPdu1XzA0PdFXLD7VJYn8TcB1diaO5whm8iJ1DHRrlWF9hCxqxbiHq5Tj
Ww0Ses6RIq4rK86Tnv3xeCrAEEcn5bGtL06xdblJ7QD2h+uwv5N6p7KIYWqnJCrLtK95e04cRMRf
9xKc24Mrh6DPFpwloK/x5YtB7hrPwp3B/ixIt+TuWDWId9H6QIMUCS/Vkp2tdTtLH75tBQQF65WH
pkYpO/9DAV6fO2HXJwmJ4dDuvXwspwTXtBDgOUNE/H3OM4ZbMiz8cDVetRH1ukpU7+/7sLJn5tKk
b+GvHZsoeCpHjc/ou3iHiTsHHqRW2NQgy2zHeKrzyMNJPE4EPNNWn5a5F/Hsju5xMFB5Ybunqk4b
Py/HCyELPy+9CRy0DPCqZubSR7pkrEgnX1pPo/ab1EqUVRjyLDnHvOSzP8+5THc86n25ysoGWyqe
0WLXAdEALRz2e7sMuPSjgje9zXzyncdQwYJSxbDcAgXMTdg9/5pjt57Ax0/em4x/8ulZjQLZV2Ph
f7hF3aI/LzHNoZmMiqfU53+mRm8aE0C0dqo+w0n/h3mBo6OaLb0jFyD4A9b5paVZKkamy/hhzdjO
Q7kpCw2u0MvJ5mTUrRXl9sRli7M/N4T5tEFqrXdHFy/+aEAMOpXrzCVsgfBZw53Ln4zL+KrLdUy3
cC1K1b1SdR8fpMu4y+ILAYUr26tPfCbYPoOaLjSPJXUx1jTI+VMWClySlqPfnjm/Qnnm3UcBNuNT
uKlvAvgsDA/fR983jhEgAGrE9BnlMOdedpbYG+rAEwoaKMzaqaW86YxxzTlfBIs9OfxUtXy+RSb3
rmASn5gIDmsFC9yyODaNGuPR613uu43c0qBR06wbe75U2HcEnXtLmfWPDde6MUlvXRV09vbAZwMt
Kf230SAOnXwhotHxjbpg7GFcIWeBzGZqVbqNys5GsR7csM7jIADQn+5zJ9Cf8onHtguEtbrUJNqy
x0by7FAjo+3ijcqJYBgOXYVUdzJmELpq6+tVfuEeP1HVReI88iryFz5QiWhX7CeW03nWv1RmVH8m
tNaFtnhoFtN3WVvfaWF098+OWGd3Y6mKf/8EfOpqF3Ssfo0G23sYInzgvzsVGMTqZwwWHC2KwDeJ
pTVRoeq+S/vaS07U08AY8H7u+1UOwQlQjySAgSr/EM64yBGx7fldK292/iUunZ30Qlq8GRUjgTSB
CrYiGwiUPo1rp0NtPmqSInpY7hZleOuc6CqTMaLhmFYg8TxEvW/uZcdMUAI8Vat8xBqdm3XiqvbH
xGzA5vLLqMZMDO4zSUCXETpTJnJU173BGJy3+6ICNijGh+38/ePM9sMfAZEWlj7Ar4z4CV+VIo/Y
0m8qWlhPaFxFDLxdkfefHx3XOoKBBGN6KEfXH3msUQ6bBK1/naNlI8O5+re6yqRFFmNG6Y6HTLQI
1HY+IxNSo3/4nJX3pihew05UAeORVW8jPd3yUDbJ++9CGtHVNZh4Hup9IiNjvFz/6SzVmGKUKqsL
O+ZyAOEZoDSnZTQRchpuT+pWGMtA5HvnWz8JAi02jovWwHQZlic81eIfeh4QYmymMhjm+VqvJJ1W
rxCQHF4Gp7Le+ZzGyzDz+TO/4T6Z3d2dDCO/Df7LOrYE3rU5tXJxDg3aZFmyEeU/aN3x95ZB0MDG
pLiAmNiU+8Md85chjafIvfSkEaV8yPW4DWj7+5SUS4nzffM+/AJtuXorrbucpnhUVuJ2dxOovrwG
O/e6xERGcO33WwPQQBH9ig4coptVwQl3CPGjQmFXUxvsLhpURwZQieohujmLS1OVi7Tey747VbG4
M27EN7aIM/lr87M//TmrECK/9q8FBn+ZJgkhCq6P+u2K5u/WjYoKzTWAf9ISugLakqtY70hxBIQM
MBRvGss4S/4AGDpUMmKpFNZYO1G9i8UiurY5Pn8RtYdAdZ2v3a5SXhxYmxVwNrJWsjwOZPz2zsWs
B6NS2+3Qmoyw5plYKHurTQjE2893m9G0jiENcI85FjjmVUkiJR3C8+rtLKgu2wlRFkyeViDvDUWK
1XgIdl+AvA7oMaJsd3S+8hKLsOfD5YHlzKTRfk0dleFqWqoitvmlLGSxsMmf6J6nbd5eyTWZqsn0
3SZ8qJEhJmUWv9IigRSifXOx71pLzNuyVQyS4mIfi1ko9mmFCW+Adj25GRUp2PesMC3EePGFqFWW
mbpPeDjQt3CDy5DhZs+dhJXcb9VtmkWsvG+xqeMZr3uudCtyZeUOztxWm6JFIzMZqL2428sq86kT
W+1+OZ5rurAisYpTvxc146Np2bf4uHgsbnYi6FNbRhBGfJ1w8wXYRe2Vg8kdkf+wAFeSLur4s3dB
mw97ujVgp8Mtc0VYgBNM3rCOpXrZuKCtB0UJ/YmS96YHubYCZiv9o4UupDcUqfE/TDnmKgSoL66V
m0Lxa0nZV2fg0UefHID1bzmgrJHbiGBUJrJUm+N+odvHfE9a5AVEv+Lwt4IQgwwT+7YjdHwIwC7x
1mVhjxaMxQrLGEhcfDN+UAyLAEtrth8I6RGcGuUG2trRbXFu8ZRj8lemGoOoCcHfDTi6lvMUuEsk
Gjb9wlsihv/804wR54SywjBT19vnPpWmlBWcCEdbrt+yyVnk9nbjTHvsIn9MXXvVnT16Sd/mZwlD
+a1d1nrUK+HJTch/wYTOSsTGFTHaEQ25oYZ7CqRjaRSxAiIPbZKlduwN8+8n8LSkIhn7Mcg9zY3X
TZu2OomB3xVwvieIzfWiRUMB53IZoLtoo/yL8gL7WgR7FKWvmNjLri5SK8zkA2q7bFA5efrtbQLQ
S9EEuAmUxVqSvjLKRL3GrJ+fltkIBXSo8HLWuF7wjuhpLL9+fIGEeSGv+7YL2E36EHrGxOZMKaMs
g8KJVXfKZlG6CWECxtrrFveRZTwlt/MP2RO6v5aYCCCR/NuyGl7YLLsM99P115I4mYL3r/q8ZF/N
gW/1v9tqF8X8hgSD813LBjDfT2uu9A1LDFNEDeehnvS7dQQlu9XqgYpk+B8mQwm6VDG8IsTmo2KX
xMdGPQqrsGjsyZF4gnP/QDyNjegXXwAzoT5ltyGz5I+BhvVHmkkFjXBDrMNjudY5t//cCNSURlor
7vUVBrjz6X4IyVKPYFUltFgtjuk3aroYZe80mASfNRJjWUmEygMZtpdNTDSoZHg5oqU+sFqnPkGZ
aEUZK+JBxUV9o8DHWsatpV1iVkAJpSR0pQKXuuDGXQL02XdhDmlGhvmvzkXU3iwVXXqhmnaEuHXN
tDSsgb6VBMfEu4HR5OajFlgApdR5I/stBfDcbo+7lzoZmFYfhoAInB7JhADoiuDmCqW7++S8E6oX
xfFqCPpZB+E+mbOZDGvuLa757WUkguWqgFx61PcDbW7XOq5cBKZ8add5yw+FGKGEEE+Omyzex+aV
edB9usGVMrM7ax6EgGkS6efmVHJV00ymwZDS/rtLh+x4iLnPCzoJVbYX9hhsnlRxxUaGEUHVJQj1
u3ycXGqYZagLW6OwzQQ41fF6kE7bPShB0/6Byr4CJpsMKQIPjeyAtH9JXgmcIJyyc8HFlxRKYOYm
1xnX5Wh5r5COkTQnqXeEnrXxTWJKoqWuAHwFmGQHzoVcuKwNHjQdX6MmtH/pPYUXKSS46D3jNvx+
H+Co/+ql85WGfGMtECh7F4PNlEydzHvC52gtufqlxAwsu0xM9W0rW8xrmX2jZboxGJd1EY5gqye4
7GfwoNbj3/ap7XEv3j6RQr82BWlLsHs3y0OVKT86xlTVdqB+cUFIdtJ54qKvceKZ/1S8bh0iL79r
OqOGp7Z+I2w6VZ8ocbjN+1L8Et9alWnopA9wAE7YkpbKAJbh913cLtsncyJpc/w1Ksw5xEJ5fdlN
BH18X+75FD1rTOu/hOJFg0hpHQvxWPocGAZSW7jk3yxmLW6dQVc3DWGm9VwOM/PeBkmSIQ6zgrKe
WU2c92mSbaZ0ZsVLG8sOJj4TfBktIBvinhV8r6AdSFnmh61c0hHpcO2xijoPeI8o7IstzJ6qsUwB
CIrYu2EkkWi8VWEJZX7yDFiBXsa8AfwOxuTHfdvtRl+zt7ZYnXCFs2IvI9nqKQHv+ZKQl7XUD70P
SkCpgk6iNMnr48zeZrsPFVMV1f4pzxbh8AORz/FcjHLIJyxV5NEmIetYehfFnCDemZe7//Lnf9Js
F71ZZ6hL3zrIOY4KSGoD3A9Zj+GkHezjZyDGCZSKBHHUDXeVr9Cu8exz+FnPRxyL822/ZyBwtJOG
t6W6Rk1GK7ZOME4MSVtru0I+UUgiRm8/ryhuA38cU/tIuMkmGsb5K30SZQ5PKvLOuExQRvvsGVG1
+9q5p+/S+iotHPQptOQg+AB3aL2Y7plUeqcego2XYLeuDFKNUWcOdIblVS1uZZrD5AX6yl0Kwt+Y
AcLt2Tq3f4Kv9x95OkFtSVcwGWawihlMfiiJhIsDejqPs0ej9XbEjVbkAV7wbfC6xabONDWK/EW1
tpl2/sr64M2WiK5xsaFyUk3n3niV4uWE3V4XCtKm+1AQ68VSHL2fjVOQfrVp+yluAl1ny7wvQ9wy
Pn9SpTzcQD4NDAgg5lraiaFzsRsITMaYEcl2HY/oU/LyNR5Tb7MbH+ZsR+GnwjK2/VRxIBBBWmnS
av0wVTJWKiffjZIRk0jd74XERUE0AZZEwbMzxqgBhg4enPKSXsO31uiG/oBL48dZcANfS84omqKg
SCDJ9Ck5b8yGc3YUobBoURVFuvjmPEbOtgOTAdR8zWEu572aZk/ag0jeG6UZdPuWQ/RVA743X9nH
vPdr5geiU0qEuTz/8tjr75To8FZDngpCAOCziJ1qbpu0XPIgNW2hlnfLX/BM2R0i+viQ94rMS8wk
sYW7KMDrFz2VQbcCmuIauXDs6NQUIdKnP6FyiyPUkg8+ca+zkKTyQV1ar0jFladiy+737WiVDwOb
0NPQ6NB0JMKxxQ3MI12SbltOeCJ5iZT/G5FY1GH4/kOv3YhrkAMT7v0QSVD/pxtC+nW+y/E2ZRoO
7K9UAjDwNuBvmsV7PbS4Qhfsd60/lFL/lG8uI19VQBy4QjwRrRa5eJXsDR/r42TpdZ55ikRJcLMC
tiQKdXs+E66thQhWOKHrCyBjEEheDfDd9T8+Fe0NrlG9RdKh765PqEJY1Cn855ZCYLtOD2/oX3VH
3gdcTlQaqCEebtEW7gFJwjw9cLNtSmCQtfy6oKT3sZLM7bZ7lkzwqaevKm+3dDsX+1aXr17L/Nnv
XnyzigA6MYbN+JLdDsdpmcepSNkFNZvkaGD71NP+dxzuXo/s6fhFOxo43il34+QIRHA9MCqzLXMr
SLwmioqJk94IxPvGRRxhXeBecsFD9JF+JvHTHTprfQv79M4TXW6KkkEOU1+OrXjZJJDzYU9yc+rX
UBMP2vYMC02yl18DA6RQ9iKpLFFLD8tlD/HzdczutEXybAl3GbOUknAaWkZGfvXUc4V+asxq5lFk
cheKsAMMAYjpZTnPlM0K7chjacmkY71AWJ8kQ7fpoVTIPCXhjWofRZjKo4yLnTIkdx6p+BvvGQ+4
1g0YOjdvzjtBS873MaKrrBAfZ35PEWbeP122nwxzbMkV31q0nw1p2bF+cQmIppO8a/Lr0JYqSUQJ
7gD+61Rned4xtef4BnAyv4gQGtQ03mP2q+n2fSKEfhKkDujWACu4vLwov7jIIZ7N5OyGPtvLSAT6
I0TOBT/a/bWFECexKLb8fdTL0lS2MNdG2EIgwuDrN/N6vZONA/8srq6uVxmyczgm8bssHckkSqKO
TPz/z3IR8JYYYi2EWPB1i+pxna6jTLbiIQ3Lrf2zWul1Rwrvfh0spnFCejgHBbRFueSMDiDOHnXI
mYle0jSfPi7ixac4Q/y3gyb6ZTLtT7NIrbLfUs7WNKcMt2+t77dqsInJpnqaIrxBD8iresbPUn5z
YLZ1EIY3QGTxHJterax9aeskGGNL7pogu5VPOrwCJV9Er9pM0joQkI465uPmkQsLLpPTN6wu6Ueu
9H674DQg4OgqgM9LLvkowZf4qUCe2MNlTGaECqDWvThX3KSuPBLTCAye/jLDSTIG9cHo68tqXEU7
MLvEbUc5ddh35vb7to3dii6h0PTH5kUZrpTLOp1hUPF/M3icy68cmhV3OeBij2XKL4bBvFzdQCkM
DsOoqPdHEfhuRSc/WF7/m/WtLLd1bUivqT7Ff9GbdiATWwSP8BeC5uSekguzOCYEiNCQx/Il8B77
3stRiLkEzX/ym8v/XuS6IUGqbU2R4zPBBqz+jdb8SMdWChwy7XJ2+dtII/lL4vl5ZZP7kenIuE6q
i1OC0yY6xUo6oCs5B+XctOsR/PJb+VcNHUvuKbol3wJRdqs7iMguolxtavf7gbWiyYb+/TzLw5sp
3KGV7UqTMk6V9TYkPvdNETCSX5hW1gcE1+oqBcayAm31mNnzMIktr98Uuo2W7qiA42pRz+fCzcJM
Hly9w0mrwNp9yeFhl3s0XmhVgasYp27NccZ051/OBHrv4LEpiAQpzxbRYsnCtMO7tpMzUIj7a6jb
J0+0RQWF3t0gmiST8UYl3nYrHiu/BQmb4sbDY201WXYk7yd9uVKr6uMKFtFrLW67msOUmRjff9Yw
iNep5gN2B4DuO26FUy5GPPXu92F43SK7I9QootqqorSKvg1AlEQ8lCkvv/Eu6Ki0gx67xIN+QH2r
L1PzLfu7bQoJZqNZPR0lVdZIK55FKDfFYNqiRd+WqDcf+syaUNzA1t+Y/6ngKh1PrGibSizUzVaX
6rngUQ65vZSazzMwRb6Cj6K9sIODjogDFN0fYu9J8rI9Kri4C+HwpxOCXy451nFrncDnv7qJgFGy
0pvwufRhMcZ1PIOYR/0ZgwBOwoC0ClzOiVEpB+2mKd12Fbs4Srufjcr7ac104UKlXURmC/lbhcZu
HN0kgNAnvQ3Qv/W3urEvspki257bRdgrUGIxYViAxt8KZvw06OaXvrX2Ax6ArJfjtqi3+wCt6Xsu
jvmr05gO8GHlXACJ/TsGLdCq6Uuk4eqHZ3eQ7znJLbdTGpp8fGB7JQBix+ZrfBppBk2CLnaJRb+T
WXML/vEgUZ7lwDv9BQ3KJo6wicyy1XoFRJTXLr96XyqdzXNqnu/gnp0dBuxg8AmJjxWJu+0wL51X
oPrvBJt/YJXmMcNO+03OjCk6izsUMVmhiLmhioDPvUvrbo6I417NYxg8iEljTyfvmS6DBMWtRpXG
mBjUxGaZ9TAAL2Q8BaA2R7/a9u2TTljriguqjTWN//xoYFmrv+oczi8JPDpTUfSNdAFxqAH3KDkC
GJtKt+O7eOyGYU+5gry+GuCeKCD2G1t3ZqUhFBErM/9ebOP6ZjQAmF5rxmDrVUD+i5KU7S4bRg0o
X5Ncj89XnL4fa0XdAdWXivlGbNK44iv+F6FKD7/lPTkEJ0OaykpO7VpFw9Ef4FEPJV5z0xezTkvp
QKTyvEe7datygZ8iEbXHl9ei0/z/lqFtClE8XwFLfJh1I+b5jhDxawxNAfYHfqcKE76uI4GljRD7
HqhwWzaqaWOVlTJj0wNDBzjMCmGSt3I4CygQh7CR3SUjDxlOLlZMS0sDTCTUYyPnsKSvS3xKaFU8
sM17HSrzLxF8uvZfcTJCZNTc2rZ+ngHBUwzeJXQd+GpCAPTC/FWZ6kEp06TVZwoZdAU/TQp6FYn+
V3rjCCpsDiv+/dLWiFNE0Fs8CE8PJ7BKYriDZqzmYSSIfwKg5EqnzQ6qlP9I2+psauCDcSC4/zrh
gQC672LyDr7nWoSM3+JhzF1syJXCym+UqGBPfxW6z2cajpcDL7nEBZOMaaY2f3OhE7yn0lLpReQO
7d/OqIMDX4QLXLoSkOXZaOf8yeQKjsCqEHmqVq7ATy7YCf5+L07Sp7e5Ka2NZZ+s5zbsiLIOfZQD
54GSj/+zSNfX/fXPcsAOwueePvj3xZowZFrNRUcmMR9Mcc/IhYnQNO+6yCQrQF0sqIAJ1meNNOgL
jVR5dGQivuEGirUUUxmE94xb/K4SvxN3BFS8cpIgqUNimD8PnC0mfg9uA1fEZKxW2PO4ozgMJvuG
whrBj+gtjN/juMQULBWyLnX2p82AifrAq0N/4FvQFpbSls+4KSXyHurklTKeuUNdPUrk9jTbG1ji
QGd1BlU9Q6nqA/+8/nzbYS934U4813D87KQ4506dNZLk/jgJY8PtdPQXvNNJWqXhqJM1VZIzXGUR
6rVrVphVU15ClU4hzL9HoaHplPweLaKxWOiqoArW41xU6yDpNmdXSQ7Hd6d+qm2ryKni4Wwm5isD
IDUS/O3pSrimyrl6zvzPpy/wI6WNpYy13LGihdSLR7AqaNPl37xYtzV+xc3acwwQNjFaCyGrxDZk
ausAOCdEXa81HetZY3qFYL3FTqgE2KgCDjT5+H31PSgo/lab4DsncYvHokfzq10RbENmGgzqWU66
KQ2hI37PhXcU0zhRPprs9lgh3+YUFtULKlaLVKee+BywCXAS32YEwSF0OH6IwilzyuySudSGyNPK
3r2r/2HJWKLd/1f8S5oBKrHZ6fxlryyyjlTyWUo9P2mGp9XagiJJkbdXKJHzdnZJmsYSU4DxztMH
upQ/HgM1e3v9J+ftfifo/RTxeEJ10ZonudtcBz8NaAXW8ofiPHHH8OtiCrdkcCMuwkATpMruoOKC
3P2p0k3eN27/r6crN8x8IOwNOoVwgyrgL40OmhtoqZwqfy2Se8QSUEiIrSMWZOS0Yi01gTbisMCU
wa7LpWAmpydb5NwcYxzX9taS6P5uNOVup9S7qq4S74DbWMK4IaPiYURVgBLabb7X6E+ngyWThvkc
UrvHaAAra8hudqwrfUF1bwgsvLKL6V/crKRvsh4yMWkF9cBfictlIK2Js1GHVOuEZUp+Q+UR7fTS
Twqb0a2iwjF52KQshLnCoghcIYeBoDDuRhEGySJBOkvbqcthR7S83dYjHEhonuumJDqcNJpqPnjs
OSLL2OSLTFu5PoGeN27Cplins2/vdxouNrQYLJ+vRs46mH3mFQqk2jwTt1Sx5iIwYOlXyaJQlUxN
8myAGThL9JnHsR9vM6Q3i9RWZjkQrdBV/igFwkapcDaL1IWAC8BunPN+Sn+CbOGoLZVWcC8joWbh
FoBA7JRGuZQyyC33KrcAh1sHiWxXU9EmFOo/f1vB3ClDPB6ol2rVBo/LzE5PagGZPs8QfEUBu4J9
NK4KXLIhK3B+ZwHwuUEbgKylWzIVsOGVSo9F4iaHqFd+GXH1Q8BwgL9V8IXKDl9DgNe+O66muDt0
7Pt/C3lSmqGfPsOzDpUdby58RkasItYEgA3WNAPmaPacozZFwKmipsns7bSG5YZXLo1qXShuYulf
HC09AIoqvWNZT4IVdBubk20v21EzC8z40gHJHs6Hd4NigY3P3tSNx5xmql6YZCUQMZuadpU/HTsM
St3314XlwNKhyWUphTO39Of6f8dXp9gq5mujmbOX8JMtNBWswlHr4jCDx1+Vie7rMLfLzToL/0Wg
4TWAWnC44KKcAcJlP6t4xPJ6Tf2KzzvXZY2Y4LamVq9DRTIgkVm9kp58ytOS9K6NuWnV4wE/Xc9H
+ZJr4Fr4PpyIBCmbsW56FxxRQhfN0kLOHjkeh0Oro5eG/nLQ8j9vespWB5GsHFQwlLFZYGbkB0Ey
2Uxzv6fZoEWBtd1cmqe7vnJLqgYoaN5NabH4tsxdwgx6YISWgAZNiYhq90QGfndqMAcAm13Er21k
s/jmeml6EOr+Px7X3B+8KekdNgcaqyOTSzwG2/ExRSUDEcKX9giIoDoMgvLqu6bOGFYCG11By47J
IF6KkbQm4EG98OOyB8GQYjgK4AYOLkNhCOnzLz051aBtc1tH2jAzxpvfiOncLrjM3t9kXMTQJFiM
bey+1Fp/skMa4wLqIJEVGirzzULoEX3Cc4X/fGLkLlfeediMm//hF0Lnc/lUjeH6G1g+yDT4HwLB
w42zFoX6Wtk6meCDT0oUW6ZpWvNk5XUzS8Kj73fzaGPqztiicDUk31Nt6QxkkFE+tVZKbwO1hWDM
Itf/mM51DLyGHGEdRU/gO4QYwBxlNZISCsd09XpW8JN5Xp35wyAhGxDuB/ZO60uXvzCG8IvAJCuJ
EPqFMO4PGHOjUrQJvblOVZtS6AjJdeVsRFTSIPB/gqSf8nEbRS7fGYS8A57ArWXScjvtw6HejJnG
70EiWm3fpZQSaxf3YDq6tR1gK3X7fkQs+Yd62WzZOwCKjXJP57uALtv0eFIoMSLfn2wZ7HWpO2tp
rFn5V6v92dRflUoIFf3jUwRLlmwfq7/UQCxFEbzB+Vho4BVjYJmUycHUF4keLfNhtgo6G7DbiEnj
0UjkdEC8+spM1LuP+3xXhGomWvXQQLx3UKPYqdEAiM9hwbrHHDr4skr8EgyPLFsyHQ3pVwjVh2u9
TE4hFGxEThMsynSWkXroOzpQVczN7TZnQ2+jWPnyZVyi0hwQo4khu5IkkvJbX0TqMfif5larwTgP
DUj6M5/OMEZMCTZ/cTGqrJQL/Wmi21gTlS0J6cOsav9dmQQYwW9uimQouKrCXIEJG8X1m6cI9aM8
x1vOwnRFXN8YgFvlyTrfU3JLzV3Rx387Xl4If+qZc11JLdv+dqLMLh20+yccZixS4HcZo5gZ0ul6
IXGr/mjyKgH3L1b0oPCEivJt/s/T54FqKVLrSCMfWNxzpdFZfL7tlIHxYTo6sTLiQx/cvwJwUM42
NSGyz3MN1smAhmNdNsm9PbWV3HoYLfZDV1fbzoHiCNaBrRNIN1rziPKdlmdvDfBxeMgKFbifcFTt
Tv/Zu1K6M1RG92frGTOb3Y/2klvWrPX+TgahtpyIkEDwQmgPR92kkspeJL9QZJONTmCsYJc/kvpL
/WezeCfw5WCOstHTrCXXxBgNXm8O0yPUYkR9n3a6OQ7qq+MiRn16J2ZiNJvjnesS9vI7ly/QXvUJ
TeOLuaQMctFxlEluB5j2phZT+p13hC31SfwabfWCn25GNY8G9aWRq9GlEDwUX2XDaQhaS32RG9Th
hG3E5H1XOIT4pN66zWQ5y7b+n5WxjYt9fndknN043kX41hmnZ8OG4Pen8pqUTcWwMUh+2LFUhmxN
UZ1B+vUzQMuLxYhc4Fhz91O/pJ5MXnM1z4w8c//x3yIaBsgyGeda2IZzTHlv+xnKIEMSMBucpf7F
t7J3ejvqmlULAAGtrg5zl/ZBYq2dwKEclnV3xga8Otpmpu3XGu9+ldd88c2L7JDCHHa3xEUVNfcV
xhI9HntR9w0y0MjrjVF7q7rLNvsa1K85DntpgHlkWiIi1A6ngHRkP79HSFGaVGEz81np7nvHoKzm
SkwOzb0ccNZMtHwBoy3dAgtGI0d7pIGLAH1cs4U2Al11CVQ+/+PUbtdjXeH+53YY0NlUKuDpUh2Y
nl0xOGjnEDMsMmu3AkNvZ3OUYRIxfFbBWdpyV2nAGZ1cKqgq8/mRart/Eg56OIz2bGdT7Y09H/rO
aWfXPlkoJoKj5Sxo+GqiCRJVLed5hx4EznGPeQSgzGWAadHtnqKdvV4/P+ska+V0sgciAh/va+nf
qoToRu83Exf/Me4G6ywQFs/XdPZviOf/x4ha4J813M4IwYzxAFAxzuUaJmN85SnmbTmHKm3tLqDJ
UxrXQA5E8qCV+gnSFOMp/xOk+fIyMhhE5WcwU4ZXcSIDQhR5IR+sOlLdLS/Wdgci+z7aIma878db
5Sms23ZJRoulsMHJ2jNzH+09O/S6TICFcG7o1iZHbyLN25B4xDwe28BTEE7jx0Fdzx4EN8CvieY6
2WUxxjb6uh+shoGlRsKdEAMgar1Wt1hxUPHAJ5KlBBwjvz37IC3roz1HT/8tbtR4ZiGgZSZo5JLT
qDWAMa2HSR2hRJJpbTXed9la5TBAxOVd1Th1Y94HQ+euE6v56BO5F+a1EuGx35x5UoojjI/QlklS
/W9In2Mk1BdlejOQGLSFX8tdBh+QV+VwuT1D9veT4QPUclRpQviWi08ruVTpoBqUwNDx7zFBw9r+
r5WFjgcd6PEhUYfdSgXKQiYw9dhqugK9Jsqquu7BGFq8pwh2LswinymjJ0NbBh5kAcCh3AtR+/zJ
+h1lvGGYO7in1nPxImvtOGhduV6AcaCO/Jm2OOmZbJVSUClwhNEJZ4zOrOUrCU5CGbvjIiG/WIAp
Jmz7JKgrXUBD7jJm+s5DVPtpoD1AeA4MnWEs6Dmm65Ye4JHFITL1UhChLQb2GTX+i7514y4ccPk+
rKtNxYgrjKtJcfwmphDeYEw2TAXd/2Drd1OAH5astod/m6drnCI4ZqY5BjUQ0cjorQSpYpt71Taf
525yUCSVdoVkwJhJR1VM/4THm3nsRtxLrnxqVnXSIWQdB2XxB8PPsoS2PLOuTawDmyiPUUP16WIF
C1LRhuuxRJp6Udo3elUZfZgtWv1lqwD8Tx+eu+zEErsyJY+JpyAsQDgy4tXAPQDcy1XIDBZQttyO
qJsgy2SiQQBnqYc32FlB7YZcKPpTzGVdymHhZmnWHyUQ3Q9D35JPBtHC8NGVxv4wbLmwAgJ8nQKy
XgjbdrYpUoibaBLfBjtgqisEwyGVsq3hpE2ZW2pcaXoxFASzkbSEV+d9LmN/H4C/4ZiNqziG5f5c
mN1yb0sftLwFUoUope/0qYMFlihgk7x+xBt+FQUCsr0yfJ0KsZY9AKH7n3rv2xNG7zuUwv/1hPGA
UzcvDgk1+7dpAlQmjXoNUvC2/Ubka9IyET71ZonPFwEChoNeM+wS5gx67iN6eSf4KXd3m26Vl4nn
hL6ToXJoq3mZUXox2AT6WB2vioAuKXlrRE26vWE7ahUJqNr2bHMloYyCXB8tAjaM02oftXS3qoD4
MM0FRm1+zttcx8Au0UVelgeml1uRkn+LXNYN+EGrtV8l990ZnsALlAebKoo3CYXWCfFr1MHJyEDq
0xqJvnTCCFJAM4/YG4MYElXm55ZK3FHRzWU2sN/Ut93Fv8HIMdeNmfyA1jHwq+BYTXW8Q0+Cf9bW
1kMGwK9P9YNorOxVApdba9m9r3Nx5ECgeLM6FRlZLG1E+bs6MktDKWnTFJMvxzf4imUCG+DBiVXw
5G4d2PhSqctxSR9761F/ddvn2aEW1f24qXcESmZ8OTxqlJL+DLW0HHpYBHIZIa6tx+Ds1ceZ2wj7
RMxfxekgY/ZuTSUCMJLQmYT5N928o2SW9XJX67JZ0KM4EqyMQro8Gb9X6ZB/1v+0yIssRofHPltb
Jysef+Itk3V+dfUkH0qHlfYs4l9Is/ZTOc6mO9WndF+/RaPtjUa3PTcStC7TA0+z5gkGwJhSISyt
6mXCW+y1f2bJrfCODlfvGD1GZoLb8jZyOPwcUpvitsH8hZP3Qhdt/vz3L6aZQJV3ABzK3iVzYmnR
Ence6LbqvhwrKHSz72Dt+Ocw+uIdeF9zMEShQPR4OXlhHRBHY/aMMWfXdpdIrtsFGHL4loUNfP50
Gr9RMHgpqrdRip1aeclD6A1kXLNZjxecnfMKxp39ncQxtF14Yux4YgwV/zWp09HpcBuO62vfe4EM
mOUwH+f8EEbteulznHmQGR6kVr+DTneI2BMswBrQOP+w65xcUCqhrU2r+ht3Tgppr5szrLQ6jwak
8Jh0lEMTMYQpXYxP23yh/VAjS6DprquxaPzDOQttHDibI+eFNmy7OE0fsbmYPk+gcaEJNyOiufYj
rsgxNenRjOhtVgR4Dhw0qsBrZc0V3a8jIvRZgpBNW1dC1TQdunl9kJfLYwRTjlqOyl5PnmFbvvMz
pLlpefQO1O6T7/3VKBYgEaUKZimamkaxU8By7pxRwWNs9HBkKrVQwQo2THleXSHn/LF2tulimecS
4Dub0C83c5Q6HN4NCi6dcri/5EBiMGZUitXK8+kO5ShKAVUUvJZVrcckSEvW5rhfdByuNud0ZgMx
l/P3G9mPM4HLG2XMwZJm2akTPVlS1CsEBMjjhKa9a6Rj6MMIHt7j/kkntl0+yE4UVF3WSDyuF7vM
foIhusYwzpwuW7M+wPkxrEM4FNIWNmE9I3hTsSGxme1zuAlatHSbd78/zuScDooVCHMbAt0twPzq
47Kl19XQ1DhXjy1EKwO91Z2U86d5SYC08MpjDXH8f7nQAAOtSauL0OXmeOPca3J0VVvnxai9mqxv
3r/HVbi94m43Mcw15Erazd9sCrAisn/GgdUepbTgeig9wMb/xPSQ1XWtpBYb3RkYdTweniPVr83p
+cHazhZexT9rTdnoNWc40IWu7zHgcjpe0cISAMyuad6Si6IQCM868DKWYWm8fvTbghsfhMQQD3Sb
/19orpuhb3/pcLv5ebfl+rh1iqxCA9t7qKllHBV2rCVxvdfpY7qH254yv2s6gav8BNdffm2KVUp3
5HZFTy3/2nV6IRw/D3aMqk/BJLs81hpTpcnsAzIaibB6CcXjD5E7itxD6Kex6WQCZx/WsLISiKhC
Z5a4wuaJFtrvX/Day44a9ntJFsYEU8ZKqXZerXfx/J5lJr6+2q1303UnvfDcCMOV5mcDhTNH2IrC
gKsIaMhcC2CBVOGxCRwziDAs1rebM+w91BlDcExDMrB7V091w9kR3wWIgF1d814HtDE+ecU+KYpc
YkKOwS4PuBhK8hN5pObj29T3Z+R7zVDkY7K0pwP/wbGvPpwWUoslkNUz+gQ1bn7z7/NLiy92zQoj
ZvHAuWLMYYRLlg7VvOOvUvemy+v01AjkRBTc73TLpKzM7dxRPwo27qEOo0n4fT6u9pQXPTxXcoq+
EzFiY8iQRoGLaSKDFQKJhPU7C2nFzX2FuM0Ht5l+T+2+NaUvI7r/lfiDbbf1C+JHe5ivZS/yJgyf
LiVn6z9ktGigQbR1XqF1KarWdvUckYpYIA9GIKX0PjxaXDaA1a/4iDyUqAGcGIOfjELFSquA86S6
0T8NEsS7PIM5QA50C59r/Ikh3fJ5dRxh8aP24pMLAcfPz82B41DMpE428QGQqdzhFYkZace0j1JW
uqwkCwdeyfQlLI4uLzsRCO7hb+vphluiiiSqC3Avcx6r5p29fpjNO/DuZi3U81cQzYO++RFkMZO6
pHiRi8hPZWgoSqo6Y5c+aTmZhoLLJ8TGMNV9kKJwTmyqJO/tvd4Oyh2mnUiK1iHCXN78uhgpy2yY
vgFUssxHhCkrVpeoLf4ZntCc4itFZaPCwbbQOL21rXYM/XvxkpoE1oDSswPRqaKBRDITS1ONbSaE
Zk2mE2Z1deUqg/PrE8q+CJx35ChKC1iPIfgZiyENTFc+L4yZniaS3zY3RmXNvhGD44Qs0D23ufnw
SKmGpaIAmNm4pvFrQk01UQqQRmmZxa+y8r9E+vHfxo0ttEAKTCkHv4+44UhmDMuRUzEIyzxPZBsO
98a3IumUibGPZq7IxNf3THd4exEKpjmp0jPoF19PVrM2/AsOtizFQBM+DkwpQUfEm09edC5+6kk9
t0l7af0TL5Ma/I0jmOZnmjxSnxr0KkRZtVXWVtd58AXq1NI2CeQOIfXVFftpM/ZOX2Z636FTHfu2
MIbFGCR9QfX/RIyqZzJpjyGBAUT22ihnKAfZG5aPSUlnS2mXWo/dMJcIYqCJHf87hV4YP/dcKhga
duOEBsOb+wB0z1xk2UjCvyCy0uYv1AejpYerjIKC96dAz7uYj62oTrSP38dPkepvWuhP9J8dIBv9
FbhOpglb+kq6OYdSexSoPz3GiMgv8JfyaCjp5tzzISdNcOv47G7TdZnv+zNNj7d+nK/kJLv1Y67O
VK3PvabWvVdv0plDbizdaxDlr6mihXgCzpWgpACa1H3eSm/KCCnEJDNw+EOgJmJJml7I9jkWw9Ri
WDDSuS2EFMy8niCZPt59Ljh7XHAuv8npF3Av8Ig2BAklNV7z6FMUSTJHFbwESCHoidrsHGFDwqI4
2Hm09Zz8yX41iqzs2JxS88u19A1YAhDRbakCP+pVUKoQJvg4L7fH1pXHUv53PCQjE+VY98r1GX2f
4sWHxbOdWY28lF1nWtf1K9KE/M9zY5TMTLQ2ccam+isjx967Ch24eHNfql/hpexX0eMhYbaHtrVk
2eibJBQeoHHpoime134csIwOsYvXARimqnIT2a3QBZR0hr3L031+PS1PZxaCvpFn9TDD4N21bKcQ
BmBQeYURFGHXNdHin2DS9pykpvDQSnNs1dnz2/dSa0uKb2M3bImjGx4csr7q02YYgllHgA7wygKy
af4k4iErQ7ERIjkEAnxFCjBmt4XTDebGkMSdE+Yaha7cIM64xkcsJF5WPx4Hh/JRRB0rSh7Kn071
t9VXmQ+k6PHfibsUzsLH40v8182135J5hpMTrN2LUM2QWU6BeOD+I8/jmiS5FOQTLDU/Wal7hsIp
oKRXXDocF3FlpsisSFEuLBdGcDtWXzBUyJXwvXcY0FtpPkUhAl+xSnx5O9q/KWPbZXVeV8TkI4MU
BxCeiReT+rbCkHNcWlI/L5NGT7QTBgs4nnj/8WkTECoFU+pIBKdNYMCkU0tcX+IUEQIUn9MD9MSI
KuFoe0i3mVWDq2V5VzZseNzlq84rU5Yd7HOXTdImz1jB9b4FTDajcq4p4TGRGflt9AudkcdKewhM
QHU9ic2yjLgjnmQS7qoIcfW1JRk4Feq85ZSBKK8R9mbyA3w1Hhts8DVChbPZuR2zJfQCbxC1CPYF
BQHjW2AgpGt8HZu5O61p3AQYuYM8RKkxo2xlnNmd7PNni9p8RMt4WkSGcGfiuop30p4EPY90gXh3
nQ4dd2LQFt18/DeD1f11ARb2bnNHDSGsFJBSz/KKoouT84r9talhN+w3BZllyB1pRZXWVkhBZpn8
fdrTKUcickdLkfRGkQVxFWtf9ARd6+0mu7dHjIn80cqyyZHfot5Ft7KBfh/HVkf3L5GjWxElTZCK
L9z0ZojnSswoVyaDiZ0XttRTGTrO5zKmSnGv6RK2UeiMWDZ3Id55HGSWyOyTT737YG2CUrWBr8DN
gPze9XPyig4gHkwSOVkb0gHAmZyuPw8NICoqznaXX1Mc0FwMXJYucY0mz9zjqmDiIhpIyz4hujLX
WPwFX7IQrZQq6/z29FAQTkq+n+slkE3k4+vVvx1nPvXMBphu6Rr4EkcEh8TLCw1IW3iwcy9CutNa
7vYRwnq68zP8tcPZmTZjkZDa3tYHo9eGJXesw/y4T9KnFZbqBTIPOfP5cN8Ouq4qR52A90QbKjqI
gJpE8Qskv/13Tg3LTewRFQ/S3Qz2DX8fnxFO0ZZrsIzP5GkfD7tWX6Ad8HxFHG2rlihLOJllVQ7n
HwjeJzhCHLGudPKBOeWKDs3M5MRXqu/kse8Ym7xDTKCu3HxnJXX1y14tK+W/tDDmudq/G88R1+lf
DFQgrUDLs6iP6txKAezC376Ei7ikvyqeiutUP6chwyVj0WLPV1ebT0XPU9VAIPPRxoxQ0TYZXoBP
aVuiMSZByAaXwBeDBKwF8OJh01HmZFxR37AseU70CrqXPQatDcmjxaMOKsbO99MYwTqwQsmFa6e+
DiLv68W9AyuHmmlBXcJiT8Cd/5miIIlZqheF42uwyJtlotkYg35Lh9CeUt0F+Ba45QvidKsgKAZM
8i8EasEdhN22mT48geAlOf3lUx9FHk9vokTQmjzqo31nSwLeCvgJvUm3Nd1KXKEKR6OMmoL3F0+B
WbukDRmBdaUmSZdI7KkA2gg79WEA0Q2Z9sWAJm1qPYFzyrhfepGJTuIaPRE+ly4QSziSDz5+vRaG
4ag/bv9OZIabT52NrlRnUiqLvBrEZpot/MKsPSdEhNEymz4f7xnImJ2k2Q3/eq/q18DZ8bARSna3
fc3dLhNljXNHmFlSmAP2S6oY5nfWD2PeSUOSi77sHifkOLCqlDJVjOcLq8CtEeLYOUp3IG/BISlR
s7R52708BcwA/+eVgi83LqAcvtp7/Uo88EXw8FwyCLerBspSJBKJNNIxrftoNqZEljUgPm9BK2St
PDL9RYkhED95v0XsmfR1jkIIM0YL8u9CMU8mmIlKN1Kp6U4pmDazaXalpzb3aJ4lvH4xYo+FQiVv
yt6SR2J4z2KuMYuy24W8qNv62G3JWMhUjz/3rtQ3mpKyAcjRtjg3Pk6Ye0tVaIj1HAVIixtqVcTo
+vefCKL8EaHVJFkjycS/mqjbTgzTWc2LfVB+xKaQ80c9lxCNv9Krm0y+txW36RZXb1j7rU9nCh3a
pGQyt63/O0wmyNTwbhr2YsF0f0A19v7pbX4oXq6U6WKkOMaZg0FntdR1VoR+sQr2c6Vur88ZT4jU
s9ywyuUCvqq3c5iyYxrEie6qJfevaaGhExzhySHjmswN942gcbuzLYFnDDrTua9hEyEYkE7DGc67
CGtHyT7HU1Y/BNRNQyt/IqiSBRSFTjrC9QCLdOx1tKdeD73YMej8YpGms8sjve/7Wy2tspgWgGP8
R2vi5LbQgHTeelTjWxqbJjz0OXJ2IU3Uh/C3EtnIwkqZ2b+0c0ScUywo4PmgZdjRzcu96mwMcQso
+x7J7hER/qEupa3F/D3tJdtBZqah9iwnomISKE8xB+DwkbLGBwI7h4QgOx7BBpJNkNtESrZ1E64D
POgHSAwtWCyewHATiybvl1b02IvJ8b6kSY87pBEcBC4pPonRqa7kgsnCgeUpqgKl5JGxJVvXON6O
V+9lDzeqyGZh+Wd5EKf9VK6SyPDQjruWndisyoyn9mH0pJAdxkvmv0axzwnvx/xRgjwKDEMhZS2v
vgdbIZKRZcWXgC9Wxm7DbUa2J1FPvU+mRQkWxRsY/S02KsMWigACDvnXwWdyTJ149j9ISf5ALOe8
QzW2u7juffxTnBYrH6LRs26Y13B5WlKNmoC6N1MuWVaes7yiQ9kGyS0usm1lAnW7eoKZRsMZ//j3
qL0SO8aFs8eFW+5WLabTJ4zrHd7mMYqq4vvmOxrDEyMkYeIUCwhCQY0YbZ8TjOX7wqgsn3YbE1sZ
jsqSBXOi67u6pk9QCfCR36xkXa+g9LZIJ1e+t1++/fR8pipLEb5h6pqxFdMWR1td6yj6ZMm7ew4g
Ipu7+eXyMmATPMkuPWaymYPjp8kulfRA9P8/1S36G51btyGRR4GAvKZg+qsCeg6hHu68o51z4+B7
pCVgcMqhiA5WZ39LiSikeZwKTfXdSuRrm6tlz9h/ZC7Zl8OoJQyXTTv20WIK0IKAiaX0IBYxnDR+
N4bXIqUpPxXc/DBwTnAYecc55eRGi2qkC2dx7Ha/PMkGPjsa6EhSJ3qLp/bBdVczfxbOhKAMRvKK
46bVkvcu/Dbgum4d2USx2bQpGTmHDY3u58G6n5nGwFb1IuPQ/fIy4HzR6+xPoPpiPBaMChRdGcB4
aH45OQc5C5yZ8Xq2wHHlrAzCWqmIRMYp8CrO4W0ud6ChD8qDfWdHk0VPXUfCOCsUi8FDI+c+pZdW
79UvYSVw2kx7EaB3O8rUbosT3lgN7HruHdo8B/YEJxngI/f1dRm2XHu70clYByr7o3COfXWFhuSo
LgCr3w24FSkbkeddKSDVzjKRRfGu0kwVmF1rR6FGJdc5XeYXIJcF2VXVQb0I6h6gksG+K4pnEn6X
rtk60utzMJSadF1x2p4fazETKxKYbu6xlzIkW7NFzzk0LNtd3/w3/CRuXQhjgJftqoZK5QNcWwJ0
bcAXcIQR8boAbV76jgPXytUE6yXqAGblCrzMT5ro7Y1E31gS0dfukzSyDPhgvpYyuctx+KjU58Ny
827Bo3Rl+0lDXkeMtxV4S/JqtxaacVBY5vUyodT6UQI5hsFwmiIViWe2Fsj0ibM+x5IWfA4UtzgW
XkaHvfPsRCNeqzDHbuN9iQuAjIL93p9INjtKRTqZS6zO7ik1jqFoArqG4xA0m6rkOXtGKUk3zQCf
NuFPEbgiCyQrYf3VQ97EOrzAlsAbg/bM4XO+O3lRpROcEeF6wErb4olvX9JcplkOLnFvsDiXBk2A
ct0OcsqdMCTEsefOAvACbchpkZtPFbF3I7c2ETZhd+kzw/v+KQ7zFOC4QR8ym+J7gkLWyYrWca4G
X945wadk3Yg3n1mJQqbkyxsnksD6iMpa3XqR9ieR8HX4rTk3KbgCD7m3+sSu+9YF3O7jqzXgpDmI
5cy1Vt/syTmsJx8xvtRGByFN8A+FaEfqM84EHxltBxczrpT5EAdUk1s4OG6ethMvL/kuswyrvDmz
7EvggdKAE3Kl4TvWjWG5l9yQkyOl4jUb26QjpGobV4dl09YAJ+BMCIeOWMHba0PvTqoweely9+ny
DjIXxuVwFriJsDZuwjb6MoWGmI+7tLFcKH27P7fw6kWfDL92lZguYgtWJbwjC59o3ihhak7fdVWL
6hQU0vwuYzaRSGiVI6Yxiu+SvRQ/pyfUa3Hz/719MDJnKm9fzX5EkmkP2CFeaM7WiXcPjcElcf//
JPZLbBcHmV4ytBBe0MvwpL15H6lr1A2bi6ySUqqt8OAwdviEuPyX0DMhy0M0JFRB00JykA9TASgu
u7CxUphZo9de+UwT8f3IsRQFBjs3SrD5FgeI7rvYHcgn/R4bTcSptyeTFmeExkXZFOpo8dUq2Ekg
l1DDa8ZHWyBJYjnYB4+0eFkqhof6cv3JULP6C2dNW5fgnqmWJm5dpQP+qYLv/EQ95gnitJlUUnii
+rBx7Y/vksSmkLE5VXeQqCQoBl72abPnqyBvpq4Y29VmIbkR4Pb5rjY2V7WFsh7YnijAJCdQndMf
5k0hxlAagyTd9uM+5S9n6rSS+zxrD8eJj0ObypcBhwqd88Jy/zBezQ+xXxzyhuEx+S06qD9Vj9Hs
lsZK8edVlrUsgc66qa6JpzwUwgs2u3kAHs4876o5jiUUu9Xsrc0YQ52R4xGxETrn4GXNnh2v/a1o
aqR/VxRK3eS+ChFZhkSoUlbr9aAAHgzF0x1R9by4YHYfday+Pq/+i9cLZ1jYZk6F+MDwD9fnPJPB
sBJZ8d7FmwwL+EV4N/JVLdKhpqXuHdwwrdWvsC2jaPPF1ze2D5ONE9BH2kBGwMCckPo+VK5qMhnB
I7JMSgPQrKO8D6Tdl/LmjmuiPBHxOW5ThKz+gV3vZikYcKWAGR8xQLNSUxVmjdy6DmNFftqjL9/L
omIaE0omQ9415BlHtZK9HaHTWrJ/MWSKcp4Cb34UnlxBDtUFYs0izZzoK2Offx/ZmGpfRtrLqtWp
Me1uHYt0eTq7KosN202z+ASNVTPKNPWX6qtW4RbKaHzPldOj+W0bOZN1YIIqiqkceZ/xO7Gm+U7k
H8wqdSdSSLCJlE3Qth+KogRQIgDo2C3eVuGyfi96RKeLuyPVyMOKxVjQACJ213sslt1zAYx81F1l
5FxO/tKwjyDhbPrfBbKZ2Gokm0e7pX6Aa4zd2/iFu/Epjp5W16kAW6LXhdVDuCwd5Vsjk0PSU06E
vFNVHOIsE1Wy00Wqp4Im2QYkioH4Spvy0AcCnlsh6Q12PUsjlsPEu8UU1G9XQaCRums3R/C1EWxn
UY/3lhTkKBRsvwMWR8XS2R39eG855JxY/tE9Qd4aOemdJQDganxvi2fLoIsRVwnND1kmnYV8M3TF
8baVpZVbBOGzJRorCNG7JYmzird8HTgnfBjZgwPwrl1aeULKg9FL2cvGGw/CpXQfwIHt5USEQhCo
nhq1X/TpBd3Ql8w5MsrON4XYfjMFbAjpPXndqf+fqgRu9awLjHBtW65hfREDWZJbW5pi/MBNr12N
F8c/geWNLKsUPrGpCckjmVNYa8hCtHvO/p0OfyEkiYyzVoQCCcyPdA+h1EPNvS3Fx5axsUDDMQh7
kLQyeu7AKtDkZ7ZzY0E2tdbvBZYHBKoeZJUlp+lwQ67dVF4gDM67VIezuH1Y4YWirzoeZeYEwSj4
SrcMAR5rKM1q905QlISlzRtlnn56q1NwjBhY2Wtvg6AF/gY8tEe3YFLWbsVHrfoqj47H5JN3C6ot
XseAwrROTMWCUNmI1TU1fnf4OWTKPAhGLOvt4d0gXdi07q2UABD30jvpcATQOPAkzQXDVsAQdlkr
vKrF3urVN5l6Ki3U0Bc7QbveRcKcEViJwr8wQOoFbV/aC3xigfc8Y8bd8YoDPio8iR4i5GZlree3
P9I0bZp0n+SEOz0zWxex3Z+HdSNBPAgjSzFVp5gTDhD24QvpMb6qTQAcolF3c8+GTZ1uoVFi92ph
JC9ym0Pgj2AseSkwlivT0Hb4Mz2P683wiYgZC07oAYAshNSh8tRxrBFl1F5PXVwuE/wJuf5ALapc
8+pOYh+lICV7x8S00GcYcNhmgXjK5koakFtU6aLwNbViieuNGgMx8tZ4/q/XKzjMlDT3uTdXB1TI
NVYm3VwDzaWTX90+AZpdHbced1gBmFWhGsBzE51BJqmXPL7aSM6AlRPdtywhlF9/2k226OChj71V
OIHSx3JWZR5orhvja0xU9CwQmcMs37DYMns74KuxfwyOcgh3aBmxzBwwN8gP03u6Q1waXeKat4ZY
CRtM7Shnb3dBBbJmhCnYirv1SAb4l35h+yb0d0hSc14ak1etvp3v7ER4z1XbPETgqmRyK/lBFJ8k
XUZDmgdkrtW0eQiMIkdGis5yga+HTN80YqRA2EIpBuIt6OgdCqekZ78CmmLsUpeeFxA8DWknqeCy
8VJqK1x0NGhuuhZhrbTHrwYHrcWgbGz5WpBqPNElXfF/4Vzoz9YrN3V0+pgqMSwqr15d6m/YhRmU
a7GYKH8GyIZYY7CWxYJp6mGdAuTCFiN5b584Ap1eHIO0NdFVYV93U28060+27NEcyUdLEDwfC/t6
BEP4ArMNtTj0HIZjsEGfiXiwrillH4HRCjhzta04Xq5BApF/jlUQFZWrkThF2Mmwj1Rfc70YiW4O
+gT42e5A7ygqXvTW3iGftnO73SMmgM7OL8VygcUna86Ipa0EynKyVQjq9TAxyUXiCeA6DI+lpSRl
YDdsBY3ZayOa4KHpmwtRHYfI8TWGDylh+ur30tB6MYJaC2NhXbIQ3KkKNXe0Ybg7Wps1QmX4oKQQ
dG5T47X2TFUSDMZE8/XGCSzttmOzzukSxMTueEoIxvJNJ1czRMOddJlitVfXljd1GKYCo5Ns0gwI
UwiL4rjGpxyZQ9VkVehK/zjqja3jFE3XVxUV9o5gkbjmKmzhw2/4kTSaAWGKV8S94KdSlK/uMg32
zZnMVlvey4QM5cgw1aKs4Y2M3QcrSRqty1KEr/FpuYBVgt9Yn+Ej+ZMcqOvH5y0yLl+xQ5gTeJLI
RNI+GTvYkkeI6xetzYJTMbLSDchWec70piH6PITKKYa0TkMaOhC5yScJpsrzqUmgWXKTEl2wDTJr
1qxChRlUiB1AYODm6Pw0ugZk5Yu5mI13xtccMXd8+3mFHZ2QX6vTLzwZ87ZPQch8Jojx4SHCMMce
U+9nHtgWIGKiY5xDuFWr0T0vRVneawKnbS4mkO7jUKReSxukldwpWreRMbqZWbtbeOmQRnROdozg
vVnImDHNNZEodWSww6q6MTd/JFy8bDoBYGqYNYDzHcDO763TOzFV2Y4OtiwMgXiGB9gORA7QS5rK
ZIW/gUhNjXc3kfaTNzH3uT8Sc1d5HS4oJ82GbZbGVZnUuLjChvTQSjfpUvHp6/HQVCvicYoIRaNf
oEMYBJQdCroUok4A+BeDHb3yvGuAf5joWnbrsWHVbN9k9eEAgY9JEF2Gf3a+iqB8cRmyKgaYB+69
xJgBzsW/DZFtytO1WVtg7sbX947o01y+q07IlRAx5osXOc/Fwz7ACbTcRweFga4Ndh4uLSBblV4t
K3k+PwAA93cOkck+pzHBPgml3URacGeXyolYNqn2gHUqcc8jEoVzx+5xpjFTIReyNdLk2h4AJto2
FKjZYiU1kLFU4c9/LBzVnSMVcSL6eqihC3yC+ewl8aMEXQDMmEmhxI0hSeHWHS2Op0CF/CxPk2Ci
yLyhjr4ERoETioctv8gDbCHisM1mnRIKBG47lOmE+V9KM/wkBt6Fxqhmj3dl6gsicAWmnnYEAqeQ
Ob0oE1G4E/8ru8Vymqh5S883DzPLZPyKpRSlVfk4NaoemaW+L+DvccN46pbwo4G/y/6E7Ipp+cai
qtFpCdNCeUoy7qEbXJ88hgu/nHChmprbb+ZRZ+GrSCKhrj7sYlcJkKcy7Y13HPYaBLdvT4ogZ4vK
ftfOCAi8P+yKRBs5sF/IioC4+0xB19/6Et2UFaWoi9yiu4yPsFQqmGbHTUeOizWMUyBzlUt4IUoP
VMgXuPd6xOCpBk6tJOiQ+ELShQmpNsVTXrQtFmKN3YQVF7YZIRkB7O3z+KQTWVHCntntCfJtRv7t
iTxAZpl2wLIHnUkxrbKJ9HDf9gqHsYbhEbbYgDFXF68dMteyGvfdHtg+nGg25t2sN++B3g6KA4lN
gtOtFKyhvai/27WXSUZsErgI2sMcosjwHICk8tFw2tksQV3Ac3HI8FUrX/4E5BWdgWX4gr+JQTYx
KvmWBpCV12IJ3sgL0QK4c4s8Kn/F/RrUHJ9kTCa0jF4R69KYMJDKanjDK7h/6XJ5nnrgDsuOhaPl
MGqhxA5hq8BfHoBG2nyoLa1tbtVdM0ZUVhDUBznEDvZAz1qMglYYryyIL+/6XmHn4cj+iGc7pBU1
5qrzupT/7FHDwS3q11YX3j8q+DnmqXaiTdz2Ldks/zuAQ9QkYbQOHH44um8FIZmdzWuGGzTU2c4H
U9C6X2V5yKYY+UDaWgt2BDf/7cBRWts+znIdUNpMw9u3BU6/XBl1icS1mdwouvj2H2tH61LThjgM
VgaQEiyWLgeINf12TwzoZe836cp28LdBJCpVVPtFa+e82RmeJ9QMyHAWf6MCE6h5wG+3XBe7gIZ+
jsMXDWqDfeIzy1hw/NIawiom//HBTNI1brjcHDMLjYdfQrqxRuUJyofQEovlsGhjeqWQomiLptA0
7PvP0Nrt/uPmGbWe4u5Dq1VlXv0e5AFf+KooevEOq6udD+gr9jBMxYaBwHuGtNdV5XlCXLVSZh4a
MEFjkBM1AQcG7uCA2MQrBkLhZwAC/DrozMUs9CLgJcw/9KAyXQu1oIM7dXgC9mMhDCJgz647Ojoy
MwSZG25DC3z/90qhITvjub4U855b4bU0IEED8MrmF2qAYn+1NO24iLorLHaYoB/+7SjrTsgZhMyz
8m0YsJ8PKxNR2oCrM2IWVlF90oHxU2Xw48rGEzwrS61BEmS4D0+QKddUB+zqTUI3GH2jYS87d2MC
TUsPDnFaFReMzYdfuvRl0Vw9I+EMQOLkgLvhoTEPnj80GqYC1xKgzuoNSPDhgN8FSsFNUrgiAHCF
ltvSoXWhWkmIvkvTunX/713LXQdwknA6quhFkeZuskTpfhxtDYd28tPQMUU4TXjK5brWfLnGToBv
eyY8U69uEauEmTGAMucsG5w8249DKZmNKo16kTRPCmLpxHQhLV0hjPGEVruKkliNHTDm0Cp9tfVF
0PLI4cdgzkRrCcpjmoZP/cajDhiGkCa3B1npJfP0URTLOlfMFnrmQNe9DJH/UdHhRmBobBYF58ud
9FIj1Gp0EA05mwP/oNylUQayIxBzXKPbb15ZyZ2XByy5B22INWQysS6BJbnoLd1D8l5Uo3tApANs
RQByG0LObNwo6X979+jiYNFIUX9dZvkRdqPCq0RcY+k0+cCzow+s8r0oFc5Vhjttm7A2jWRoDh7m
oVoiZDr/rrYIuxgdF6DbJjipSxqvhsitW7gMxjjX/6t6k3EJushI1Z45r0LEYQbTXPjOjwwuqrl4
62GontvIUPaDhIIKJbce0TZwW7vd+hTZa54tle4AHpAiKAIitypxWcyDvK+b6wn9Rl9Uo2w1N0F0
RgK/cH83J9Z3+XPqMMZVddhNw23A1tTBMOzfBhrb7JSweOyZi+DSCb4hcQHk2RmzX6k6Q2klovcC
dghjOZTrah/OXFdiAtplE+otdpbUGTuMbP7W02cBC7pd15KEWKkG7aI9dfM6mxY4GzsalUL6BN5z
eRMbP3IMnUSwUJqcelidu7t4Y98qixU0uzaoG+WZ+GS7/n2QCBVaIyOS74wepK0UMu3CMSR1i/80
MGKOih5HXs1IypIbkTzBjP1H4eHAl8fbCvMGGTMEnhhYw3kb6ObgFaPyZJEfdt2wLA9hDTHeig0A
ithxW9we9+U3nXXMOavtCLa9HUgXhPqktDGb0ZS/TnmVCePBrxNh/IcICebCr4JWokBG2iOADy41
rZZUmI/lIpaNEyDKNmrBRsci5kmDtaNgzrPszEgb7HiDjpi7C6QmquAwIalXt22rUZE+WtcfjJgB
KZu4lAS1MiKyYPqlkLPMZA/EBmWXW/AKhO/oRIQpZq3U4d+QmrTjbpRJ7rc5m1Pw2QK9opYNIGDF
yoB7pOMSUDtg1dA7QBH4szrXTWeY95n393E1cwFwcQ8J8Fp/YsI3/qy/7l/V76jl82e/d0/AjRvJ
38+y4H7pXnXi/OyzogivXngBNhuyd5FiIsUm4jbD1+8YO1ZCO74fNMwFwSRrgMh9pGkv/CCgby3B
JVLS3S2xbmTOrlizjRKF6Muy1xXFfsK7DvM8ZqQgNi940/qAsROZACFgd/fyi1pOh1/jIXpqGSG8
vx8od0W+7IULoPhkVsZFbU6ULsBaq6Vr0vnL+iEDk2jyFMi6rZ7x8sm0B1EZB1dDxh1zkxgRY1/A
Avb3ULNL3sO9aWbnGJYbmqsl+jQ2tGwJGfz6KKz0vqtcRV8NkK4nTJLN2013H5Itrb7g63srmqWU
KIKr6tmKwCfM63i/hP1oNUtfyV/c9ZsrBCTwOW+hRLeufOs0UPE067DOqfU2foJWWHxDm3cXBRAr
S8xopHygnC3wp0ascoSeYryc8EcWM+A+oDepRFKqzp7853n4sU34Bhp5/KEVGT8I22BD+3rdCeI3
C5MT2WhtEWSnQamThLzvmG17BXnimT6hjS78FPM4Jcpvmxq/os4rLvF2CeSU8N7NTQgsWOuEJit7
gdhq65AJdlXYE7287NMwOPbpBkiXnhCnoGID83eFVuK9RCZZEPMAhl7O2d1LXNPjL0qXuNSgLAak
Cz/AdAjLtD1r2ut5c0lR4d/+lMIOnlchf9NyYZDBmv3bvfuside63VTNg9y72MAHbhwkz54hxt+L
QqA079tk+Uj4yMgszumQObSbP8NcGCmsQIoo04sK3I7lpbh4TR2ioI/hSWEF3AtHsUvp1ePEVTvN
tO8otB20tXxR5LbMEJfGbdUm25VBItIUiPzo5mUNCgH9pOSocxTbJ9ni/IFGZn5wIy7nGRbUqqGs
Am9VrT3MCVCXZY+ZOucqB3MQ/n2AxjPtTUjwLP8Hai4VgcfpTjKnkEVWqT1BYVpuGRcLPxTtgIL0
9P3NRAkT+A4KdIeJwyGRQhKwSxiFO37DusU+BjpLhzGj5HvTG0pzfEv0AbQ2kV7900Zw3W8yXgnZ
7SRanlUXEyCLRNaJnaa3F9YWHyFO2DnKPuAQJ6EcB+1ojBaUbM1P/5Z+gLVBLXk4xdL0bgNecprM
U3jkyn7Oo3kX2yDjXNiLEkAR3TDNAhOBvEqXw3k7MYAU/3EnFDEfPNkslxNz76bUfw8ieRzvg82P
ffpTfuEWCYSAAqn6WBRXh+7lYkQPnaeKunjmNBzZGBzo7d8gLWLdpOEquzRWoMjzNrtfDuVkrIf7
AO7hxRCPaoj6i396J2LtvPbX5RT6Hsn8rDHPx3dF/KuqJiUUb1d/52+sRghHGilGR/scvNHyVVLM
e5PmRnFwkEST2vTmX4p4ICKRMl20RZ04ZxvrR18lfj9UQ5zCFMScOKuK9X9PoPP6kcFet1MQvMp5
zUnU6htujPyvePphrsvL11KQ9E5KkgGhFGcZiUS+CLH529eLe7aZcZLgCm5Cg7LL+eEdiKjaTKb0
n2DjfrUw8NG0MwBC2EvtjdLCPRRyGCuCcD1yJ3YBF52ECrHPC090fNSxqqz4cXhPbG31VZBKOI8+
F19QViaXbaIbP2IGGJ/cpelOPqars4D7kcN4hmZdYr4Eur+vJ//GlKjrLGrFsUEHQOvgGhphIs19
VqsF/nplS4qQo8UIo2khecB8w6nr6255eZiAtnfjJERjJaiGVRGrWk7Bzf5H2vJdftbqmRJSz5zG
cZYyrGviogsBGe3dDKOn9W/+PrePhRZs9hb6xy2DUOID/M9Wya1+/CSVPsUASlhLvCC+Qr2HxV5c
gWaMNBFKBfkC5SHtAmradyWsXxPSoOGvejjlVMh60CrQs+pu3OD9WllEDAZ6HDeDZOwGS1cFzsnu
siTxZDJ8jxwrzuhy9asXwcknfjAC5+40ex9g0QIjWpA71EVNKDlkyDOkDW3bXEKxoqpzSQ98sF1g
rOYIaEYw9iKjT1BN1nJJAUSigzYTi1puxAWM0jZJ376CUSciH9SAOZNuAmQQoWxmC+SWSuYg11I+
s9AWvcgn/dzXxSyH8ainswscpe3kTEnv6zJoy2+1TkQovc9bB7jDCrZ5urIz5ol4Suyapybo3lJ1
P23Ic4pBAP8aKL4ac8GL4g+KOepaACDdt900C7vnzVySI4jm9EB8R4BX5uFZSzQvBFoLEfVwLZ++
As/nWEwkAScmjiSAj0bgMv/7uRi54/Kz8qrvEZj1BGU9yetIyzu5beDj9069x8l0msg7r9doLrb7
wRqv5Wdqmo4Vv5jU9VdLypoQ1U9/+Nzl45OKVM8uEgGKUgnL86ooAJYvb+QzaNXzKjbGbqQ8F4G0
FgkCLyokKeH2u5uHwY4+5Uwtunx/6NDHM+Sa3Byh6qfhZaZnkBdH8zAFjOZge0E0iXPA/D9HKqtr
xl27i0JWaUs8fRmO5XW0m000zF/t6SK4aC1LVg30TdjQEP7kZ/JDbP6YxGGfJHQE6tvwPW3otXDD
sn5BXqnER/0Txg0cXt0pVpy5529vituKlauczLuvNCDV9J2Z9TmWDkcisKrUiifmLf+Ujd/IWI7R
4fmdA+0XycJK6IRbatCIg9P354znd7RBuVZ/vScA1Y95kYt5m5mgAI+0UV0BngcAyoFVQTDVHTCc
Yt5nkj9YdHwTU8aCpnzBwFnh95Mzo6xF1ixHtCIhep/tuAhX4gZPNs6squGWNX6M51zQeDe8HnoE
cokN8/PrTSUWWjmCi+XUc3CY8Xt0G5KGACy9NkJRxtfkCq4hkqrVc3QNDoScgEkqiUIJe0kClXva
6rji2DUuoi4p57WyH96HpW5qasA+STirROXNKLoaOXA1HKmBVTMSkUVr04xJLVp9QBfFNZEBwje1
nYXpnHQ3GRJIclLRqtGJAEn8HDP1m7AGSuadXUgQWKOVpvwJK1ZMH/NqZstphg4ylTumdPNjzv+7
VHmRgFNsJWX/jz4P8c5YGOI+8jH04CXIY+3LX8OUBE9brvYCI+eH6dlk6OkF1pGiuQ6IqFI0AkmL
Vf44kHepc9HVRxNlFSt3TOMjaQCIvpTXd3FDUFNH8PvRDzP4L0DHUHenCZrBCRaW3EFHWiUNsPNG
7Kj2BcoM6ndE9IviZ9wmQ22od/7amn4yJGkYq7mbYpH33CMCIG7fXdlv/8UuJmeLTj38w4Uczq5z
09W9uVgOxQst0GSoLQK7xt7+MRLhB3aE6hCeA4xY2OeBHOqGWyanAiMS7Gw+AY41OrFiuZQ0WtWH
f1SRyXJPWlsOwo11T2hBPiLEjA8hm/hah5a6e0LtlJ2qL3XjmK1vUVKofz8YDS4Hj8shvQH99XxV
2EU+ykPACtF4+v0klJDlDp8oBIkB3ftlYiSr5a4lIGYkE8LdqqEzqkY4KeXKuewIWH+HSjGJFR2k
4mA4DkJpJ3Mcc0fbhEOdOHrfP7X0UEzOno4DydoX34B0TKS9xc9Z/jiWbcL1phNeDtchj4ibw/tZ
C6D55g19s6jv4AJEOaUsSCnblpLBJH/0fpQeSmnjIqb96KVvEo2aX+y3AlJ8BB5V5LefszgpMwx6
hLFu3o1aeZOk9b2K4P4xYGip6IEVJIy004LM6mrIXu2kkPy6UZHRw9bXdWbNu69PyeBFh87WU3Dz
HgP1fs1Sydmh8fKzgnjK2lDvrgIeM05z87hBhYr22ATV52ua8yG2seG4gkAvKCtQnfdsn0uaLEzg
nEp1mfFtRqIZ9zJ8yMvfonObs6d7FMDfAubMWgXGm4OnfgDiOQYCExbdmiKBCTN3LdnCRP5QFHrV
+odbKNvIWA38fp8jFC0/oswaIrBwLhT3Twd9fDtMQq82pOvDYJnYcgTTGLRRAwCQBzHYapF9aPqx
ZHx4pAs6xDKnEBw/+tEyo+CWLdgcsYlu5iV2zmqSAvPcVJ48Ij9q2nRAl6cSxP4JUtdQFWaK6zOt
PhScrAc7iMcX28tv0pr88X0ZxmISyZ+rqCpeaKP4+c194M3NejhW8DkBbxpx6EUze6VWpr5dM3c1
qjl6E93DqABPdOXIYi27NViWUgLqAYcOpmcrIPLKmeq/cxn+iBjT6rX+iVOmL0i8QFUorRGrLssZ
o7YkTxmuyWv2Y35AZUPOXNvRSu4KdOCUXRmMuicU79yY7fzm5e/xSVQjt5NDGZQ8b7mGDbwsDdc4
aWKL95nQyXbCOEy1oefLYfo02pYd0QZYhN8dDpHEHeSOXLSLxDT5shHOq1mI0PYzoai1Xx0uBZRV
jfcBWW45Q8sh/CWIrabtDZbfOiPyJDBUkqbJSV35rRIgpVHvMggW0gwkQ1TThE1qlR9g5me5N4LW
NdDiQuhAMqpzPU6OBsUHTddZQABPLDZ0nI8iYc4BS3ht0eGlOD01XJ/74SlXItUnrTbUi/j1F21U
dvaVL/GRtqPrbsQvi7MSyJl+ceP41LkuP8QqryTKJXUcVUC6aOeuMymFCZicK15MHNT23Q91iMWa
JOY2tdEkkAZGH3LNGvCIPuyMKV2hysncMjOmvybVb8Rizk9cq7Tlqb5983SldLR5uW3dRDOLhpSP
fcn58WxKHkV+MHrvr7lrBl7UAb+KY3oCt1QAG7xoUgdg/XpitDk/srpPa2IM5zEMvxv9uUcSBtRc
t+a0YwUSXP8WdY2B8W/7Vq+6Gc7fFt5Lhngdgk71FqTibtNZP95KQUyS4cSZXR0de9J80A3Mz0y/
hvmy42tHMkgOmA7Ox1xj1G/3EZDrjdP6DaJG7OeKmAEo86Lac5jFT3qfc556q5zFwgRJsrvjGr7E
SViEF9Hb8lllPPgcIPZ9o5FciJHEhNj/rJwnCay/oqAIP3P2LvgvdgM8PmEcQ0+2EQyPE74yDHRr
1LcYd5GDiwNmBqBOHpM5WSSJtPplGgoY937e1oqFx+nToYaQs5neWnyv4jZSisASBrtrMLEFqnuV
4pZpLzSywRd8RkorSx9A+hAyzrwKxYIwHI4vmJJuNyCbp1RYUav8C/7z7fduCKa2JmZfjzCwGDdM
7aTcF4nMkn79V5tb22EualigjaJEZT5LSEDyiNGYIfiJsFMPt9rPrk1B41fIVQ5AZMF/Cl2p85B7
VmSZZ/KI72ESIXiw5dhFQ+/pRFa/nBHSTdKqLSqPJL+BUm56y5rZD0CayhZzfrO7/d8lNmOgj8b0
O0BqSvIla3gfhKky+7LGy4I3PzH3ydDFuReoBOIOVr6WN5YnRHkBzJLYr00izWz9rcERK+qyVHw8
yXx+ao+UX4aw7bn4eFFjOKFQdSFCMIPvk+0p7AnriwSG69La/06ba9Ndj8tt9yywk9C0gKDNIcW1
J8WHmc1OBs2VsYJHp7d79geZYUG5xf2v8fYRZPKz3WQwEnrQI0/kJyF/RJ+fe4VtH36Zp+C+9kto
P+Dp9q2THieQf28aDphKshJH0ldhGz60NK/0MS8C5HpQXFkI4N//yE6pk34sgQO+SoPUgtZ2H5PR
+6dg06oANAeOSsnYOLthJbAIauwDRwnh9aIoanxflUxRnAMW2M4lInDI15hTqRlI4U6gm3O++DBU
C6zoGYN/Cl9UlPODOKy+H2IXCs9ToQSvcQgn3n1er2tzhW2KhmkKbMmJtaQmn/ZNOEIa8V3ZqtRj
xhiFsjZ64rL0aM6SzJuH+wY4BkU2Z8d0ocVS+peWHgnSOHTe4ghSHdP/7rRea0T/70hC9pJBgC0k
Dje2P82QkBI/O9xEjchAUIISpfalJJ9mbOOkNFas3VwdImWCCAFyidRVATQKdOuOVd8hy6sBMI7w
t8EjJT0YUhlxjyA48wc3FDxkze7riVXjqB7a5UW4LKIbqKEPyxUAg6LZhC8BmzBBThuSmYBNszdJ
tSMPTDNPIfMMe6Q5uckEoYsLu7tR4Hp0f1YYNSwZxzZYsD1RAc5Gj2UxeMaoA8+fJ/1LA0mQ4pOy
WyZ5uUlhZWekhW+2z/OEq/PbNK+Nbvlsve0XWZQ9aT8Znxk0j1xhQ0vSyl9EuGXQVkmuVHHZ8Fyh
e7AtvBXKoXq+yKuiPR1Swz3AsWfNCARlzH3nyRQuuvyWIqVlTooitEYIq45XvyDbBVVcsjGjSDI8
MHEUsD3c3EheaGfqsXiDeJx4NcJNqLhEErVx7mg7xgGNPh1LROYznn8jx92WfghK/8XHTGWHZKBP
a+ZWUy26Av+UhiHtuntZeSTgfKfde4HE7duBktgHD86jl0jhJBnD6tCsun7JRBrJ0Qoj4fd1b9rP
Y3bxrW/mZRtpUFjp3FX5odZzlZHIvrjD17G09tfnTyNuq6dLg2yikQYb5EiR/sdr47FWGYlLgir9
mWhIZwEkEveaeTQzydQfapxEehxce/HJ8yCFsb6igmezdb+vhNr9CmR7EeA88ti4vMtieHQcp9CT
16uRdmm47lG4uaEWP84895j4EtC838XUQhpOyLv9oUoQws54NF9aDQx61jrv4jmkutcsakd9GBi/
1scYvd9nd6CG2eVT5kza9/Wxs/fAYjZsaMIr+nMQtRQBHW0zQtiJUSBL4YE5BcHosXRAZtYqs9IQ
x9VNS3NyEkrLsO1FlQWlWNtnEmnOEVLSOGCYl8J4laY/UMTnpGK6yFvP73OoeFBFjWx3wQN47eOJ
sWRfwT6gtVYtOnvGv12Sp8VN07bYXBI/67VThkj4tFETYH/lKd3DghMgw7IbEzI3B+SQ7Z1+41WB
V+7j6xFn4h3J0TcL4R2WbvTwF78XpBkdJn5gVPPVc6aZRpIWDZXoID1H0u+/z8D6AJIZzHyiEJt2
e8ytSREYBnao7PX4c9rZcj10+4et7WT0XSK91rUJZrY2JvMDcigX4tSeQcpC49jPOFZD9fx1wJz/
vVq5GWVDAFoMWfsWlux/uGSWNxBcbvEjWI9cEgmRmIw6UUw2OePnaTgxQhsQqRLAiUqKNea4Or5s
z1vO6ytTsWfAiODAvALh+be91tp+urdGeEhhYHzZEwMM1IN12Q3mOBzRlO3vuzT0SQ8l1CpNWymW
U4irW77Pb51zBWM++ZJYzU2miM6xE+51xDSGM77M60b7f4ThsITi3kRnZ+OTt9eG5gBhmAXn0nR7
BYw1Kndg+wrFnPkIvxO1akbTrrilehV8Oi7RJ83M3oqKNMRKU37D+IoNCrSdVRrFqNVSSN4Jd3eC
dU32hlkmPYPBTJSHf+cMasJ/XqBYGcwtC3sRnxxdTWSUfpeDRIjsr46FmqXpQKIjAsg5ufLd5Uvj
ucZjonZjt2060fPhqDgSUPc2b7zECPn7PHOdmpUrYKGDx8T9nQLGeqKBeUZ2rVEgDHmztd3GpGRb
kzY+bBVmOXHx2ZmKkjZpoqpqyVMYujZCRuZdIe2x7of2uKEAYUciyBWnnsANGaagn6XVomKsOJM9
HbmnSl+BFqD+nq1k/Ss4HZ1oeSKJrZI+UNFK17BBY4IhXtKobmUhML0QbH/VkHsZ5/BzDwyzr2Oc
0jTf8jfSmnOVbXNoVhP+hYaOWSYIV+tqiItjnR8Dr+0FCQNxDanof66R9PNyTYxODK+zXrUClv5o
qRM/Jif5unzXQRQnXswQ/B3Ms3QP7uaQ9d6LoDei7AWMBqloPNOSQunNI7rxXDDXmgHYDaeq2CI2
+zVL4R9nbSL9Gp8Emxxf34P0Zweg5U3UWJb7iBCKxglAz4gd/UGR42O7U1vh2FgCEdE673RM4IU/
TL77UFXQQmI4WGNs5JEWoqg/VOpIPSDCXJ/z39o71Kyb1HQll1EYRuv/rOGpRz2UfqaZ0DQCclZo
likp43ljx1WIaQ7CRkutrziWoY18fAkE9uAERjiN3rJb+l4kFQuWmdOeqk9WraDY5St0U1JbjoWc
oGjivCMw5uHb+l4/lWL/isbA5s19Fhk/vOzjCS0gWwmyyRUM7kGHFBVyYg2IpixCz1IQ49EI2aI5
MsHjdYVu4uzfndbFLNhDNb1MbVzKA0pNsES6Msc/2mkSZ6kBObwE/Z4vwYK1LyQBySlZ09zyVF9Y
wMIwUWhByxVXhmoZnlg77FFaCqs55e5L8jZVnb9if6Hp8N9YHwUSlXQvDTLCwqLBIOMPMBCwUN8t
BCCeH1ImhiYZd0b9Qu76dKF43AoQ6JlSKUiDScRpcPh1dZfAUC/rrRCtWVvwrmPzoX1zk59sP0BL
wVBLYS0gGUO0LEMPp9EpUzJvBdHnVk11njqMtIohZr3jdR1x3jhk4rxUHS91KNRDzaBb7L+Hqops
5hpW2r8SfyJfKpmlb+0MfXyePwhbLjtzAy0EJCplIuUM/9xfvfg7nsfct8eK4TtK/PaIxDyBQREF
jmdrYiVkp226nsSDM4t4+5VqwauXUS78DTP8toNNrjqiTEtFF6/hIJcpY5vVna1yvCbLIri63/hc
BL8O5uFWtPHVg4e8vFlrDmPapgUBHoIa+BgLWf7w+KNVMwgqNvSj00Td7Xaaq3yObCQIBIvmNrfs
WjwKURBZpWjhV6mvNEbogt82tWbRPV//PO7nBriRvON0+3TrwdXJNUAW/rj6qM47tB+JWg1D2sJ5
SgUY1xdyuSBwixm0iaU+UyKX3yHnz0cFUuRXf8JAJHbmbIWXVTm87V5K45I3m+d1GdAkH/tk8eNm
eJVx64pZYSxyim+Zihy4pxurF7jAZeSqBC5GWP7Kxhx816Dw9xEGbB5xZA7XiHbDikYW7gcoaNk1
VV/2DqmtsqI18VYikgf0iIV7yQoQamx0IprN97O/xDP88nJ7U2aC5f8Kkax7Ri15taFisagra1Vi
rJBtujM22fioCvpe237g4KqhQ8Mhbh+4o4PXEg3yUm0vK165mAnsOUpv2A4wfhZ0GGXrIkzDnVs8
5vHnh0U1a0UL06O7mzfK0Tqhtf5TDlltd2IxS+i2w9qDUJaGuILprzKUlSFr7N+XBWZntCeiwFR6
rJhR8zZMZzyu7MC4LITyhoxWUB5RA55Nf0h5LHtewfIxLsvUqfD4du9XkR1apdEDkm9pW+BobXWR
NY6WXZe54F0fq5Y2CWlJuiOxIHCxtb99UI5K66NFc8ZDV1LqrjNXxaHFli/u9NANmg48EE4NTl0V
YczyDjsOkSsM/K0AJHkmmZHHYVakDm+wY4bSvXYhBbCMydpGmJ/UVB1qpbJRdN3zqMmQ4Oxa3VCA
zUDrHR8MdybOAWN0GqLBa2U1KV6nLvHk5BVVDjE6eg7s/BpipJJpEDKFyKoTfd0Hv3ACpWkH10WS
EQPW8kqb2Fs/+fJr+rTnwL5+q/C4elNihpzSemZmNis3hviLI1UFDOiuV2V3EeQMDy6ZgBGKv5uO
oZcwzID7pYkZRVEOkOyHqCVfUUw7t7SWUgXSHSYtV8gv1uijlTx7h+U4FWGoQRqf20s3GjM/yAAl
ahmQhFjMigvt0JuLnzyxRlJ6Yod7580hLypSvXC/LitmSvXvcFGHxXM45hQmZRpaITj8DXEA4TmW
vXQxjx36s76P5ODvkRVartmLgU4/RiJr1kPV5/0Wdr4sBHSZ/CcgVV8wtwMH07OtLhDAF9W6oyEX
dcUDa8NIJLf6leOTssBn2lcM+34IcLMfriPUcBDScs113Ya+RomnSqfNNx9oPD/YIfT06iIaaKUz
+N5GS0bz/7uxpciTRUAAz1UDpEiYTuh4Lb6EVBb2OqYwKnaXfKRlOe3gsRTkyS8lVnWJOq0+n508
RTxCZgjc3dLjpAZ6hCpq2mhvMUIq8ustldg1//UjZp9rilFxQcE0TY1ZWzu+ySy8FO48K5jZPyLs
js1l77YxGgbq1RsrAO/dvNwwhQq2yeeZ2x476ft7M/feCDsuiSpfwIE/TWOLjw7+zECqV0mU1gbf
fde4I6IWaqA2W1YNy/nIC0+YKSO7GM9jZig7iCKG36w0LdjPJEQURvcE2BWi9v7Ek8CUxvcd8+7X
dvCFc18ostdDTLa8x1vXE5Foaua+rGDGuMW5FGsPxFbFpkz00UD3KXwHtETyv6Rlzx30/heRnVAG
Alvv5tUmpos/Yown7dlEAM6v38J032pBt9rQp2OrflZZIhp0LCNEHvTpgxE1lD6mvYGk3kzIFqEn
BI/E0Ukq38jvFE6FDsen+78B9l5Izoo84FCKQQryIufKXjP+I5wUn+fnQRGBZJvzjoajODSMt0sa
Ut4P5VRH3G6hazQ+GuBzj0qGCC0WBBfvbxio7aWp+b0ZAHUi64/bkbFTNhYdFZbEHAIVF41W52+Y
StUGABOSidB4V0ig5yZobf6AreoqwBTWpSJ48jbOJvjjJ2wZFLCMcBO7XQP3Oa7mR2dZMdP9zS02
tN+b77O3Wwhhj53enX2Tj64SJ5P0iEzI6UjwmkEvgrD0/+YMcKTKJTo8GGmJDcaQYVd38iysqcLz
/rF/jL0qnJVYrfwfqA/vHeIzpVF+5HIxN+M7SsYi3Ma7Oy4yZ/5/t0uOseR7SYKr1CpLVEwFh3jm
YebFs+AbGdY+FBSRycBChb62PN+lSr/fFa5tebYOzQeHd2aUvNWfJTsGIlkroFP6HzblbITMYXCq
+F/3Nh1mkdKDNd2n4Y2l5hXuGQvIhrRw8RCjame0OhoQoIaT58v2C/yZkP32zB6t//YRxQ9wSYAx
As8cERK2XrJiEGy7E+bSphfMJtpL7Wtm+/2NArsUucOGP7WPL0IL6jqF6kUOkiuQK1FCpqaCTrKN
rbynlQUG2eVqOxXTr87CifzMWQrtEq+jcUoh5OQwAJGXsksuUmaLQ88r9/RtcbDFvGq2mpYFE3bO
jQEzG+oeJLH+jZvqeNfVnG97daf6gq1GXyXhYD/+mAeTemycVRBSMQiobUR14wJWhGyUsMApdzCZ
607LxPoSQe55kMkVxyDDD7DfCmu4XDg1f6i0Uo2Gsa7LfXMtFLjomyxi7DVRnHKB7MwMbYC8epLr
ylUdSY4Lj4kzMCLiSSRybPby1EdWfzJYQvTqnhSMwKAZNMviHUu6sDs6rrnPsNccU3085gc2CMMk
fff0ow1IzuZuE/SsZHH6bwwg3FVZg0JQXjWf51zRB2zbUWZly9OL9caYuaJYWE7hiBTMYhdUQ6bm
lwbTI03t9ewKi9BKheqpRJf3dPdjD+Si9kcbtsZ5GiQEezV+F3gXuXWUrxL9ehP0unFei5p5/fm2
qSPdjv+Bv5qNRvZ0cR+I0GMUW9xZCY54jfUp8g6skYM1NImS40uPQkT5Mws76a6zi56OjnKl/1OZ
g++WbBEr0Ip4W6legkgc41tTSkRjwnvG2TqpaeZx55EuYQPxT1YP0mVilDkWu4driKFEIRJVoetB
x487woKo6aqRfxnCMb61qdK5Dlb6r21FcjlEqCvyUapFbWcYlVeJzxmnDd82gDhiNNbsETOzrxvf
3t/YSA6K2erOb5YsZSnYFGUzx2xZVxujKbz4EzMBuVxp3pd0Qx0nDVzs7q9HdQFGKKS9PgoXzzQB
bX40rJaAx6hQTSRdcdJAVu1C3SiMRnAa7bQ7cP1So78z8IOPxQ4MSL3aQzSkybwJpIfbrpGzBy5C
bOb30z+xhUabicQmY8UimVcNlCR2FRqfx8vQxEullnN2tS/81yEx1GUZpEyj908c7DwZ17peCXrU
LE7FrBNa/Wdsjdj/Aej4Xv6/Eke5izR78xGC/IQNtHCzjfWHLiiJfK8cSOQMFyZhof1D2L4Bho2J
oWi8LvjHSFpO+wJsCIDCQP/3HEUgAiyCPUNFykuqPlKDf9PQ+OWiT6HVAnW3DdgFDTS4fqBnGrmA
eCCsLvyG+ym2OFtISKek9pNs4NYVDAiCCW7a/w2mZRnoWKd8r18OejQEcHrp74kJ5omGnKCpoYhv
lrdsTGAXhXO0SNA4zOvMOZQ1Kqhht4RISm1Ou9wcHTFStKVnjRPYikisAi9sMV+9+xjBIEvqzAT0
8jfQZIeRAXCobFDDwOJ/DmF1t69jaiYJgW+NgfuXuwo55Ny7n1Atf4FfiZHfd4fLmDDQ9Rx5u15L
h77PsJTpvPfjDI+2z2CJYYU2btEwfxdNHj1bC5+qujd6J7VNfZTrSQRziLW+H5Bn8aJ57Owx+AGN
UsTKr+LG6RY5b2k4vtW7W/sOEIamw18Pps8XLhOxahZRmWTXWaLOI0Ix+xQeGPRBbqNZyancXabd
H55rKYymcsGSW63f+2vtMbVRe5fmNNBdQg8jDIzOtcr7gaNUxXMDfkGMujaGqJJNLggUCI3euhhU
7XJqq03CFBCCm6GQOqqKaC41PsDmmZgzG8OuUD0RxTUgppUWTq3mYF01E4xXOqLDJj6qPmyWAypj
WcFFxlgj1wDUcrqUGYyrh1i1IjY3Wo/us0e38vaqy6HUtELYvVwMcll6tkT92Zw9aSW/3DeHmijL
v07LjHABmsrPcyddl5Atnw1DidMGMA5bCKAVwthGQ/y96Ymb0SiDsUsLtZU4hDeZ2EXCGal3KCMa
vQJdTNU1+2dHQmlHLF8TKzgvgcjwCrm2K8wpC7dif0xD1ov2ZzvCzjKHBFRc89wTkl20bv0VucT9
FnzqHJ7itvtw0s/3XAreYCZ6/mnxy9pwbd4CnroyFjeGi52wo3AjPzMFd6yitvjSQTZm4fBaP5Fl
ywcydxqryHyQRL/oQREWz0PLpNI3P3NSoqRnKde5GPnvo922PqoE5+U3F1OemfjDX5HcAbsPY9Fl
XOnMIK5FyIxxoS4L7FAPN9/yjoJ038pgSBlAvz27LRxe62Z6TzBwdfDISlCokz43WvRzjkGexs8l
hWRX5BHvzc800V3l0ZTwRvFPSyYTS2UyDXOUX+wDTYidNcNX97FKV0phmvoDDw5G1y/6QG7cgSM9
Y16AuxRczNHPzyjUNwywPtdbuGSiWTPG7cXGI33EtPmscM8x06y+f2p3wGAVMM41Xp8pwsq7PzH0
DXbjjmVSCMAUxcYNLmnqV+km5vFkiewhPcl6P3/wCDkI1uI6UV4eKi30x4pEVmfLpjpYshrLvBKy
Vd6tIqo9U9ksywsZmRRLIXx9Pzds4lbXhFfEPW6P7NUEVUZc1I45lRtMfmwfwKhSpWx9P4OrK35i
eVMR3O3nFuwSXe695iEKStWfwR4nE/s8la4VYPzu7UvaXT+ByRxdaVnR3lGxlAf3t9q+g+1M3fuL
1AG8n3Sfnf04h8gtAewjk3EL8pQWpZgcB8UDwPrK/9mq46eprTo+Enn457mNJfMW8TRO6anwgnyo
OXGuQ0p8ILLRDnXSRYlW3tzRL4Q3+1TlSo/Q/s2knSbiqQcj9cNjronzIr0UCxBsn7tIt+HHdn25
JaeNxXlN4FNZ+K8PiJa6ewD+08W9s+EtUdQLWP+ZD3D3zC7IcYQTAuY5pVAap0BCDpdKkUG6IHOH
zooKcoeOIpHneYjdTFVD9sO6HDg4ouq93SSjbXyYPC5enO71JfYlGg8UeZHtax+NMf3FcBJZ0e3s
sSj2tv9lCa8HD6WPElzhjPcFvUbV60lo8PPTlC3lKo63TnNSAYWT2+dqb8lIbeRhD/1rF7XeInC1
BrGakbBIji/vZ/7PJfrQPerBSfa3JSNx83RVBzmJQsnGd8GbElrWacH+utS4SHL7KwrZgBBzxkhx
7Gy18DYwglnEup0pvp7aOfVfieHE5vm5ZXrG5zRoc+JGoO+xXKkuez9nLEdFDPXjz6iaqyldGHrx
L22C/7uV3cimMTC9UdxZN7fLy/ROJguxxR8qYSCZHQCF+6Mm98FykHwxfosAW4P1g/u0qTeDJGOT
tiV9Vht1WD/C1XLV5ehqO16GgnBChZMxmGTubRn+fcYiLvzdo4Ull7D6Kc+N81ZcRTQfYEd0+TdN
AjyVpc0o2g4EZmfycW9BQRt+VpK94vqMvIxwOouopPdW7qNKzJh9RlnK5zxk3BjjB43Ltvnd6Wi9
1bkiZvpuRErBmGgWVnzCv0WTu+aZ4rglns0ReQc7w+97P6dD02bZ2k7urGOmmf/Mhw9idXv+VNdu
8FBQ5jn18ve9ExqJTXPunjYuK7j9icvrE2on5uk7YlyP8TIGXejRKaaFWlCXbZNVigqdNzMe4VOV
Fk2eZbJLyf9Sy5ALE+UOQH9SWm7dctMcecXmyYB3tdhnNjp/t02vxYb7Pzm0W5DjxWpd066fUL03
jSDQ0AicSRZ79ziv33dlsd/qgIFL0FPaCr3igCiRBlOp5dgPVfbFYluRqwlg2skqTD3WVnXk0hS9
ETHkdumrvpAUom80gR42JCj2ETAxlO0M0G1IO3WvodWEWQ3Drg8YaBij7mHJW1dc28F1whsgYeSv
mho+lBxmBJHVanoKDTjQKitH1Pr+CkQGl+e1e0koOKNjAEHCVFnt8LzIKnUZLovBkzaOEWDRprfx
rjjHsTqvghl/7cjsZjpplrvyaWPpp7ha4KBpYreolPu09LatAP+tQ4R+Ep5m0n6EFKNtUoU8SUTb
uAmERN+xR/c1NCnTMKPblBkNuJ2BDkXSeLmUFs5aDmYuZsAficuKVCCmrFHgUsjA5OhGdXVV/bd+
2FA+0OySPekqrx3rKE9H2jvT/zhaHIexPAXuzdTsxl0siC4aLhxsADsmXY+jLPq7HAjdnWfzahr8
dPqfM3hGy7qd0uA8cAzBvSltNghNoApsKyLUMfGVnG8vWGsYfaq+jY70zJhNuDIrA7ZY/53g62jf
1HnFnTvnit10IK1O8k4G+C+9yAg/z3Dtl8HZwcUXIaZKy0HkyMXtxpUZM/TJ/03MK1cH4gHyxsA6
T8lLBvUa3UWA41RREbMcoM+R1Cgtanvj0KcAPpg8Wim9IUiW1NdDGVHrtanMacnM/FWeg9eeCKo0
nJwXaqY+sGXwCFlukFbTN+riXBuEbYq4vEjbNM3nr9FnvKIoqOimrCntGdqkWzEzvCiHJlEvZxVe
47n/2UKG1wxI1q1Sfm021DXmXOTKf83Rm+kWnqyKlBnY+BQC+rElxVqyV25FVQXd/akWNommBaLx
PCLSCtOl/7iQEDUPV98ZnboOauOrz7rNrdx8a03UxsBflypbpP6aMR6eP8kjN+Wc6pZ/zx5KZ0QD
zJglWbNXzxjAPJHlCaFMvudJ26z3wh4IcpyD5vwAXmGBiTlbOax3LqjbO6lPekE+PkHbG94AaqBy
4WdTcZz5Msm9MWR75UmNrLzEAvh7UYRwuwCsDecmZx0ALtYg9EuMRDDK9BXdiMxkOtiWeTGRhZUI
vXAZjnvHMQhTMHdNZXrzGDbZ5jTLMZAD1PYWzt4WqBESduIMwuBJ9DY3TncyMfX9WuCTvIwMYcS5
xfg3ctGSTGYbmcaGcOqftnwKizELb4hzc03Fum+Ispw0oss9l2tUFKpxf9eggX9phCQ05vTBVWsu
Ts7Jogn827jUVGccnjCpD0Gp6WagQ2LMMH9HyA2CV3Cdov3clc7DHnLr7/bo3Y7ETb1h//7xzmC9
aEWZ8GOIvtTNWV/rz9yMkSCg76EDahKHXRpQAqCtdGNNHRQd7jRJfODC7vi+vqPnljCqo1LYEQMo
Drt69gnti+TtjeBrDWewTXJsNexITo22ZJuOE08yj2z2CgvE+WqfFHOFQRm8HSXuifz7UFj1FazS
e8HwFB7lsfQpZYfglH5SgCqrs2H/Vkm5/waSgqnFUzT5ZRtjV/rGw3lm1yhLr0xUGu+nTlTj2lQK
16BE/5YVG9QrpWcAtTpuyNn1DN9DabDHwRmHwyduWsHhYteNeXLgavISmY3WbOVk8igQFZ2nBusc
M4RXKngce0bogslvfvLlGHJ6JXHAfZn1j7PoGUaCdK4H0fWNjclzO36n3ePLSxal+nlb44oFC/gc
bcZSI53+jE7xIBPVQqIoJoTCD3PTyXXx2nfGN7qLq2XgyCfJFYLKoGu/sYxRRhD/QrsX4yMOwQ2Q
aUZB6emsaiZfFkU4kZnILtpsK0VWRaj8SF8ezeYFD431lLiffaaSKEHw7VjGx+ls7I8rWDIJfWyj
a5PaJtK1al8ma/serfY6kVEog13tp4JAfnn2UBRVVIWubzbPB1TXnR1IsSjyl/M5NRjffRONvxsH
TLlyPt5fgKK030lCvcH7ILKtBqfkMjkTCUuUhg4zAOuGTndkjGjG4vjSiS+mTnhNq0GgMpRb3sLR
n8IqJomLRnCOaQHmKq8aazErC7arrzYcZLvUiD2CsfPb+DDChJGh8t9VXn6pHWsxeV71BiS4ms8A
sO7hJ93IzlztX4IyOwr62fCsHF90h/DmD6Vz5N4BPuIuHim4TvSitUFJBupda5p72Y0jTXd8SaBc
ZY4v26oKGR+K/ZWRO/BWLyeDu3eUtBjmnf7oBWGUZCMiUh83smF1Zv9+4CWctEtpBtYPbPFgtiyw
QVZvNsvSuZQxI5IPed866w/cJY/nsSCgVCHP2+XYL0o9bttPekkWJwD5DoyaV/dYycI2tX33hJyN
8qa+t55/t1r4Q1/qzn67DZySH5vdlxbW2W/eETDQN/RJjXcyTl7FEICSqqckEloqL9GS3UCLJ10p
SxVT7lqDSbcF+JERC36djy2lG11nELIyIA+15MG4KQrnfQqdBNi6vgcS48N6yl19CuuXftIFRN0S
jCeWCPoZ+43bI7TzV3LcsS2DiHXDm8nLBkEEMYo3XgFzMl0p42tj8g0qGPJlqApFYoapqKF1mmpf
O2fJRPKp5WHnj9dVL7E33OrO+W0ac4zpaccuf+aYwQv9iyGXdYeZXwWyZk9v2sYaLEBjDpYq7oHd
7mBAQ1uYtTAvclGHOyAv4fPSfMEKAq0q84rFYbM46KDlesXv7XpNSZ7zO2t2rXZKw9mSPoY+h2oG
WfUsTg8DFZdw+3ajPVefHoap7ZPZXvBODct6/OOjk/osWtOx6u5LrZCt8K7a8sY9/A0eCUtipNnY
cmfbVO0FjgPrUJGhPS8KtZuackcCACBgSuDIET4iglJt7K1yvVUIZSg0eI4A/WuPbFe+QMn+XKEN
Ep73cWVnEGicMuPwBsUHuKqo5OnnNK2lnkVXADCD3fd7g0/oSzvu0W0d0Jps0Zv7vBU9GHRSyxbv
5p+yXMKm2qneSwWQUzL9QCEyfCUgmwlMhUPufaK3ei4PIrgD9TWZNIuV9xFvh1kSZa+e1takPWCC
eGftLwM9G/he9DgNq1oAIArTq0gZohgnOLGsM4E5wtEdkyJjaZ55l//ThlG7yOxJXSxmUcnVj0Jr
vZw0sFA5kSWuJrv7FcJqrMzWvjfXYG8OMsXu3pRJODh3FMH9/kFVVnOQUNbBPYHF8E4301psnt75
3qiuSp082FIIfyNg8G5hp9GD2jhOOBgz5ZIHz+D3/BLtSJHorMe3k6o9V3EGECFjrL/+nWGHly4X
N+m3JyBG/RESr9tfT+x/EN/bAlktiYobh2EhSVYUS15o+4Mp3hO1TOeJBR48rdm9kANFfc0PrZXg
EBORZu9O0eykZL0jzZuQTxqHeAu7NNJrKn2u53ilqhYTWc0Ty3xT9P8M2/P4U+l18E4F08deoO1c
B3wNqK1Y9BHJfpvSONwEQsGhSFCG03+op6luPQoO1YySHDlAYpKKNea8Ns0TTBh4Xe3q9j8YXjdI
Orwrs5p4rM5b1M5aIh8I12YgyX69aPoSNDLc4d/bGfvegqF6pdFkb/fAF9ZbQKAp+BIJbmjr0QKY
KB0be4CrEt/UBsFlaefwdJqHKIDcfNZHzqW7v/6NZ5fhlB0bTABSjWRGnYWhnQk+I+PkOoqLjI2I
P0RlQ8AHCbH6xwN+8cL/GWEn3LU+qmiWpIQa4r+Daud70ZOZfxHtunAegM1LD/Bb1w3m0JKpHEnz
gvxjA6PwauZH9oySkoLWfiTs+9hjmHVSPYgFapJ9L05bbMx4Ef9V6NX3uVSTdD6PbAY9sAnofD2U
dpm4Ut9AsXCLwiVE6s/RIGR71P11fSrJBVhUtiHj+3tj1Ip/Z6igDPeLe4BYxkybDIm37Ok9Zxir
FJDYiizjPGuOPsAZQKUiZiJ4JT9cli3UYDeMtTjh3dnRIhLJJ6fLzAA+ncLHXDnfDxsV/jGTgXd7
zZchslXRo840bIzHOzR2NOZMalTLgW3pjg3sgk6VpLi+sr8wUMOkfj23x9WV5i8DcpzwlL1QUU9E
EjBQsV7fY1w8ZxyOLX3G203KUPI8A32Q7n+QtxmovdhA5rZnQymcXrH1VgOMniFw6EXZbNSF40O7
tQ+Hit98Bg4TfrVvzSWGhOsN7RvZrDbBXhQOGKhs42g0iIPS+p+SDBRcgFWSAhn3B9B6y5OBkxV9
y1VmnSY7skJ563FJxbEJRw8FrsD/xRKFxGcsV5DZvir0801+DD71MLVUMWkuZMcqOpBZyymiRv8/
ncLGHwLwK1lLKYOZCfz+g2cuCo5OJqrK0+drbtSKOcOc9VilbEgGDIOzZ5ip7NhnKRMwCV1j+lTH
cW6Z8s9r0i4Na5szWX+qM3hbPTbPgVaganDjOXWM+IVMH+FxTuencZt6A+1/df6IadKvN1hqfGKc
6i+J5SGfI0SrBhmBIFIpGIhKG8CGpCZnzGupWnwEdYlIcOvLQF9y1+8EnwrJKxENEaCpmElcD048
PlDTm0XuTYrhzUzxZa+bmiZfZcyNlgl35zy/Cl/mCe8LGMfJSnQBIAabPHDFst+AQPRbUWlxoFq3
K2OyyONhC/bwxDcyuwyC0adOeF+wdOoE2L02FUbXAiu/GEmQDxRGQRHmXaR2B3foacDXljXBqDkE
Q2uFLmtPQpHnB+ghmelg8rh57QwKARfBujMMDGyXEzLRl1tBmsH5XLxesQzKg35lnXkmO8iCOY4A
pT5SeL2hoWGn5R4K1hpSHKJwG22BzsSyEliWRFxjiYhg9aBwKsGHU6s9N2gCVxHYG7WxTrfr5URa
zWFjjWU57lIN/2RB0SaxlHlLUAAt7r1G18CwTWTC5tW7yjbJdObiV6bO0D05AXuSM2z3IczKcK26
717yaHVJ8zYXhqTgPLlZ2rADHNXeDN6qWzSTheLAAbMJQGGB1qQfJ5AQ2SVQmh/FI0sUUJ9eeq3j
t8EpGfScSc3ZXbxAkM/qGNFKD08dSniteck404uwFMH+Sgp23i3lFf5wig+YEbDmowi1TDvC5G+1
CZMbzvSKnVcC5MXG5ofss5F7vbdp3JqVo8pMLJ/u+Zq5QHLoHWW+jlhjDF3FP8advURN+XWTeaLo
QV1VsaEdkVA5pPPvIIEh0p1rNEG+T5rW50G8g9ccAkQrexW0EXQHXabJ1OgvinGHD8StAoo0rbMm
NSF0z7p2Q0AjWRxKB7yPxj+V9coJPy5qKjgi8uQD0eBFQ9WLC90AqrgU4S5e9MVUn6KyzNCWMh18
6L2fYocMukYfnRVYwXsg1X0owiwC/nbncAZzg/MW8nKgWVfAakcDmr+gIfoi8XGtRHma1SGJzyQy
qhRPX8kSrz2UQ9XBADKibiaZFkdWaupykT/+xMyEYnCu7R+oazslI179rcGhH/F8peisyW3u16DC
rnoXjjixcus1mGGYVZmQQf/nZz3xBhwfdb21UDoIAXI3rSyuZBqIr9pOjoPkV92MiF93/C7rNluZ
gn811SgfhT6HU3fGK9haxis9JaO45hsrXZt98Hv71ntxzRXG6LTxgTrjdOc77UN+JxiQfnzszNvI
rJx63T/9u7Okn6FSl/mxLZYwuqZ8ALNZ4u79Fl8IhSt43fv/hY3JhnxnEGD0IrD1MAfl4G2W46qV
Vo9gdUEESGyB88G4Zb98dLlqInRZLeXsZ6eXxOguWhMjgJNUzTIFmdxTA06c1SleZSiv+rJZC6p0
j+ILLOGDC0FMSwNMzArijnLOmbNtG0Z9AS0x98/V38jZYa99JFgRwdCXC5mE0Siz2l1CDGD4A2Lz
TTVxCF7eqikbTM5yBi47kuU0PrHGCv1uel9zR4vQ13QLm0KiuBdVg3utaaBNgSO3zyJ5hlJ53che
YBvbq7MFN2ySfNN+5GhMjS4Ma5i35M3uDlDSYg26R8nH7391IxGc7/NPfPVaP5aBdwqE7Ai2I6pi
kjNY8Cy8zIZPRoZcX8amZeASNdHMWzEQ64SNzml0ODPF2XVnxXw9mtak05LjReN7qKZTYAHQ6RT3
JIvO7dYKMvnwOyjDd1kanR/yPTg4pbfiuXdMVvniWqW+kZjiEqf01YVNYcLsX16ug1+CxWtEX3de
vHIhfK6F10bXfWCVNaAG+c/8eOIg9loSVNzgj8fjXD07IrM/0nOSB6f+c92xG2pwY6wpP5g5f1ZZ
qu+JAvj6GxAFvvxF6NtEhDHxeJlxOAD8MHMFL2/69rAUt8r1S/UfL3nl3hmFarlV4vBgcAjX2ON8
nFqbIIrsga0AAnYWcRmFOQ0PwLhmgR3nJlHeE0EnHCrK0b1Bc5DlEPxqdLIQ/jzP1Lv1ph8dLGS0
E2CI6ly7CUejNkKBTPgsHVY3gF7GtBELR+gxIz962q6JWATpuyylJkbAU1sfQ4/hANSM7REpTF/E
IKdhPnNp71kUexf31ADnkdGn1hVRWIMLE3rYQSl14HTy/ZNvnA1k/ZPq2X8d7cevw6vUsFKoG75b
bA/ErMaSHnZvgEmmzwh7XaiYJZTtS1ojczuvYH6Dcskl7J6gRjPmr402RPYGGG1lAg7lZOfsN8El
CEUuJSO0CmrVB1BQWWidIPkcZJgeHSqu/c9htpQ0P9W5Fdde/v7/h1l/IsO5INvbHjLmIEItYSa9
Lca+phDhb+amBfhgKynS0189ujCofoD14Dl0HPS/xpn1nJ+CAr/xda/eGuc37rwWtt9QKFlDBcUs
+Hg5NjYO5/enKxsMpxeAb/KPVuGvmvTwpJgsd3hdfpllfUoIdpucB+KzIiH9FV2hk9Nt5KBeFhvV
HtTC8gP9m65L7Ht17QZFDTveuNmqx1shgTSAReV96SALCyWIEujb3+qIQb+EbU70XHUP1KaEeZPU
J1NC8NEKDMRo7HpOASCvugNcP0mPtkojrkh8eDVcmjF6OLNrP2d0emANDe4RaVrNFnOwg+rdNCu9
lPKO2vScmjSAXpj2879vo0BMXvsxm2JdJ1eKkexEs6Vw7i3NuKpgROmHlclXGD6XsDP/UF/AS0Ls
n14goL4nNfaCTjU1BSG3ieD8V7eljm9ICpK5vZ6mS2xr4eVDogNjFlyN+1SxjwTwS60zgHs7z6Mu
dTY/JuJKJf5UKiuL1yHtj4Qao3Ei33B4SzK6unsAJ4JHXzYl10IOa1bZ8lSgY8SHpXCgdoZ2olMz
vHK05L8Q3xUYJK+KVhWsENPr78xrZ5uygVOmrUw5KhkY7kcPa6d+mIjIqKkuGw5DQ1CSBPyFu8r/
/m5YBAzs/FSf5DD+KFdFLEyhxgJvNwCFnqnwzgC8SRCXaHXydWN/bBhEALsyBLI7xWCp19Nm7sd9
42aULjjL4TVH/9lU9k4QRFGKsSuuDMhhpQ2LKWqEPP/ndjbGs0q69Fy8oYiIJj3sLclII26Dofbh
AOiwAUQwyEhRV782JQGV/fEth+QGthxS5nlu0zP82wFqK8smEq6AKWsfJ08M8FQGvdom/t4PpF0E
ExkE6NII0WypzeMIFwlQ7BrbJe1ubdNKOuNWsbUJtH0gWCJAGX9oFlw6ipLGXjGIcNMoOr5ne/35
oax+SSpG6kQ19jlYfCYSXyGLdq+GXBkTLeM5n0X44XiKQdM+RzqsP/A9+fgWl9fqGQLH6JENhxgK
+03GQEaZnfjNij8037deCV4UojVcxnKJC5njbeVzD9XwiV664gjR9VJOxka7fe5ws2tWcOaP1JVr
7GybqeLhR4/q6b4cvAaPWC1dNet8Jig6JIKZiRCStDnsyCmsMqTlkPcQb8YJTqrAUmek6x+rvGQZ
e690Pn0lJO5YwRYY4asw0NXGumrfXbxI+4bjMEMFFpiZ/aeGamvH5M8LqoLBstUQWpUwCM93bE70
u/PzEXXJRV1RRBj+crnVhpCWa6ITXttf0kB14CZJshHre4DyUa7EXj6O6D52gc3g/cepqpjUfnsU
RcA2XiPS4rPNcvmoUVuTN1ZTvsv2ml9HQusjuXZIzMWv5W+cc9UPBf8PAzyLSxeBUdF6kOtYQ0Wg
9xPAjpm5MY9+n93uj7EY+gKgArFyvegM4jmKt7ffR3LgrxVUQbfSE/cv1BBFF0EJunWnSnvqibed
Y5Q6u5ADos+1/JuYcn6YwpMf28Z7ht+1wcqFK0SPReRBjjvbf7NtCQbcACSC1Pzpwb0QQ1AuZr6J
xE06lFMbyj5X3i+o+Ux/ZW9GDZQFmkoL6t2ds3nPigaj7eO9Qvv1xYHe7W8p4SWr0otpCV2pA4jx
mF7FGHhMrp+nJCfbdR33/QG75nl/RHkqPN6pjBW/ztoSn+2fCK9zYZxd1yffLEt/42HS5yJ1M08h
6wCuG9tLnlL2t3y2mUkP5kQsIOGUdsyDJ5+S70PFZ9hzerv2n5Y2FeW2N2w4TeT8gVyAh751AECs
L5TgQUVNkCn+KBvcEWOe5H9q4shfJvQAdpRrbJ4g7rpFT0yDfg7n2nquIIQOk4x0iusjhVTFmT+q
/jnNl2K7pF6C3doE6uXki5yI6P9oLMOdSvaLBERQWoRqOvqh8fT3ms7fdpwhDMnthZnPW/gKjYfk
mxCuq9/mcovEUSQdfEwJTxajpOS69eUNaafpMvCvrkbOadfLnh7klBIPP6j3lTgf+D1ZFuOn6fhC
E7FnvNar82IJWZK50DrwZfInwfgyOXBmuJ0bQGcYCTFLdcFNB5EXHF1wHSfX77bzZ2SLAVT0Uref
oXqwuhYK+wuEjaQoX6KtCx+prP4MGTqTiKtTEn3mlNzB4k+DhIckwwVUc46iZ/rAhyK39u9KUali
7WnGLvyCMvowbar4dD4jpLgxWvNWQcnZP2PjIWTn7ZNUosevTGsNpiRFaF/uTnVPIsQY/4hUyO42
0k6myjkloBazf8jhVcbG0Qk4uiucR3OeTDhBIxAobYr0OQtVXeoOxMVq1YsC9ei3wjAmEl4cvAeJ
OFhpTJOYXBuy77xbr7smyrqyjQ3aO6z6xfBaVD9x/wVT/FMRlqhi7VFk6/K5uIUjVGvVtAYWpBFu
dgSfpV6WUD9PPTPOTQNVHRlKl3P/YKc+H8Oq41qlo2ys5S/IWc8G9fQIqJgiVNLJh9VnupXLY9PI
GzXc0BGkx/TqYV7hcw8Yp/wnNmP4T5CFq+UvPbamf7kryB5vqYONC69eDAyRMIeEBndEeSI1g6p3
k8Wf+LpUD2f8Ihoc/ay3Y/7ipah0NLRn47ITqylGDoa52K3+8uKMW7lZCfVcwyt4FgsB4rfc6lx3
a3me2/CByphvWqQatPOTsyiH7WYEoEY8R/SHc2KWpqcGxna6dp+QAOQKHwHkKKIgUVspahvO28et
E44kyVvzaU5zsOhC4PFK0mqryBYGUOjxsUm1iNTI5/0ZS2Fu0pAKDiVyKIJk+4rocvOlEHZ6Dj1G
AMNhwHOljKg81ao+eOQWKa+YXvGat8/uclSGYyUuLNf+j4Vpe4B67zG4O+3ocijxxDgzSsDBAGFP
K2b9aCeeAripq/wiAkQtd/Rnn6xFrXvuFtmgaxqF/oFbmFIl75gwsjZENhYnO44z+kPnlsqBb5dw
QRlSqFIz+9pGpGedZgf+AqYr34GmahbdrE6b+EzjtBys9F/xiS2JkBRtaNzcIH4wybTEUHCFV4KL
AUkBbik5ZwU/xDAeJfMDL7VELSc55EoCyUIEe2AvY2gcrJZ8gECKpwaDftIzK8jy6o9507+LTzbz
/Buh5RPT1bKNSdC2tHZJQNOLL0cLA7kI2uFFBy74PYn+9Zl9G3NGmCyh8J17OVj8JkirlLbLvRWw
o6Og5EI19g56VsniTCB0zDnXx09XnKqrq6tknA83blMCvdpRmAY7OYuDGkYBhzb7f3d45ffzu27U
ICW1c2lmlBMW80gkWgJOcYwcs/CjaX5+/e0MHbeAjwEy58gEB6i/3ZKe2nsDTybnJJzXuaYIl+dr
QoygC/AZqDtWB6KnWxt7qF51uM/CdvjMq0dBOwTGzuqetW37TxPo6kC490vdOFZb66y87u2N2In0
9v+IvGZ/REuGQhRWnaC5jirWNnAwXvo+8+FLXOcEINCuOHGCARj3S7jXRv3NkAvOFmfK4GI31R7q
XyaBuvLDV0WEZMIRctuGJcSu05xK6OCCaAULKhxXgTWJmqB84YUdWuCgOf2o4jzzD6Tjy2sUTmDs
CMicpARG++S1N9k+q/HDjNz9zjiRe+ntrJoP0D9ZNJhthxFphpT/vEmdyQhE3T+/PzUmxinhgfUV
staQyTwJUYIHRk/osVr3xOOYwyUfHD5dsKeDG4FSF4JTURskhpscM55+VMYD4tZ5sXlv0Yoi1H/R
zr/sqJbB54kmNRPooSfWCpTuK0bY5049rcOxuB5BmgqiE3DaNEMxh+9RXT4YWHmPm/F9HDJJcC/N
6A2u2luD2gI6SP9QSSuw5Q6AQJvXVm/t3pkJffjhNOoctvlgHHNDwr+qYas3s4YlAWSobb4xWgIj
pyFMRmHq8vwqL9QnoMbZvnfS3zam3ed1i6p0fpd/bqz/aWqSR+nFV1jYoEDnQMS5ZbRgx310fdHR
yrFms/xqzzviM97GApROlBTZFebflnjB4CJrOCx1KuI8r+l0TVUgHA4QyJuOaEG2oicsH1gQhDVS
DZDtVkFHXr1p0FZnY0RQPDQpdp75dXDbQ9JG3eCtBmH4pMgRuD3Xr9gujEHkNBPWBt66gqZDNhSO
hPI6Afq3z6/kbAO1p1zHQBOy4KF1tHyCjZ6uAw/L80q40q7Few+yCJB8BIBdNxkqxmTpdEh1mRTh
FuhsCyB64bQsH/409vo+mzSRWAOJZz/zSXzNGnHcDlqyJeR9bpGbZEbic/McXxJ+G6bzl374nGAt
UOGQNuXVxYTejyStOFYa5bdfBT2rpaIC7qiztuN7BGl43XRxVVDWTZNzIdw4XAFFRf/Nao/7wXLT
PuEzcuyqYGqGKNRUke0TwPraHzoMFtS3K326xRbQ9MSP2khZbSk7EGnX0h88VPMlohyYAg9NhjcI
P8k1B38oIUCGZgsLTjYYMW12/emb53zzz2CHvEywiLQA2Ij1zJkgGnUzuJhKxo5HQ0FEs+9cxSvN
9t4lR2jxQUKz9Anw8QwjBwdR1UF9OwJ5fmzL5ETKrXQ5Ld7eztNluLyS1C9tnoKNIWD67tXiMkvm
yQYnucVbNvOFDsSjrp9UEK8mQHBbtWWRD3d9DehYNuAxvWdIr3POK5eOfE5IoypKb6Fc5SdHjDj6
5GUWqvzPcyX4G8uOai9Z7b9O0z666Wd716hsxFhxMcAacIT8nTMzsk1/MR+dEgn6tjeVFnw99Vuo
c1zJ16UFHNlCesJ7wPH2bgt1CfUBzXuRIxY0GCMUGAite+JqMgV/oqc1TAll58pAGZjn77Yc5cSv
OG0x/yZFPoTXWi2/Y3+3ug3SC6pgP3YbjQ0QTgCF+IzAZRX74NQBfgErjjtmRpe6gRD7unbNIN0o
Q+PoJiyAf6ZSWSQ5mboIRIgCpSeY3Ns8zW1zEhWNk+zrQJtiFFCgcuEFmP0kpN3qtZGD/dlqU+ik
X8tVa2Jnnx9TbhAjYPV6J7Weyf+/88Xbi+Pmnrt8Pn95O00Sya2G4Jc/eOgr69vInTP+1KUxUMHN
+szT1JotJiyNi/NClr2EcDrTxXr9W3IY5v8Saveo1A3rAaNpFJLsLWOV8hB3RueQsyGepqBJ1/xJ
SW7MvpkP0Iw/H48PwCNC9OcAA2+E6ZCG8FhlMcZzc6kWpWpTFPfLpcnQIF4D1MEy85qFvrwglQ40
UeSzQyPJDUBfHn3xpoV3jiBkJ3CUU42sEwo1HaNvNTiGjHm94N1NxZTSrVNiyXUNqJuSObPjbpg3
Q2T8Zs+OfURld39+XxD7MfYu/HzJdi/wCsoarWQKiL+R9R85ZM4AlD+tKL3Xim3Fqar/ZCcPIUbg
UNxsI0fA3tY98miQBoGnEpiihXHNp2xte/PAYcUYEfC2A3O0w0vvXd/TOctcFPB6joMOM3l8NLwU
/uhFeFyTa6T/pusZSNwNwGiUGEuyTcnlm/rSNcMlcbjLxv1l5+tGlAB5SUMQ0pNM9M+asZNQgg4P
ppmRHKyouO2Zm0kiS/e7eiVcqLNHFqxc0mMykhFcvlcUSIOc4KcK6nvXL2IHFC2n6b9BxcBaPIdl
YO7uLSimGw2lXVI9duUA4YRwfMpRHS4191fxHQx+1/k8liloHK65WMkBpqsnELD9f9wZ0O66OY7V
pSRfX7Tg1RMlDOH1TFzSPkAbudIfwrXdJjbYLA7xKFXB8qou+c3hzBld0ZesrFLg8aiWlIv+8Hnc
hJ9v/Cq/V7z84C1cb9w8ViMrS9roHXVFjsxRJDJYqrgTbVfxECfIae5Imf2MD2dgkY7yUTzdA8Ql
xLEh3J4LtEY7bSZHfau2gExofXxvw+Re4zGsns2zpqM9KO+IcC9ZBQAzd6ePc1xgEGuv2IO82i9b
39ltC+XIc8zkkWdnGN1WNek/iCAKGRniq0vrameintysN4in+e2cjTBNlVE5m0zLY6eq0NvljG8S
Za7hdh8OZ//0Cnr/oS3ZQbBtCzOzNK7Cgfa89uOB/IIVQ9G56UNS0yJWReIiQIW/xhq04J/sCXcz
cuHRiFYwCafzpwUtHThfkqdK3KReTie3lMoQ4s6jUyEm9JMpqmpy0bchwb9A1Lt1SA8FVQndyB1K
1HMFpy7lUxHwY/0Ji+aigZVIX4+M/jvILecJ8cnSn+Y1u+I51yWEc1Tg/F7/6C30x2YcoPpeQnys
gIg7RvurMtU3WKCzbkAvWP8+g8wF/23jSV9LkGXOgfmJjJM7uw7O/oYyRJXV922US9G27oTztGde
HFzlEtQIq4gNbn4VUcY+YL7ptYbGr+ZXKIgAHb02bi3VZ+Ani7ZKX0qw9lO4InWljbEIZqZhg+SB
6zuHfNzZnV5Ls+JNiGCgYIqzcB1XNfSGeyHGT8gxXMLUT+g9V6Jao5nS5Avbj4MTFpYVmeGbKi3i
czin9mp9+xCHgaF9XpXzhi2+qBnLGGlnk5Tdj+XoOexWSFxKUt0//HSKlwoYv20Tlfb5O/FTXsGE
miokxdJ2oJZE9eb0l5YfYx1GCTsJDfBVkSGGJeclE2guv6EUCnvgLLaJNrWTgPD88v2NdWKlKLnU
VrqDTyfDlHO3LAx6hxOa/GVHvMkzMlhfaQVWq30cofQBzvzjP1nRXyuW5cg8zCD0QWS3gpvj+TtC
KHQx7ZPok/60ivZEnmlSOCAlhb9uRQNSHMzhhXahc9aSU0qmqMJFmdyiESZUnhDVEoI+UCTbuv0B
Ylq5DozIcWX9dozAP8BlnBwXg/StM6YQ+asq1DjmkbCdgSePFU59kDII1lauV7E5v6gHz6KmVRGP
GaVBXj3qJau5zQuJ0Su0tzbo8WxftcOjNEKNjKQR9tCQca62I7j67Yb+MIcMKDeRWbcNjjhwXg+j
SOszz/bhHhGRE+Dr8bFk7uNJ8CuDZ4VMxmzMIFZcKHIvRPRoowPl3PV9GbtnOJ3g2muONTIqpuEf
9jU68bzk1JlGPr9LkVSrQ/jxJ0M0lOMR0vJ8aiEQM16CpJadlzEUGTchWu7F6+tpJL51MkoK8PQk
mTcWr3UlgUJYRZW1jL3vhUktrg8OBTxRiDSS/VBD7sPl44YbckV2V7K98dSytI74Q8jIjLU5v5ID
1xe7/l1BLhAMVZVs4sRk69KCX7TxHUi0L7GVv0KslYvuPgt7ekafjWln7br+sob1KO8JAaz0ssQl
7AeTj+Og35aXmyVxstvrmnSwUHLM8BrzpXHt1+89M6J5Nms59BA8dC10/vpWEqoCQ7cC8aue1qzU
zpQp7bo3/prOeiZOZNfHAAEu413VeIs4uA7ThKubGmMPiCXtcPFFWDaIGQmzsSlqJUXMSHap6G/E
vwiQkYSG4SwLAXlbx4CACWkpKzaEiPPcht8ld383a2M0vJ/1P8tzAXE3t2XfYZ+BkpP4LB6IyIlX
XmSH9x1BEKEZFlydY+H1l/85ssrKGqmfaGP+sFNwwpAXEEw5A77cu3H0lNpShQe/utBFBdL0+Xz3
8nFNcknbU61k+tXrwFjEKAEHoOL02qVe0B0R/HCY43CZFL2Lf0e4AApqR4g4kllzMvx1bkj7fU8o
Atx+wgmiAxp6jFsbnQuOVkGPvpC+ddkT/J7+pTKgi1SoAL5edrRs7miin3+1qCkXtszmvdpGYOuH
LSBQxI9YoY+72Z85NDKht6LV0vi+vW8qMtQZGWiOXJt7SQCmEOhYoZdFgm4bNpPVlXKFt+XQms3g
UKhLSwluH03yE4SxchOh1+emK0MKxEg/VZLzoK3KfqXTI2+s+sdf/DimuMIha+dPlcGJgMjd2sNT
Sy3KjYsnDWGD3nrpnW9wB17HzYk6c/cCdH3Ig9VRNc5WpZd6sZ94H+2KJDYvwPU2662v3CEQM+r2
TRPvFRdaIyGsbq6bRUswzFBdXnOfmmcmRK5B58/gIucj9uGCw0tChnPHJNzsme0aeKLWvnZ7rEan
ay1rfaD1h5I7xJ19TYvYCtSBonXyXJzHDGNkmCycE8Mlt6Rhg9on15lJsyG5CYNfO+Ua4lXP53NU
PKPy7wgbB/5hDla4g+k8hNm1mzcF4cbTORxYcuxN/Bt31phG4LPXkatymc9mN6ipZp6JrSRdgk2C
6OeLlHaJW0qEVWiBZ95tXJM+0wVSWZ0rf4fznP4LmP77l3FSf/Dib8VtTFaje1VGSqCFyNOdIqge
iVa3NyUaHh5zMI3HFBOPpMFFTiCZPxV1axGnLvJcbhuzjiW/qLCJBM3ccdHnv+QdT3BubeYqMo+Y
nGKq1PKwFCzOhalvtd+9J1da8l4AYnoXAFjZblW9OCYMQ5vG9zaYA3z/OPIgEaKkfPCchO89Y//2
ZtADLONMKoEOjJ5i8LUPkqUhDe5/du4vCucdNhe9/L6u2RsoKfhBtZj+6jzr/wiDqMaA4uLG3saG
AfkaDM/f2P4Gc8Pkzwyd8POKlWWHtTei08cfLm0dgRjpPoS88ThwlELxH5rDXnlKj4bZYj1TC54R
RCOY1dbq4ogkMcnTmJPijOCDx0SVDvDwKmUD0YmOrwKLjLBK7D0Nc7lISQGIU+clRqW354nnXP/2
V5ks9hId6+9LD6VF+W8drCI10zMejH6ft50SM/v1IDiP0oLrtxPoLJtCMEOVpOkug4CN0pbEpcU4
efkoPaavgHUPMFPvxeGqdN8nAwTq+AhAJoDCoQLuBC1P7cfJhAiTlwgeUD+hhIgxoIDEl4aKItsf
kWigzUI7+y/Ayl14T3Q+M1d2QFZyJGtvP011OrNf3G67gxn8jbUU4/vWe9ISUfapcpe/Zo3RZZUT
acwTuAwch8ACI90CQ/rM7Fhv0H0hw/fzlFjToCjny0IhTk7Yr4QDnkeFOTWA9l2Hrt3Lug6F2LO3
cGkZWGyGakkOd3CcUXKB7craG9WgIvENqv7AmOjVBT7Bm/MjP/o1fhJnc8YiLMk7yR0/G+6VxrZa
aaPCOK4MospO9DN8l/LR0Zeon3vovnIctz+Vp5279rX3UTWuGcypFUsTMimC9zFLfASRbOKVY2go
LPgBjdVWrommrIjNzF5hYQuBGAUQU9a1FlNfUJdZfieZX/a0l1b3AOgreJrRMB7mEsCt5fht3APs
VI0A5dKkQNBAifDuQjZqiVi0YkQrnEK4mlrJ4+nvw2wYc5JvgNzEuF5EavbcH4U6HY5RWQ6xMGMv
q+TNBayhpGaYEwdw9g7M9DAAod5dL4EXnWx5exW/9ThU8DXImrsOfjot8ze/dDQv02YznoYNzDkn
aqIb8irC3rrK8mJ8ma+DfauyXuuh9tFZmxz1WjDKrEVpenJ55CMxGGe/uIpQkpYdLNY8dnCygQQ5
2ZzTtZsOHf2xJc628BYxaQpWfCssxvhnhflLLCLWCNGXcAFYjHfrzou4OOPN6atzjcDXADCHUm1r
nAb22ZiXYPtHBysNWjPqVKfNLqGjeeG4zr66vjwqp2MM/6cvDYQ7SqcJFDdjEOm8InOFDuZ0LXjA
McfgygJIAUwz2hTqf7SUHFO7ZdVQ6X9Q32u9LyGQ867+fBn3TQtFp0IidauoT9GR6BZQDkOt3QNx
UOsnElPSzpmx3+0MJ59elIr5AdsfDwX7Wq4s7PIjvhHGzOrBBYLE3SkvwsY/Gzuo1lm+k0bpHnQP
pZ7uLPaTkIo7mUrcBlbxUPqF8H7tzfpAJ1pcMGkIlUU6Qb3m6aFzLUgxNdpuvALKnG7VV+HRnjqI
lpduI7rhZQtGzf95kKrnANhi+f57V9RcqU2vIaTQ8d0N5yCDcjIwa4rAptTShaURNkbrylsC+C99
gjhcdKymaWE/ecobOpb9et3IWRgm2LcvdDrJlO/dZBMeu6rTJnqXzJi8UVWwiOLYQxgyvFh9UQio
XXbnS800roAHUBfTc0OCLtQj7QKeUCbiSiS/MjrQN4+2iBg+bTiXtZyjBN4OZFAg2WQ48JPr0+NJ
ebIqpPBZ00zAZTIshSU/EaP910O7lJBxfYaBddq7oqPt7iodUcmiHelFZnzebiJYljie9MlYbeSG
MrXOfu+PWtSfUFqnCzXlkEFbmaFWxIBeGHnQQ8U24FeZ4NXsv7fOHST4wRxqFtDbd+LDPdlKETGj
y4aU05K+dFYFkvMPtRcH7P8vwWWJpg8IBFj+Z2bRJG3f8EIy+d/Gd06Z/n9wjUtowjRG6VpVgHjF
wo5j0NpuED7cNroys8MFmqnP+1IE5pBurOPEbQleZngZwBMjDVACZ3N/JBPyJMcEOE6k55LFa5g/
ODfo9FxAmd2kCZOT6O8VLBeZjeY3xu/oAYy6NR4ooFV2bJUrib13hxPrW2w8FxcRALYJTBXOmjjr
h8Y05BqGlPPLiarIeg3CDqRVgopt8lz6Xbi4phWDiJbqeLQDuBR8V8VImKTJnewKecdczzcTjPfT
gjQ0JK6L/krwpIr241qmwc5wadaq0LozTgPi4mAQFrdPXQqcggk/4It0i9o1IocsVdg5F8BdYlD3
3zeD7EwvjS3b6/lK5EAzKy462ua07rEAIhtIFa0NQxbhcX8dGSiZeaawr2KRne6Qsp7t9aaGeCQL
EQ8DLJSph8kElvCccaTL8oZSiCiyc6H/dw4hA3D04sHOfXtmWpgPVYbs/Iq/VxlWWwjAN2D6S/yN
+tq3nfJ3DtgFmyv8CnY81f36qxV4dxuMdPuDsYpoBObp+FTLjJERh/sbMur9VL17AFEs0Gejdadw
56/duDjpr4nYv4fZn8MV7GCoGVRYiBJYdzJFW8SXo45rUQMJX6CUYmh7VLsKEdV8S9kID/oFIW0c
+nyQe/j83hYRVP6v05pbTqM5xFZfHW9mn1+cLXl02+UGqokOKumB16LkHZtBhBSNoZIkmLLVY5r+
4l6r4A2k/3eaGMafrfEJRRc45OqZrgcMnKPgOiTFooQDJJvznvUOlxLFNorMVSUWi/XcUTYqH646
HVW5KrBYLk6eCn/PHFHJQs+/b33QeZy/dGfk8YVSQoEjSSj/dqOfMJxmg5EHfkH0v7LTxk/NnRhN
GxKiejpqHPZQUgW09mWHsso/IpZW6RRveXPHmYcL8HdJN6wChsN+OWPWYJeywhkDtzn6a3EpxJ8R
SYgbtTx9kMzhOF+eu8NBAKW4WJ4L8tWiIHnD/tdL4AIWeQTUUqyzJLNQzI5zjf6xBf86n0BH62bi
I4Ab3Ewz/IB0HjdPxfHrFC6Lpfduy1eZ6423zKFw0sEFagHR9aFR7V1NUzbNJIG6S3RiOL5RptAT
8SE3QLOxgyYs1lJZwPLFCyYSq24xVnnOhHMjj29tsv7H440uIRmi86I+rSBJymRfPVevFr0rWvSC
iY7tnNXYbi4RoHcVfMId6V7i8eNspS1phEhuPN7Bx9LozGB0+v+En6vaSIYDon2kPvh91Tos5Tzu
tJslSu3t+oAkA8GQ+xO6YBSdjAwx86vd8gtyXsc72vPNNIXyP0lAJwNuutUxP/1B5kZfio9PQ28b
vKDocLfkrVHmdBXFL0Xbq7y+/kNe30WSxXl5kStd209PO6lOEd6TuD5rsRhhFs2YlP0GeW9zZQR2
NwQZG6kViplCCXb0+Fmbq2OOrw45+KecJIMuB0KhjUh9GCPsPHrW+5eQzBvH8+QBrAjm0rkzsmje
SZLnaprhwmEhGBHfi15rwsCTCH60SGqBfjkhsF5nVaHIzGIr0tFaHSfNmdzq1zePzx6vEGss42EJ
w/ViWYeXKYDdIIMBhcS2ha2So0pYoJrqJLKkcHs4nQti6zfbhHXUuRqV9UQbJqrBQPkdMpH27Ns2
kSXjpxCvf3/SvtHra8fPOKkb+0i0/aIzwQHFQILUvOdBvnGk+hLMlvTeTjVM6xew2sjq2KO23p3a
oESH4/7MIyTiogCYyIb1UpGHuDDafyR4QyOvDfCR9Egpe8s6r1UegMFsryQCHaSf85jS3xR2ZLTf
NLr5mMi9qGUhOgvSa6Ugna9khsUCJLQN/EKF8v35mMBeldPS8yZuTTPNfMVfblcy6Z6Ch1w6BYPP
Xh0+A1dvfUCUB1GWWJOQZ9WcGaUh7WZEh16eSbeg3gsIXAAgaGuJPcVD1RuFlDu27Wt9ZhAjXL2Y
Oklz3SoEpGasjf0wZA6OAY7fEpA9S0qlUsjGdqNujhkybV//pGux8gw7w0zJ93mJrMLCt4ljWHHD
/+V2wWHpnZXUXITsizt4SDrbHbFdxNpqpkQQDwH3M7ag4m4pEx6ijRvQHJlxY3DjFG8ScF++0c/d
cK7fvusQ3K4QuFz7eglpzBcw4qianmt0qWt2z02c0fR35lZfU8hQ8fcsqLb3vwbIdVleFIOD0TiF
56Msnpf2G7yPupEloijljHfWRcIUSnLDV3IZtWCxAyhp5Fqwg0Feo80FAR1gLc/LI9wG3yEShH0X
4N22PF5KdfLSzL+jvSRvdJUWsU/g+4d4B54TX3hzZcyvRVYaUPp2ZLPhHRf7Et+T2rftlGPcs8FT
TIh2tTQA8Yx2jRJUhiCwij4xvGgcv6vrpQ7dQf0gkISHn9NbkR9IB70fNdFua3Iw+0HyXr5vcXVV
1dzpSULNCVTL9jIGqOBqWsKOtXVvXZIOmo7ZGK+MDJ39q+Xi4DHHu7ZA0dRpJjaC6Sa8iO63fb/G
49fY9VFn0Fowp2WQlmfvn6vcOv2XCFsOrrCPiZYyxqDFd2yW1nuvlGb+O/jBi7LahxjzWMa6gXzf
r/Ufas23iJf1ngJjHhgyWsCV3GfqziQeF5BESg6ouSEZNNlmVw/+jNpJny0vxBWy3QlpxZigHIZJ
dG5jRrFiLEWHS7GZEvYkidMdnWcw9gfWnnGYqWF+nj6tywNiR2qf9fnpVIaHcwPPo1R40Xc5M6Sq
JuiYRtCui8VFLZiNT6NGE+SLz3zPVg8Mr57ej4EvVDEvdWs9dxVgxg/cOGDM2VAkg1worFF7HRCu
S2CtLA2hvf/pCWwND1b5rER6nd0LSW6gi1PRVZfdKmt3jxD01WUQioDiIUK1FUcwOGNPmKnaIUrt
hScA2l9wiiqLwKo8R7TyhTT+oHU13m6SifMrd1TUp6S9gbaXw87XQGGD8laYsgbthNX61wsmavOW
OJiSjH6tN+7K+6IQA6v/KqO7L2D2EvKJiQRP5bn0yVDJCaQinODDkEyy/XTyjIeMCaHPYGzQhDa9
ptCxzYtq4LpQxJvjvwNlkHvA45wnVmJ4j6R6yEa/1yQAmCngoyCzkUrghXhSk5GQE5/HKygcNF5c
b12xtiJfz16t6dczpivg1YhGIHSpv5AbculB3jMrG9DOdDUEtcOVU4z+Fa/VfKJGmO3xoHW19fty
fEUzyVFAToWqsPM3Yp/PpkSnWbsZZpeu1DYwzK68t27+nqCTiQMFqajf7bNJjlUrCIqPbGPJcjeL
/rg0HIdpSNObeAdOblodg4NMZKU5h6YNevQ5cUtXfL1fbx/K6xRtbtyXN3UjCM9PLd8e2u4gLfkQ
xhsy3ozsVNVbG4PgQNE+9vxrZWNMZrS7nCg6gBf3Kmy2CtbZhHEwPVWgJK2p+AT6Iu4hj7DIi0wj
gU4PFRKT7lljX42I687aFrUWHI6umgfch4ImBZo+GrbYYu7547Qp0Ff0kKtm602d/yOyiBkDNq9r
SOT2kGmUxo/NetGKhL1BKcmUIWHXCn1kZPpWEAh3dZuCWqJoCY10PmRSymDPebn1PMqBI+5o/lYg
GMcHhytPygbMAf5BhQXBMK0epSL2KJtNp+Dk3U6oFtKDyej6kO/7CBV3uBh0WhDgdothUE/A3vBj
jFPIw+6WoPvsq85TrOLb2mniB3nsmjga7RnqxSpn9nT36Tvj0QXx0lnm/x06CTwbnVwc0oSNMsqx
62KuhRICk8Dfs3C+Q9av1Mot2dx3pD+PRH5YDu9a/Cq+sP0YSmZUsaTtwN3yPQ+6JBY++9Ybcc80
axnT00OV0lwLhx/eDYGjK+dVOXp5l3NCmtsEFKIto3d0imFGGI+szexH1eZ1edZyewavqS/Ysxgn
yjA1ZHwEVYqmDWf2pPV+V6J1FNoFZr9upeEY+m5t0KXQx0/CsDv9lsTctzJhQDR6fulSnNkCWK3T
yNJ0WaVWzudSku5ZUXkUjd3Zn64zoVCFoHKntfYtXwEFKb4bfMdeowXgl2rqlWvzAXYAwS00qEq5
kWjYajmZX9aukZXDVdIMR11CFgj3TfrrGNlIwBhCLpTXdKgTLpcL9ca0f3vqse9wdrQQFQnFBdZO
tDLEENUikSe6P5ztEIcdGstlhx5W/fq8U/qfdzTC1FFlEbExnt8yinghhr1jzUHqnb+zKZZklwmk
hDZ9R5RNfmAormvyM39xTyyg0O8jAg7NThYrdp/qk8mBEzv3WKYX72OqR279ZijtoEyujT9J6FnQ
EIf0HIUeRSWx5RAwM5ETVr1RrI6Re668naetw/TFzeYGLlmVSbifsM90/VoWJBpc6m+tro7YU/aX
XtSuTaTYmLz5AjZt9HTSHrbwu37qaieYspxGZ6hEHtW+6YUDPOVUDI5QLwtKyBSIC8MeLa/XqWz5
5qZHS9inKq7Fwx5/+5QZUmBAZipuvuFXBTIB8kpIV4rL7doxBwsh5lwPbr9NEQslMCSnDLyJEuWV
sbPhJEgqXTIzHwdV9ksOUZTUI9ey+b+dsZLjmHTRaEW6ELqdTAe3W2b+t5YpKb8GIoQ9xCURCMWt
A5q2jXiwbOB7na8ntR05B4uGNxDvBKA7WwMtorLaM4ecA6+gAhfsajWTjAC6fAGkN7LPHTmO+6hR
yDPaASmtzj6XVTUrkvsbly0iD3zVJ7GsOhxMwGN1K1Zlgk9sn/reKA2BoKQ6RFnf8+dKWz6pGf3w
DbDbVooADGtIoXCyyVY+mPzXYNRE3N0lc22I7xohlf2KlSYEWg+HAo7x74e+fVCvq/uTwgykUS+R
va2qa7pRwkw/DbFw3EhWO4OSt+OhcKULXVZR3ch499s0zVEFRVQZcpDvoBpRs5BDt1Dop8ETclb4
wVU9wATAQtJzvE/FUHqEgHENBmrrMAZnhngvwfi2UQMotENxQ8IpbPljRshx3r487xbZsgNGLl/j
BpLCouuUt3PSN9gynqjZTkNpIfxE4kppXMRU9D6SaFgqcP/kFkG5wsLcuOK1S8hiwVAeRtIr1qbP
BdLeM6tZgS4BIlwx4BuztLazxm9vmKCHe3WaRxwx6BDNmGQocmBKBlnPvgLK9ltEIh2Oy6QjtFrX
NdvCVuDOX+bPdIaqeJZS+8EMjCzwOoQhTHkl9RRG0q7gaEPy8MIWqsVyiwAHwMMXuv0giSkJ7zGN
NN6cYnbFZ5HA7v59Va0AXQlqbo6Zv/gdqHgUhjoPgGEJkhKT9hAQVlgbkJNBJSjTHkwQj/7QCx3s
9I8RCPz8zwJCsjvYP0x8pTcaqm55SnLvw2jaRizVwkVD1wXDPnrjRwi+YUCvIXN3yVfESRb2Ec0Y
WWs3ihB5L8bkM69ZJ1MnvBPH92k3n54IKGSgFdi9ZHSfTkh2gtxXOEzEyvlWGg33qShTk0dGinlU
/ckD6ket/8MWzd3La0jRWl3BB6eZdo6LdtMweyPucBDIjjBxBybRyuTOZ0+lbrXBp3ksm74hqPTv
V8cDo56h+NFZ87rae/zy+MzykAvq22VUWabJRJpyQns7jnnGPFJikxYpWTCBw77Zanh0DbbbGhlr
e422Rwnl9GGRmvLNSFyBLKT1O7WP5Tg6htnhvVkO8QGCpINVBznMVwFX+o1LI1FJEPpNfaQMeIr3
jZzj7rBwJVUULHCafqBGFzeCEEE84qsw9gKXBSYbZ+Y5cD18tcu7e3O6Zb1g9bLwPykgqFkGqFgr
K8xbME4d0Z2FTpecaUY+vVFjcLfxDtak36LOF7UPbXNa4sLcAt5e4OvKBzvdiaKkCPwmCoSYFOVF
K3MpxsFnATU+qIg1Wcey6j6zOEXpRAFaMtX52clk/+bbicFdhNlOsUtbBANQyzsppMrZi0sNzGMs
WAyF42mQfMFqrb3tJEVtuBglM+vR1lwiro78IALnz0QdWFT5ONjRVzgBAX1H5G+fc3ZtDDLvuDEJ
x7uLvRypalrNDypw+5qH2lY0dtLaeOHHPP7NBIbHDcsAxcboEQcjeC1BnwmKO5FLJ6ek6wuuRfyi
nZZ329UoK21byPNi08uOuRQ0XND4s9wVdXTrVeA5K634DUuBmtN5WfELvSySV8ZZXbyaO6p6HySn
X2juw9DbuDiId5MdMhexNjdZv4hqm1TJ4CnIbPArhRYG9MR1wBsgLW5tY0FweEWqrAGNDOCdB02G
CtLZmVjV+XON8TVow72rlUT2gDDr4YSxY1uSpg4iexeM8uqZ+BBwKVmgThJMYi5DNYL6VRk+13SM
4+lmusagLDHmApbawsl8qLtD9X5tTtmLAxoxiZghtj9KYoWKXIdrV1izN0GsBboFcccogwU992LC
g5tV1KggPiF01nR57YuJHMJcvmwTg6WP0Idtp4ZXzQwBQ+1MuB3m4356eF8YjpqZUjb1BEARRT9e
R5IjnZFb9Dd6Wop982ZgsecOZScbAk+jTh6cVMBl3ytueO0zGC3ZiFgF0WCuMWhFmtd0+XO2Npm3
/BlDzwDb9mfzM5UTX3BIKOEKXR10/WLrNoB8+vE8pAUjvTk706n5HnRi+yANuYJeNJhTAZicUgVe
FUHiueTHoAFEktoFHXFBfC8e8LKBmAoARm+rAvNOqUw7IjazXHkV/EfwjBq/4HmtGQ4Jrwmbei3+
yXzFIjzftTEFoJXzyd1c0SvfJnT0r1QYzytK6XNNjCUFFXFGnJhlRZ4+UUmlY078X64+RD0Xrevl
/JcegvqtsJz8HyTSU03O1XNfv6gHMz1Z8dp0ThEmFJxWKdIxJxEcif4I+S0vouDgahyIDu4NWN3O
5f1Wb+mhH06ksBIXqJmXAgsNdmE9aEnV/j469+nLyrDaUmT5VbXFVssuB1suhsAZ3YiCC5BE5D0R
evHC4gsOMdJHBKs2ezuTSoy4np6VVXRHpN2vBJQMxLNgpcV8W70oFpI/5qeONCDxECflt1eEtHPB
qO6mFZORFU3riEAJyvpuSqDpQyUbLijgG/wYx2UOArpPP2V8n7ewe/eADCU3y1+5luATYNilVV03
+VDPC++SWdnCGUuj10T5Nd5yHCazhP3QRUxpfcmbAzkxtJZ0NU00GjDzmTnDHp7cQQypSxcERyvc
J5nuMGXPfftwscOYKpo4RKRc4RsA1aM2meXaVv6zMAyMd9Q7hq1Mm0qim1AFqd6qxkglV+z187dQ
dpO49KmavTcO90reYXURqcJ4Q5YFD8z2jMUVG+ze9/v7tQbvffiD1EAqLAQCa7iH0bCBxa/ohhWW
0FMZEUtVoYCsEnR/PrEyHgr5UEditvzFc7lEij9VL7PgUS5dSb3U/7XQcsoF39QFAzO0RYvDdaOM
d7K/hXLW1qXS3DDE/jgkvS3mRphxqtke4E0Z+AXNGw/klLyYYKXTcxy+YXQ1gKMt2sl+lx72JB38
TSTn0YmEAeYhI/xfVXA3qYYq0ohG1GIOaZhySYXPAJ7VBk1OUa3Pg+8iPJ965Yf8YEA4KHd2DkzG
7yeFDf2DXK6hkeF1gmQmd6pY7A2Z/3xbQUGrm7ZD95R9FE6MS7VCpjGL9enlBChdq7oyyiz5+/3F
2112LLqGDJOvm9kjX20QpC5tBFMT6VMKdj+491ev/Opdds5HoChhNEFlvVjazMrhKxMiwv5N4XXC
OaaKYBq2mXuiZ4SsiZzbIEg5AC58Lvvsz0kRzLspgEs4iucJGdZkqQGGcCgJlX8FN6hpNqil0Crc
s+rf5JjAGseDBGdgQhQsy7Sk2mz7NodfJdXGl1zq9pV2MxDTU8rNT3XTpAM+Q8X+c7uaLfZSSalm
W1Wqupc2olqNvdi1DzKNfEMbDz7ai28OU9kgFHz9UbI7InLmqNExOqnabYF438AjkvzQ5pfMFkfL
yyU+au8LQOwkhgSuikL6Gu/QYkwA7B6FIp4NTw0lF9srdFl7olPKq+qTQFSl2EfIQNauHcXbY2eW
ZRbE+noMwbx5/0sJxR+qqPZ4kO7stlbIvXhHwiu1lWFDya5VZrTRNDgZnMTUpxQ0OEIRtMvCTPvA
M8iKP6il/S7Rbe9i/RgX/mQA0UfcQizyCYlT7x0X0keHZ01YBXtcNiPlBYWzVqvc9R/LHQ0roLi3
g6mRvjjdOg63fXoc0Ghj9LeCz1yLCVSw0KV63LZOYRswfwAP5/+FcGJ4EfMPS4lKP7ygNpV691k5
X4XTQL1pST9aoAOyprIRhI5PJxBLhiHKn9pUnKCTaFk8eCO90439yWDm6wy0RZj5L1+rhWy+eiB4
7PZj/QsXcK1vHeuMcLZJO2Ib8ogOgLJG8qbqqF/+y9HxiX2x3VRvACCFffrFbFL3wmQZzJzAKuwn
r8Q3yzF6XumX1tx7Q1U/VNCr2+YpFsiQfOHS0N/UuerjiFIJ4/ji/qCRk5/0kkMbz4DS+EoYUQbk
ClSCXNU66EbB2unLbb/TKiO7+RsjiG8qyM8JZNJW+To0zLcLNEcJ3dsZPZatWIcFZswT//syRBHU
Tiu3XbRgpYVucVX5ns01GnltKv7OZqVxA7BfhR34lRGmb1zC6Dqv4ginEdjvqQXIRMjK+07KX/kX
uOBKvbfs49l4NeL/yDm9qrbch5KagFZ/Rhc3JvePaTcYILZp0BRFgqqYgi/beBlq4r7grji3U3df
oT8ubQn6FEQnuyV5WOQ7q2pySSfvn/jytnYg9PoeHBHgxNRPoNZWQts5T5aTjxZmYXKguW/trl9I
rwoshYfYzp1uPQZ0VjIDKxKYDs7HXuNGgW+C4/Di+pWyvd70Ld4NEkSLOMO8p5CP7mATMsOTKKAq
Gtp4XQ2SN6NXwvZ/SevuTniGfdbmbOO4pFfEE434m1n3pHF9BNg8aybrNukBJiI7F2d7qFjGO4lr
H1D96mPvxh5ZSjd9b2mKXbcGscwgPZGwUAM2uGl0A+/6u7qFx9xLU6XxUNPRkW6mhdG+U5MRAa2Q
Oya28prEFzyvRfhM7G0G7T6I5DSZpiRBM+BqSP6KbWMY41a2re8iE6OkwW4ELY7krzsXe8QC81D0
90Wc8PZ78PE3TLokSjOhKfe/nKf+uNWCwX7ypSD2wpN+1hzpsvNrhz+x/G+KPbkAM1QZ80irzn5K
HzpolsV+96nU50eY8TKzJeeOhVOwS1ixV9yavqw4/cVIybbON3ve/EHAUXIWhFSBQS8L9lx9j8nH
gHHAzhgPQ305OSSDQbtM9+KSyMCd4EXZwa2nGvg/FN2HTWOV1hq2pU7Ume0snPjsE/UrEjrgRreY
5pv1CUHvtr5NG9WZnZFZCPt/guHAlIb11sF2uX+Qlo+L0Scuhs0LMPCVScLVx/N8Vpy8tipSxBVc
hDWNoByzBY0eNSYcX18ojpDcZHIWVcJI9Zt55qpVotIbB30oWey8e+6k7aGUre9x6FDdkZie0C5n
D6Lh0u2/q5wWHqqL4Dd3zZJ3M8dN3RBBxHHswLKBjU3+udwTXFraAL98CQ4xSDBGdJK1oBK//xI2
mrM/0EOQLPFpGCCEN4YxIBIhN1uhyShBdXzFjvFZXIT02fS4f9CVaPymUmXqMOdJeQUW8K2qI2Xz
HLPshsdnmfMEoTrXecDUfIxD4oTI8arW8Ntmeh4ndc3+9jyd1Fpc1Iywbm3IZy0zqproFK65ttFG
CQPwDM/7LdFUjOYXOnGC6IPuuc1AaoGaU21yra4Dec5mNPAeOCwJvlWh4xh2fpn5zCpuKZOGny2T
wWvADX7GyAlxaKifP1J0Hf4hqe0zAL5vMNc7acUuTyK0/C/IdR9aD2rPXZzPaRVHT2KK5OSVyqtZ
yDFWcZStDhffKqAxe6NQXcM5LlDy/XB5K7byZQB9nMLH8bihNNuIPs77wovghZ0IjzbjqsqtLn/O
mzmIHokAJo5A4sZnJSN6cjTDNW6uPJuPKhqL1oHX0NUBsqWAwvz57MTYOoX7Oec/7Mr3hdrpl/zc
5bXD4R7IJ5cFouX3MY+d2BLViG9782TflT8tATgnn6WHONtBKAmVnJZi3oP4UqvOF3Xf64nNQDch
N5h4XE431LubYfEC+D4rx+5XL6XkGg9+/NsYNqLVrSj1QBhC4RZp/kbfL50NZQBUtUBOQ8iIYIeg
dyoBIey3hyvzKHyQUPwf07/ixx7hvJTysTSrBlldNy2pzcBCJpxRDOKL02mPbsi7cW50w6+gUMpS
bY92hUvGKJS6F2Y7aWAaKvfv8a8liMv7ZiZ4XQ/KWgwtpSN1h9Z9PaKkVphTHdkUJNwd/CFv1TA+
IlTfHfeSkCM94XAB1cBiMu/oIqRK4wRcEG6TdDdJbBFvyhQBZhS+evqxrCIc0whf37R8asvuFGd6
3JOSxRfwWv9CZWtB2Rr1AmQKGe2ZNkTOnq2weOL4GSkRr+GtAz5C1NTLZ1/iaAMKOBSRZp6PoCC2
MWTbuAO5vNll2hgC6f9qIThfBm9ujHxRejXwKWB3EtyeuGHuhmlbC60YbYxdNcqtNrSqgriOjL4c
9U7kb0I540e3bCiLjtUk8fX221ngd7cKXB1DeFx8gTdVHavqhQ3hMFGK5KhW2TEwI0Upfp0f0fwh
dgmF5BnTEQb3vOVTSE3vWBcuMIDuDQlMJ3K+IySMfq7wfaDRTIcMjOwUeCreUYnmJeuBcsm8CirC
IGw4VPPkAYo1Lt3VyudkIqtOU/rAyOqpZzp4QYVXhtaTJH9BRE6H8GE0xHLCLyHJvZECrOWyEz8f
gKozizU1F8l7dm88iU1ZS5zv92YZ7f4+0CMNqcLPpbHvBtxIs5hU7y7kuHD6lu1kVyYKJgAT/jFv
NuzufcQvg76gbmw/D7rYGPtd+EiLEKWOvi1ID5hP3JWPQNC+4Y3TBR+AOEldOamFax5zVHCZwTlY
TGo6Hv7/6qTngWz12YiMc4R5QIAVpa5Xj+BeVcO+qbFuXBzpAvL6iQqV/+Sutl+iCybK0BABPJWQ
pGi2GTJ+4eXjY+9y3eVP+RPRGVRWREQWq9BA3C7LhyWxAyUihHGvXL6KQLTfeBifpyye71xbm7tU
J+hPjQuomOWVK97nkZqk5UQD7VvJdSow/8PGFMS5ncISXZ6KLTHRDbkBfcepnprXq9USykn3hojK
aB5Ju92qG9ictzwju+ldcJ1ZDdFLBJJSyYfNHb6KQ3qleRMtUmjk8FQBfYV5kH2nWLKzqoErruf6
foDxJPT8gu4eFBfr83SkN1yPchhMPj0N0vDSLIbSzlj3oVqGUVcOoCsvSCvatkM5/bjZflJ0zL08
IL7gGYoADQtBaXw8Xr1wIODBmpSm8dDZnTux06ybykBniQldKl8S3N7oQbPL/qCwCxN6fL86edX5
03V8uZSI5oixN/rvyPtPYoH3aQXnTdnmjBHUqD5fdnpGc/RrGPpYxxxi02ahmUHca24VblymuWw/
ZU+dmZ9+ZQ8NOb02tQG+MfqDe5F+2B9Ot8PWlna8A6oirsWsg+AVOeZatHKRCUBnjj1TEEYCtJAC
HYfPiM9nbXo3BIAWXo4DMk698EgRHYbcrHdwCeid7QHkfSsB4mFz2QY02e+IISILBtiG/V0T0V2j
F5WbsBQcAwF7EILS5i9xTZ6H6XOjGhWA7npEbBkvpCMhkH4zYZW9KIo0IYpGv93xYPyrORJI7u2U
YHtOGZbaI5oHrJlLj9nHt8dweJomnr5Jyvds40JGcR8aS4PJK6xyYrmJMn4rAbw/zwS8j6rwvC0B
f4jDOWqcMu/A7Nde5827V/G5NdRLJ88p1RHAdJQgiLgbSaxiTug8IKWNuXIBTWQ94xhtsyyVKiqO
8jShsOSRQFOTD/liRl+qon0jrU2pDPtE8srOUbrpvvzOT4Oxwz/JE3epudlKETthCmUlwMx00I5m
cmG+146q9aCn55g+UD0xKzwWdDihmm7UoZRhuTImAvW8jHocrjYbYPu6Nd02Fvoa+F73F2ZGtUBS
+v29mgr8XFd3fMSwZ2sEJelmqAoLzLk8rxXG2IMBIXHTdEydCqOmtGTUavXFc58vTb7SGQyQQI0j
lo9A7SB/sAUd/AfNF0QdUQQrQ6DbvnirTcrusbr/wsnpFBJ0wurJvLZ1vM9aYkWq3hN+/mI/RWm4
NYYa+mFrqllkEy/WKBYm4x+FpcDanhrYDzF8IwvcJ241qWh195Y7OXCnx2kYAYS2RTWrEBulr8sR
9JYGas86fnS2lusmP3DgZ1PfEoBFszCSc7WaZ2xnqX3D3fLdROiOb+2EbIhg4jmsu8pqlQDvohof
lq0mRMf0rSg9JNaFQzrbdUriX+2En+xS3fb4nJSvxzNmm9toPkryIXggdlMiWeaFQ1Eg9ulErbbO
DL/8NB5RtlwzDBjB3joBCfX/t+uEDfSMZ/r2iNQZTnIEihPm1Gs95zNCm+Jar0/veqOCyFuDZpgw
Y0dycWO5f8BZYbxFQZaWV7A0kSK8b2kn855dU+N0lVABsVRbakN7Gf2EM6Evb07XkFtJAqfsblc+
+ZsdTdDB9BLFILmB3Wn0QyBW6dP4yqYB6Q78OLKI4YoeG0dL9airvE4vNeeaOAs3JT9UwnrK5hU2
HFt2cNu+cRVzekmzQleYPLjYHG6HMLdlx/JuasuHTXJgZgZ6nwPgOJ5W3Fiz/P8TaaN+7SQbj3Pl
9KkHycfyC0aGFERA59AHWixjVduWVwE1aaP9ryibmKl3Y4Af7EUqaKhyNKQp4wB/Qw2iIWD9xkpW
58yxhyy56bJpDz2yx+bGKR5uVrzLSHCxGv2TpCIbKKaGL6aBN/uL2cQLkvEsPTyuVDskwThJILdT
e12Jx2MTFBRA61BfDr/sBnvrXg3frD/WuycyjETUdzqrh6b9mMD7+0C0Z15EJHAs/KzNAgXqA569
bTwtlWqaVr8KgMibSghQZJ17vUn2iKUfUF3oFT1ZLbXG/33pyeOcewG3y3tYor4yoy1D9MJUgHfq
SjvMmHGIgT42aU1ESexzyBUA0pJcBgdQYlvVlSzbnpetg5KgC+g/rFLCe9D0gPZdNL2p9KsPXSez
NwFT2qv71xDrf4q0HM4/ei3cbq7tUNhGiu/flQy/TbI06KgNK+4Bp7iSQNIp6SnBuQ3KunC4f9qs
D39iD/hqKTjpGFacHd4wpy5WuNDINdlf7rHtZBsmChf9fLwRMkFwldNxF6HW5dMFoqjUIgWKVMk7
WN2OuWa2wQPXJ+pJHDd/mHcB4D9Cmz0nBSxmF5TuglJ3LaJGY2J1J8xV/zssx9omLD1ZLEXOnlvl
A8M3vIw9N+X9jYV5zvVK2GXTkpIsCdBTRsLtT6nAGBAycl5yXl18WDqH5spyPfK3marfNsXir783
MqQbBqWljsnE6QWBBcFMvSd5O65GUxj0KuYRNgM+QK8vznXx4yxTRSijBJLg/WFZk274v7wJt0ki
qNNi1qO3fHRfkeIVA9PAS9bSaKgfzrv4/gktpFUvS0a4ytBO4+bp8U6cjK9oyM2XYOq83JXnkBHs
/yb0TRrW2ykmgFNKehopXoSplbDK3PkxLQLsAt6stToTY6pzxTaZVfCdp/xMJlPchsUIHy7Y9bdH
sQVLNvDOHkIaL/5KrZTK2R1TFkkjgVCp6KvTuFC0Yn7JDUxO6gFq23AEolHGHQ82YyofkI8d6vtj
gPnhYi1kwJADpCKI/5+CnLvIwkcqTnRa6CjLgU+2gRz52+IbeDJC7qIkgH2/J5XEYt+2DjSnZDRp
FWmkB+1WiE2yDy6wajHYVwPW6cPOpQR75ETXEuPi1RR+h4GBOHQ0W0laRMgclbueukgRMkbPYXqW
rDRZ1zsqqUPNcpZX8TdFLUu8dYVoGaRsCbsGmQi4QFWY9Ay+DL3hMgqCHMVDgZJiUDHlvpBzZLCb
GNUZevhXoXZbQ9elTz7iSskTjf0FBxrs6BA7uY3Z/RkI7O5/1rCS1vj4t+OaRRPfArpBfFG8xm8Y
fpxDxOww+6TqP6AWqOsor4dNeprcgCY01UyIG7E2LGWFbVQtkdwyF6ffQOuCE+q/g4GBvS/HRdLC
OqA9GKC75jgi6hYcZtN1x0xJ9TeSf7202jtEyIiBmdhiLg3eU0MAHmEd5IL5uBap55R4RngaX7pz
RVZjRzsJljNpLNbiZgDpr3nDnWBApxMLr6PUb42EkWqRbNU5YpjkxnR0b+5wGr6xnfH1l8lQ0AyC
QU+Wqg3bJL1z3bYSQuux8U8oIioTO0VO8KMSyqGMLpE2yhKpUEK79hmTVF6tkEaVyhZj/abpx5bm
c6x89JROZI9FUfFZg9qfrcyZl5LdQIko0A6pTmiejdS16RbbzQVa0Xu9Jeh7E5zVY3FiBk2oUEZ8
eqgoEdDD94dGMmgmxag9l1VHjP7nwoim3x7XDFkbUGzT1FGBvyZbDZdwFBqBeYP1SiveR4+sdDmH
wh92us9ebYhkgSTH0tgFMxtBRWjOJ/adPm+pUrbG8kuPs7WaSzzClzgLn7FLsL2XDE8z7akS01aX
m67ncOXShskrRjaFkPRv1crTmZsU0c31T4733uVEr4kK6ghKWw7hnYgFhS0I61xCWHfjUyTNV8V8
r9IUtAmpg0nXFwKWlghhDg6rB6WPxgCiJsmiTKu0w6nFp+ySzEl6fIGhto2amoQ6IHjcDUTwi08t
dv3sAHXtMCQsrQQjoOHKjdS+jj1hprveVWZX1KGNljj9rb220EIYbu1gqmcQT4xP2NxEz9MKPlx+
k86ph9yk5r1/FtIsKfZfM8gY3AVpcvPWSBOiK7up0DRxfu6JZ6vNR+Tt38QF8CVaI+oAhKN4KcEG
CNi5DraVr72+EHJzydz+w1SqYDAgb/8wv1Uu5m9DSp8Pmd+4Q8hXrdNygaPF7xayFhvvECaasnLF
/kOonlq5PU/X/4DR9ZOgmCFy6v9z3p1afBT+5qnOlz21m1WCKNfyxHBLb6QoxSI+CcyD4pe4kcgR
jRgyXhZtJHenIzGaKcnnIpeX2YQ9Wxb4ixu0kJ+yGpmaPxOUPcK/JuLcHWinWWzcCb+ZrTNy2UIz
JxQIdzcTKUybhz/dxImXxlaM1FGn3gboKipNegVnSF5G/m6Yn72RijDeHdbMH9qO6KEGue4AyJnZ
8YqHqRNWElzGWzzj7aj5odggG3S6pop2FYWt+W/SzfJ7EFUG6ViOzyRAsUurWctCA0QJUu/A1IWa
MGwp5ehz7twqQKUjrIAjFNVeO64gYPxlP1MWklwbxAKMXCdCBpfx0BXj7jEy4gziKaPsPWYCEBNi
Dq1OipRvajJiVqtOEkCV627a36Ze6eEBMsCZlx573sY/z9HxmYnN5QlHc4Gt66kW1QDcGsuISyyF
0AG0ZRjfzJMsiHWauIXEItXo405Szy7QOsFYZTjtL8Z2pUQ61RWx0jL5F4GcTH1ewxIjpDdLR0zu
0dSqFKxadYsZNMhW6q6+394lj5qmrsp5EZQZFk394vJSn/ZDvV1Rqij0zBgrcwlQ/W+uidqnzeMj
g2srw9LLkhiWU7Go/XfcNXQyKnAw2bia4dSm1oEq9AvnB8zfgneXQNU9movJk55XpwFQgyTfL9MP
z5K06wKh+vzyqlDI+gSP3sgU4uTmPo6XG0owfvuieV2PvFTN509+FdXJD5QaF60TAEqrA8kQNkZC
RamqXPA2zkXLa6oUAzNCJ6Vce1ulf/WNGR4MDjn4zCxFPh0UfzReTEEenLUFNvoYLG0GpiNSiGgW
nahiqIhlXrRTUVtKL0DAetpQTWJGO6aSOa7vvQgrgeUFxJxNv1tqJv9vxI8Um88X0bku0xU+IEAc
wXUGRqAlDANipBIrwm/f784oot8HzWF+62SvCmL/egCY0baxTTRcAv+m3aMT221Ac9DU3gXXM2Hn
LSm+zuqgASuTlmxt6/y5B6czZCI8QIR4+Cg8U+gW8NlZU87vgAnacoCI0W+YsbdPH6BkavmNjHkq
SM0hd/DrftHV9h+bJ3LlUUfzI88sDkMK/IINmPXw8b00DPiAKQzRl9owmsJzxo450fLCBC1mkjlp
D8sbYIkcGVlrKXPXFQR272bv3nt9AGLV30PdHrMGrt3apokjUGkYMpwl0vcyRfZQeqe7I7K+x3Pz
IsSERBt9JuEkvepa26po4nSuhdobu2+PTKRTz2V5WlXCnKF22eQhaXELQU90fy5I4dZ5emOLoDzN
bVoJ74urmnQ9SY3o79P9/u+ZamOjPXdncSxPM9iZ0Tp0XQbg5dV1bdwyefPZv6qOnDWPvx9p9x24
bFcWYL7AbhBNfYjXf4jgnU2T9aVaC2DF1lfp3RNUPdKQs8gTv286yGWcpq6FsKAEgzqnkjHNIHyY
5IsNc/o/PFkd61Qw+G4zZ+3lHkKqH3cQC53fiP+/yL94IFb3V5XOsh4G+dsOwBbz3PlJhhj+yurx
hEsHYgG9NPaAoEgrFyq3v6A5xytbJmTmjXmMOGTaZAgcZDFCydU/kpbQuYoDCz8m+YxIgIWQQ4sm
5UeM6PT1Iix0BKT144XvyuUvKxXEh0Ngn+g4CBLdrvSpNfGFN5dGOsP4qmk6Pwu6yBlz0cpV0Hyl
qdGpdukxNnzpvMqBjMUkhPkJvBoA7JODCl7agGCqDjHXh6/2+KVP/W8METAPitys9TrmqNNRtiMO
jZAH9/NPVlUDfqpF2UEfyfJw/wUFurBPiKn/S3qiqNGcWDX8s+IfeaG2JMu/uVd9NDpviR/5DKpF
ovobzNgaLG/77pVQUyRkHD8qBA+tSLLOlr/Ti9EQ2J0j0invWvyPoPzfs5i1ZAddxlSE/SLjHUSB
IiLD+MAe8YBQnFDyb78X6AbAD/f89fb2jprwPnfNK3TQBlE+777mzHEW5jdgG+hrgv5M1s+GWzBh
XInnwmRMFJH0N4hRuC+VTlQEbAC9ohNTcV+edP43sDgMuvBxoCwFUR179ZHoPN8u1Tg/fDeG/Bba
tsKsni8KJN+X8IOiWpnS85o1DWRyd53sKQ26wXPSWOIuURgY3OF/gzEQerTANdWU0xYpEpiK6b2A
5iZ/hc34Z3/mpyhKPmco/7oKhZWF5ITognFhE+1ivwFOCTueAUTze+9pwq9QEoICcOqjCPJwlaFH
8lk6D9p6JH3JMw3yf6ayjOrcKs9xK7JasSHlwJspgO9X7nz77yndUlm5pHlxEIfKttEHeye2Ym3i
DeZ/Hvn9mQHCMpzk3B6PAbSmsOSRdnjdmS2/joQzogXhgCjomvzbn9dgWJL/qBxiauRoD+bMz20O
yf8/tFYxK4ot72x9759kAPyoSXHwe39ee0qpMaZk+SH7q/dzAy5uhStu9Z5XZqeLXq826PrPn5Af
osuFhgLuADU+GlrhwjJmIhjG9RaJ4M0G2+13Z2PzRPIZNg6f1DMMBX+xM5DcgnN9hYOn0883HYmi
8DJHWHQBe7pUz23Okr2e13ZFQ7g8L7wGyQNGmL9WMA0yC/NgVCz8CEqS330UHxfeZlBcMRakgN3L
5luda7JK08qyFWmY8z/JywYN2ZyC53O6LqzVzw0ti2zZEunm2oFVD31b13ESAKVeDpIHVI1EMabO
AwKiQgpqf8FrqWauC2aPSp9Dkye+7rMIIqbcOxfaQrIDHHXgewHE21EwRvLNOgTMS1KLuwwVZPYf
+tCNZNkN5nireyjymBlxEafI+fDhZTdKM9ZKfeGL3BX1W5QFAR36O9pR6SgsZoGHX9lzZKGjQgKN
X8PMNECbgNgrnfX3JKCLktnMJYbZtYLhaI4QmZFfuB69sJbc1qQC4iUrVockkuTasQb5QCLD263b
QAB/13b3F4DLYvWgqu60vAL8bu1Ipz6nG4TJ+lvxclgasfAN9NQFpyFSPky/gdWZlKz/MF9JWEDY
n4UHOQxo2mzkKjX5SKh3oXNVMlv8GIR/LVkqE7Bpje41SwXqhdXkwFF3t+7kL1xQgC0K+wBCaCDy
V1BjQuSn9akUPCCPhcf68P4ZMYara9WT8Bcja8c102P9w0sGK7aYilHSpJ+8E/fKUkhDSwnjjKxE
PPNV7975PtxmW9FGyEtP8XQHN3mlQ4ohCM6qg0R9zk57a4m1d62zREZIl+SKwHh+jAKPLGncxLpj
v+ru0G57mv2e0zIqRGcQh7s/XceoxmjITXWY+r07RqbbGFipJ2aqrzYpoCYCfYgrIfs63Id/aUXP
7nRFzlyw+0EaFpd/yDX1I17N4BYRS57/ojvKZ5dGU0lGz72xNA9lta40rTwka88wOFhvfoCRvrkc
VfQq7O6TIIZuOgywjfhh2cObEJFTMGGrMmLcGZcC6IFIo7ZrQZNsPTBcheAJ+l/5BOkruxIl722d
t3pT8iLzYuNnI3jB550ogdcx15TKG+d7qxNeCp6NFUQAozJ7VcGJb+3C6Gr3iuUZVLGv/8lHEGj5
FLCOYyCrm5tQCu3XwcwFHXtq3faHHK/vAxcwJarlLhe8fWp47VEJi7U15DZ7b0Bbwywa1YXnLFWr
E6xfCzr0e+MSM4qea28QXyW7xkUIKXJadZzdjzTBsZRlXiKAypzHH6aS1j6QyOJISuCFKXy9YZIY
e9phSwTtqUvWon2rQe2QJKUkB6WKMPRx2FrQECGbQYw/zJmccnhRNE9myE1qRLGCmK8EYzPzJDmQ
T8al4U7GmwQM/mlh94VnY9kEawarUt+K6KUy8V8ibCUJ+YZABDtvloXywHrPBU/msaorLuCudWla
ZM56LgKWajqCGmVpYc18Ja46SZo4YvrGE0jaD7YQiuQojJHYZJm8ZkqOA4D8zKeDwzyXnl5edLKT
kHlrgodJxgFJ4lPvOazWdLRvHlw5zUe9KerpPpslUZj/tAOYor33CThO4tIIUObbB86C6BMWcCHk
sucFOnaQXGO395n6hvzW2cDIx0O19J281yOnKPKHk/jnlO7EzniseceVI1Kiosy5eNVvOSGlsC6R
N/UMTawVL7IovsuDl+Ol3vI+k/25O74bRVZjLbmTkPkRsngIeyB9FDrSQ2Ud/tmFdi8tJxwLFgeQ
CWFJ78rmvza7HJgZiaAFBSjShmYctZGA+DzLFXTreYYCD0/HVo2naY6iAtCWnWv2GPj+NezU/glS
slWHB1Z5FhDbRpLCCk3bWBJbxzjEjgRcDodjIleD/WLFbLPM9+r7+Fe0ZkIFPs+ARQpNH777hl6z
Lxr2wzSrZ3ykCg9GyL+ukv+1wxBrT+IIJ6Hut3g5jObzhmtOw6h+7ITH7qtV7VK80zTx+IZN4zC3
XYWFB5RYFrv9LeHyBRWhOgHpMdPgnvKDogsfeQ0wxlm+M40Vja88o1OcsAS4GXJMEkA5esCwsbs0
JDOEFwWyPIlobfcqafy4GGwp6m1SUcuIXqs6cjTdJNDidGYvJ58meWyS1szgUVLE1uM0DVcDZFpM
Uw6HkddfLhGsyvycHbD30+uoodGnfNfxfP4U38pO+vjAjOe7KirsV3Fl0Rs6n9uWzIKx0+g1A6Ty
A3y06Q4n8MHNv6sQraf84pBu6X5fhjv6b/V0iOcr3NBp2tGY33hRKpBWeoUL4s6iz/e3k9ChfK21
epPB+0FjqXCUS9rmElG2HAqfUDCHlAXqvSA60AkxmGcCp8BlbJJSsqRofhCJY/QE+75AIBn4udBJ
AR4nVZcFfDlYu2FtmF5gQG/bzQBCD/BDIvUQx5N5E1VA9DIl7aSeLaijo/6uybT/M2E77oHqtpIN
xqmRlulGqUthk4xjWjBZ8iG9jGfaQACsXeqMZrkPObq22OrffvpYNkB3Svi8dxlTjXX4wdq5LP20
ehtQWx749OTl0n/MFprS7Tps8ly8Gfboa9++lkSbDoGbQHJw2VuK/oFYtHXlscm8+EFOn1nizb0w
T5qsqUn6utAdx1fjvw9uMcdDsKJE0l1BCB4fXaYMd89liRVM5J46eVliwxq/gPW1KmwR/azUAg1b
sPHcsWzpN4nhCFxd8o9/ZRrmGzWkPJv5mENrgtoE57SI1ljD6e+UjA5N67+7v872U6tPBzOGs3+R
Bb/tVFNnoPoCPD1ZIbRE7FGhINLwEPaWaLuTP9OMU2XYywdGUDDmLMiTztDvzRtLQHjZaOFEpDGB
UIFj0UAFRjttMhaW/TFAIP3rJ35XStJhfQWwivosQMmRjOUNR8eTQiko9C7auklKKuCullfD4ekZ
jWZK7KSAWv0ZQ6lLGYJPYOp/zw+WILFAQt3XEFQLn1O6wiEF0W5+HSuMrXDB4M81ClsQRabUnsYZ
qJdKu12L2pGqEFPLlQzI6vA3keMMquTYOp+2Rqp4tIUKssqXJEk2xI/X0uH4LxHnuDZqRRGMxlSM
ybnqszU0bTat/N+xPujYED7arZxcqqPsNLtScAAwQ08vdtBsaHY7vv8dqmrMkphiBQvYVgRn0Pgs
3gaAZhwHR+jkYzElnjn5lJo7uij3GI/0gYfMs/dHzW0FLKmGXRBHKlIE2RVZXApq9BRcAlDQIs44
yp+AWOVG0/DNfyNsYJjQA3GWGnhYFDCFtk4uLRlzwdoDU24VcdPHlfHV/FoyBmSNkMsVS0STuz+u
NRLs0Q5TzZ2a3DbyGcRlBQCznQmwP9sMBCeJzsOgmvDTAwVgUWqB/Q1oHCUn66wDbx8MG4BsJqur
fXxXj8Qw54t8OwKX+mDxwLHNRmhtP7UW++wZQXrVg6TKovZIGMEY2yMq11Qc8hj8+D94B9UZCtM7
RlFp2julU/kT+fVgzGH90OSxSZFISpjNyStatF3XEuDphdH80US2EOSl25DCutAyLe2PnX8Ub9gT
zgzHGJ8eCvcqNZq+RT5qZuQb4ca6JDpEd5guEbMN7wn3WwiWHPfGTSqQ8bPhNh5ELR+pzMFRcRdw
Gy0LSjiaQV2Pff6Fj83G5OqvZAMgfiX1q3HePkwTqCcVOB6ahpmN/iscLDF3C5BEqipsR4N3whzq
B7aSMQQnJROaD7XYpykuUIvxHEbuPEhvXX+cxSc2FMfAyrmmSgQHXKnrPO2mMcOGrlGIMAYBe2jE
+JXGvN65fxa3vujn1vVThvVeEkJdND5qbAjle4y4TCWu2UopB49WOqq1Xycn0gd/PDr5rjUBaXYS
UU9IUzoI2WLR1qZYy6Ec0bd0Gq6hbMzW9qJgem1hVGE4+bMBhDO7LL3ju9IPVY/knG0kV8haKdry
UYEFwT0KWlOlTZEl44/fe+2IJJ6jFcu5l3HX5BmpJ2/5AF81OalrYA+hp78iH3DEIy3l4Qii3i85
7o6KjB6te9Uolmd5QskzI9oGy2jDZaThpthGw7WX+DnimqRc+ehAzKFuRSxr6cf50KeEN+EISYR3
IKEy96Gfs72H+jcUdNS7p1/eZsYz4fHJ/pJaPi0m8sMQIdP3O6UH48tSRnVIszov5TdKEHDyvW2A
r7YjJUT/uQCKkQx3dgD6O8ag4Ex9NTDbu49rv3Lrz4WGl5huDHzYf2h0/OPskrOLitstFBzjpglz
JVcoZvAfhBtaB3QoNNVYo5h+NpMjE8NsRWYRtK4GIiaBv14TrkPfy4LkH5iRt98xTnzS8ip7FJl2
TZP1fIYlsqPIFjbyp19XanfiMQJxJc4ej2ZNUeBDRUu+enD6dZO0CByx0DQ3F2mQCOgxm93tbo3H
HIGspNSopmXYvH14ar9Sk67gXvnDtPxUUEpDj4TWhrl3MPAvYUCRxQyVihvFfybbj59hKC+xbdS6
i/d1zxhxq6gJM+IlHDytuehmOzmh4pN/2a0Ypabz4O7SjRhO7d6tt+XajQofoR7CSzkd25iINOUy
EEzIWE1Qvo2TRAOhVA7PyOR53P2uaK78a8VTE1OtoiwGHv75S1sA8S3zgwJ4fL0DFY3lki1791T8
Yb95foxVh9B+2SIdxtPfxoHWoWwYLGeqeln957TZCBmxPwGRnlWDM3vcI55LSUMGKeIm2qp7YSv8
mJdQoop1GWS4nqfYBEQ1PU5tnKhhFmu2O3a1SkZNEL30QaFUL2lfXz70mrR+ALW0uJrvobhYuJdp
XqhlFgLw+KDBD6NQquEAcsmRlz436oqqbDmblJ/PsMIEaJbTUmfRkspYERsU5xaQPBfUqUobD4gM
IZ3ToX/CrBghc0+iPxMu8bC/tbxqgk5kbACYTN/BUx8cGdfKw0DhIwk/Djb+rBL8ikdK4Y/zU/Gw
vt8hVAtg5DJB1vfAvdkMEQsQHJzBlqjctOYbtJcUw5Cd/aQ+MqlblHKnMbYSd6Qpnm5T9MTfgRz0
U0SbZLqBJYXydOfcp9cnpzu27ILbOyRXSIrOGontS3fj2a5MnJDLIOY/NLhaPf5Ocf4gnABuZwOv
QKCeBSsY5j4DKkdiJZUYScIrBDCBRE3NMdUrTgbP6z6MzVSW54RwDQzIey+ETaVEd2v45+zxlNsg
n+q5B5UoIXh3JnLkETUQXhNAby/3kIEOMCx4ZgQXUjbu5s+Wn7iXtIaD7w1FUryx9E4HfVddgZER
JRcg/sxFhtf/V10dFiUNPwed9loJ/s5DkOcgLvcyJTAV/1ESSLpQwZ3srS+8AvjPpMtGj3GE21cA
2n2ujZVJ4TI1znrpXbwtQfyJSBP6SgtO1IdyCak/jrRekHhbH3whtstvYWN2Jz1lfUnG0bvsEBqg
7Xxz/tQBBoZSB91UlxYwAu2JRmYuKdBtWeXjPjNaXiGcR6nIyc6ns2bjbfN/TPhg+tXeQstP9fp0
Dg2ev2rPj91m1b6PGmkHpbkzMMyxxT489PzuCykSapjvmOT1vnYemwcg5AFEVXMrrr1U2Pzfvbll
qDpKED/7CkJbK1SZZHgvgynpTxT+1aaBTngxDKAyfzSDjKBor+64+BTTFcN6P850Fib71ZMjmXSI
4MyI4iTZaxy4E1jcV1b2whRgV9xO63ScJS/u8EL0Yux3xMkSCx9lJyW0nIh4ttUuIAHuBG2mWrWO
t9qh6Vo8Mgm8hG/0dXNYkQIoQGYDdBypYojCoQ+rcSGZc8SJ47lRS9vz0qieA9SZVbweuqILxurU
O8yeS0XClS0XE9FszWyUAqhHyzSBDNpmEH4V9CxiGQXoQ09v39r+Z9vQMz1eRkJ/SeSO/aqrJru/
zPb41rLuwOjyvccRT2bBKMa+pzF9FIAPzp85zE2frcuN4gSd7oqrMr97qKFYfgHteq3W0mjhK8DO
4e/N3bceufILTfBanqqM8LCJUmmQwjbISjKDDrKaLj2UlkO/iV7tu9mkIi/9iEnDNAUACxeoSQg5
ciftq9Al6E1AyPTtpAkV1+SN5oYCi4JgxfEZsssqxy8KqhuSAgohUYgWBQXikY8fEYkIx4gV7tzG
Ho9bfufnqHyU0aTuPRwMkaCTkPbrv4fviz706j4dOiJkU508ibcssTe48DNEKqs3z4r6L4hyKV+a
NawJkJob/eQTZcTha7vP0946WefAyRU4+broHXWhzh8k30fSs6Fqkp8wWH2bREbxrO+ToS2p8+QO
6GPA+wjUEyEtyOK/9inrkEuabXAtADsmoMfVQUhCCmhKuZf0TvNpw+sRCn6NY+pO9Cx5RaQVU9SR
EmpVv+xD+K3w+JbJvoUi1KeYimcR8wBhvlqWmSOpze5twGtelaDNE9rZSfjHjuLJybWYbHS4f+YY
QxajgSSkxfkpmBwoetAw03ucGF/7ILdoaJL4u+1z2U2KazzJWVG2GnGWjFEMzLKxn4LjEf5wxnsJ
A0lmp7AWHYyEjdSs7nR8M7M7EJVS1jzQEc25gFNiPn8CKSBm9C9TF9XKYMWncF+YEgArFocYJidD
TCBQ67rlXNcsIDrrOsK3Mqr6DHi9SA6Dapzk9lAwzFp8kqZAc1wFp/YkBOGXAC17iwIVVf3f4XUH
CLJQKFg6ih4BmVgikWX8CJ1B+PNls7Di9LNan2PPDezpdYFaq3vxe5ljVMw7sr48dTsgi/+WyCBP
5N/CvzGD9MAon8TmwjJtCH3xP2websCCKgtRZ+gFOXx7M9yRl8PdjBKKo0cWa0jeUjgGmMSPrq6P
+WXGxanQ1Cma5ZXk0Op/mYua/S1kYtFgOowwGbg4yGts57EXSudYwJxj2PqKBYzsYI1uVtDf9XLM
OH4VXw+muhQg6biVKDKav4g1THFi+e8jdXw7648ghFcGhS6+e5ynu1LQi8uXHic8nqH1VjKxA6nK
MXTOxms9g3pSFxtHYq0+tjLKRInx4uPWgKCcjNCCLMcPgD4yJB6dJh1Bo1Wq5LhquMJC1+kTWrzH
2QOtr4sw7uUMBZgbDXxpqobQgPMcZOktDmzXLZaGKGZMICoRK6u5EIYUSUgXiJIeIir+uquLg4ki
9E+lV+1o39xwpozcbqB2iZ21VInlI+St9o2b26Q2NjqojFBHkBmw3e4KXonefGEYR104QCj9pRvx
x4ha94uW2/KQrrenIeu0rTiZszT1oWgkHQv4Y1STLhC2iliZrlUnQ7Mrz1oXTcyO5XZMabTuuOAZ
tARbqNMBHUDlkoBAU/B03RMZA6nclEEHwYrVxJAeWZwjfLJW34ejcMDRkJtZYIY6pk8WuHiQ9sQ+
mDkuv0ug8RYHVfB3e5MIXicsR1j7FOq4ypL+kYi12t/SDhnu+V7/neBwevle4JuPbHgRFg8HjrzP
tlWAzEY8v3B+BvUyL37XbSIioqASGKOzQd15s8L8b2h4EkpCxPcHMoYFCvOy9aO3Vy24QTh/Kifa
vwV4B+cFolJYEBa3TykvYVxa3AnCPN4K2wS66zqaDh4VI8AapBa9FYywX18fHtB9Au9T49pypKQ9
RrCSvpaQwpdnSvQq9STeu22cH+tDI7WiPX9qgeeix53nQENHAPHUGS9pfaPaL0wm2WCWMF9p8XJI
Z4iIAfALM1jaePX6KDyKYUFxQgrkMCJChYt87XDJAyw2IVIIyN1JmEp5PloONL5RHHb87uDDiywh
MJVxSc0XKdPneKPtWLZPd+6EAP72BP6vGexsw7/YAXEBnQYjF4rNCGPndpqJ0KNomexBKhMkNm+1
jAoy8PxfSB32EMzczt7ZXif8iTYaHHP89acbAaVnDqG5VZCwLL0AXS/I7EBdzJYNsgqeBSCAcGM0
Vh3bMQGCCHHIb0BLT5EYZiQCvev98rSVqO5dIm3cLHsBSIkklnx0xGw9BKHuTw9djJdkHNgcHB19
6kW4LUA2GjXkWRHI77DSBZcqvWZFcvycSWf90DNAc/6AJRh/MDWaH4XEgAoQMuWBe7Z/ACeiuEWV
SEScDsCjq7T218Lvz1F16yGOhrRN+Bf1Wnb64BVd1V1JCl/j3YZ7dPtCanJRF52+iJE/d8lLobCb
R+MN2xQ+PWVR95n7ejVnR8079TPVGXeEb+Dfb5/YnvhWFZMLOcT8UrDw6JDg4wIwm58vUJeFiYDU
DJcghtglAQUH/NvVP7lE8DFPRODrCoet3Vp1yVPVDr1ytH63zl6imKuFLuk4b45ZRbBX2qk5bhkF
v+yHhEYW5oM1suHDlfkmm2rwNSiMPrzR98iKOTQQE+5ouvG0jWM6WCP0F7ejYDfwfKiTagqEqdbx
Pm1n/FC2TJ9+0rhzPyza9C8n7KxfrAMWi7nBqqbaKgUDd05YKBN96jLbiykjrRD2fdHV3hrS2l8z
cb+RkzPX2Te3x7bnMfCPNbke3D52xKL85H/m7GJUaslOAZ3HL0QDOXwgAuewyRoDQWLeO0OIPr32
I1eL9A+Joh65ZlVZxsu3mg8eSUkcmd7TSzH2yYgQ6gpp8fceoysZFzQr805h5wq7mCq10ZiV9/wM
gfGHp8xbHYsvSGMq7BV97jD9vM51yQNxi1k+jfZf3VE/qaDlxaq0awJvwW5cmlo/ai8LKhjYj2aM
Q+YDBTyyd7siE7icMstsEObYuVLibWeymsCUE0FhVjRWI1gSGNsmu74Hk9rJUuI6iL09391Irvpa
nH6VGVPvyeNBzFIbUJrMn76ZZLmAzMfadp6WgQuUWS45Yndnsx3KEvslY/BlbJ6oNS6ewAZFQOqn
mCtGZX27B4p+x5KHA5NcUZYVnnEAnTH9n5mVb3GM+1nGfTZ+ePGZb6wQaqH6fdDxrcITUTh/tigm
GxxLXHu/WsKq8dLDuGVRNED0dATobebGG4XtklG4FmJ2caFHhbdQojGxK/fHd4SoHuNrYaMGQURO
eR/2+aCqk5nVurrkGRlnUjwYjSKYA7FBApWVORo1PTVNSzRI5tsDW4Qm1+T7q0TZdlNqU4u+eW42
BuL8sKSaBUbNxKVfGAXDf0Zp8neOzDR2YeQMffolkDPT74ZK7q9QWXJoYKi8P+Hl42TCnDnDg2iS
SjezgDItQz7u3ds4Zabl7gxU+MkHsPSvH+4wM7A+5sl64YGPmW3L0xmV1p30LM8DosZ+RwN0ddbu
J7K6vGqOJFpoPj4Dvmw/I30VfKW2fzLfubFAitB9KXlb9bySDwhPN4i18ETcSxbvfsCOwTK8W6Ew
zL3jG+18RYhUK1/AXrwaU/en1DGCBjklbssK9qluXN6ovl39iq2PmQRxMMVYqE2nN2QNURAl2YhA
zblBr/zct3ojbX8auzcytw3xqf2Ffi0I9bPskVTSTogb+gZuKw/GLdsqwN1HaoeCt3FVWtBDYEaE
jwVV7WK2wG3nSMeg4CiNFAUXJSuo8yaJGQwxKNvR7OQsDgbQgZD+3qg7fNBGnKqFV541uVSJkXrL
xQ8WkCyvQO15gGv9z0GYRYgCzielHCc/BiinqXs/152qjcd33Nx5i9P75Br6P7em+cyPQIN4Pwu0
WIOZpy1u18MgLNzl9hhYDkxtD9KcJkVWPS+shb17n8M8/2c3eeNXvMioel3Rorp1unyHlJNh0O8F
s5wE5yTjLsRu5KUTNzf4kfJvyDZM2Xi9DAzDgpJZK1a0dB61JNgnhEQBlxMFgbZTwo+NmU6A283S
If9kV8sVXLGMF/cp0V0sxrP0dQDEv4AuFLlMY8l3b6jO3fkvoJB4BWu/yYI8n2P2m+yvZIvVhtt5
wOx99bRRP1o2YQ/9VRMPU4nob50yrWPbFCtGQ39HEtlShKTvep1+pOC5ViDmxfNxxPz1eKmJj6Dm
APzNUbx9XyddcqtTfbCANhEhkw8hncAwaIWrfxEmwv+xlGtCPU7anL0W8cvWFEVptowDAiI+1/NL
K4tfvihlrKvDd5yjS3PwhiFehQanI5ayyPW1abe4k/P9o7WGSdagYrVoCa45B9YZEgfo5U+shCvr
38yX7RIo5OH3iBr6+OzSZH3ZayAaLsJF7MwZjyYdbtbclWZIa2WGv5wzeZYdGHziwwsxSKvFkXwQ
h5A3xxMYNox47hbRH8ZE/Ni1aMm82lv3YBO8ZYqy6sWpxjhspF1vojk9hQ6XVzEUz1WcnLoDNtuh
A4jrHGMD2o4Bwr4ZgaFf1IqtXaR0VIuI80u1Z5u1WKn9O8/L0H0umqzfP0wkS3Ynfj/X4YJtZzNq
qQVqoqcH7XZUlkHiz5/7eHEYVG05UVgMecfVxAiY3KdzNgdC/53u4bdwsooaqmjtpHHBXL2umFMf
n5LXjVDWryF1+GeoI0/UGr0yNY7d3o6w6EejE86Y09F8uo5W4blruuCdPI9Jw5OHwrvRjLe8yhrV
E7WS7iUzLFT1xippOEM/GX+Zob9hyfWHjHq0u2JSGylE2dP86Botw0IA3cU7NFOhkZDkoLOMZc16
TUNt//b1Kj6yZX6HDIIbl1aVIn2SnsNwJeBJxn9zw5WYaFL0iiiN/AlvdeTnVEfJ+VVZPN4Bx1aJ
CiaAzoGcvhH+ePD2xKlu8gMthXYp+hgkP1QL+hr8MGMUL1hT8xXFJPvvLLlbX1P2lZfs4yvCkWmN
cOGIR6qqOcht3W2hCEiAI0Rwooj9QnK0UbyZ00aFKCdog6xgBIVsUF8Us0Q5HepWx/S6gFPId31p
mBn5ZTdnlP8u8LmxoJWFN+nnT/98h90pT0KPKU5MadaVuP+qXS4A5tbR04AlJI8n6gGF6XL7YR2A
bHOQ6tm+FFYEttdv2T+i+rWqmsKXjuvEkL/IknjkR3mTRivIokmkdUvSHQZL0GeJxuiUFY63IHYa
h9+7v09t5KKi3AKnUUUPMY7ShJRcLinQyPax4Y299yIiIDillhq9zoJEofNnZ4KIJdxfRwZxkB/d
O5FleKE2LVbRXlsGgKS+bBhBW4dwmgR3ZHELMoRlL+eiBmUlomJYo/txXJQENoEC7fMe7XHOqpWl
/iOiUZZAUZc7wZ1TjjBzbsBO0naIgcA8xXgUtp2fkTrlSmYETdAFtQo8dDExN4Cry9Qk3MwlWOoO
QbxGDtCXKSO9tHFWzQSfnbaGR9nzpPM8I5C2xYA1xSsoTeqwO1UBQjfUsC3jP1JOfBJ+m6NekU2a
1gSPvhog0gRD82MsC36wh+XLvZRa9C5vDcA7UX7m7MX4iWdJqjxKR2RIjpMXBA+LgurrprGpoKva
wLzI40Zi+CdyYdFMc9g1wfbW0wVVFx92/5/Vv12c5fTkOldEtfgn0PmLpaIS48NlYwmfcs9uAFPH
adCcD0Yz4JpucAgFpjGdV8CIWmM47ZNTHTIR1uQViYfg0owMxLaL8rcM+oUEOj8c8ytwnM1exMcE
2b0BugQhvz5Idii3B0t3dX6UO3DoE/G0mxwl3/83sHnR6bGZTjVYKvcN2Se5UBbZqghSQuTwVT2n
HHll0+cJ2nToPtgzjse9oyJ0xgpB3cmbyQn3YIqyNzLRiNpS4qj7UfNheos7iJ7PuR+deyy1r0Ny
IMPc7Yi9wqv03kqikdrIeXe12Hh2agUZ0Bz6yydl7Ov0lzNzKhN6vilYEoZ7lj3+uZOwbfThgGJj
UREnoUXuVAThQuUnglGkkfY5tn6yrdzdraEErPF42e+BEc6RY//P356i/WHBQaYMIghqvM80+u+L
CxKIYvq1eqHhHBqBCHPhoXpLR/mEnJ4Reb8Z9eSWeKyd1ZIZfRALeysEcJGsxHaYkVqluy38eY8p
KRk6cH52kP3QGBrNdoZf9fykFHpvf3yr7vSCh79ocF+fO6+RM8OYcaSrR9tgf0WfCfW/2lajhUlv
QxBL1edO2LeP9VjRzqvM74Oo51mdhwkK1qIYt15EDMDPa2ZsRMFp5xUP6vrxVp2BNyL11l6fOhfB
5TimDDlvOvL5U8QcBQSmjenaDUJ6EMHreqqCZSNI1UprZXKpVr2KeEsb057gmDLX1sBMzjsWyRbc
hrQfOv/q2lbPgAQeQZS3YROJ4f0/4x59rP12fHpsheus8sbpy7dxTD2kfRtO6awOK51DmzMtXsJm
7pvV5D0shm/i/oAifHcbd7duMdjf3ar0zcuO3bDpUCJI3dCVmlhPbLAz9Wx6l284z00lR3cmJuxM
Hlx46hzhGHHSC9SVRUPsF7k53uDXtTdCmx45ZR2+8FDYYchxBBZoBTHIlCyfGONy18Fwo28iMIZi
PhlMDl0AX+8xEU7uVngZt9gVGVCZbUcu9rQoifjFAeojmPnD50lLALXo02RZKuoDO00sNElXglK8
Hvti74OVqnFA7PJj4W1D4HOWBRxIHn488oA9c6QSQpTcEVVOZ/dO4LE/G1M2PjbNL0u9mt9+KCUM
DDwCVwvCn0eyrdZgGM/htYRiZBgIxCBdMqOeNihxjP/YaHSw1x7iwjiRNLTbq/SMIL44vu1X81Se
UH9i6YsMCwraoCV1WGFRZzQBl/N9AXxCbZC6uch6f+ozcF7anPThbMB9agp+5Yn4Uezl7Q+WwdRq
hlCvoSITX4oUug3GXFru3FXBr1TYBtMwBCeqSE7EQ7PP0Vvpjcxzhy6X3ayC0n6XF7NSfgQSbIPB
Wy75ii6yGVdX6TIH5yQ93sncYFlkSyLI05ZcR27OnNoAQ/odc7C3hW/L61lKTQlAMX44fjmdstMc
IcqRT76BiUn6cryy+lps5yLQQu96BdS0AdiyNhRujMwfJPafs5oUTgsyygzkBkjPzbwb0Ul5BAzS
dRjDXQP0uyPufa/v7NVqg22zRBLfKyUjAZ6rOZLnTrxJyJMvN6EGkE62YCOAbLPpPSlPjC+9xaD2
FznX3lOj3k2PHzWXDgWBdQjw1TJlpS6NQl127vzNzPSxOv09CRsH57510oB79g3vekcj95gMZVwr
8+seTadh/c0MhoDMaVn3qqDu91MUotLeE32UYbWRI9/9ojZ8rU+XReDFe/27ninXRdkL/Gxy3Tj1
QcrJKah7/WOIUH03T7869Poy8IU8vw/dAmDkfZHdhvi3YeL/OK7EvfQNTsMYJn72iBAbvnGARybJ
wWG/daF6M+PRhZvDP+IiBrkRIIxIHNp1ViEJnhciUyjwUMaH7cYgZSYTk0cf1VdczSpfSww3fSKE
1wUJhJdAr4Pq3wvvHjxCH39Qn8LKiBtzQSuokEDpPkGizzU9X4JWmacy9nJAp+JK7i0OVW2Knxsa
txMrMFMBci1+q0vegyR6rdQnD6rhoiiuT1G+8n54VOMxE9Tiui49dtOqgnlSHJMwFOKIcw2CYqUM
CZaFwjPXNzUfd0qequhyoOPIx5kBWqwhfOLA07c1f9FNAjqChv3R+izJd4+TPgKO2ThySWazjeDV
WoGMYkS7FdkkCOCiszEGuukGL3jKprMyGhF4TzP+SUKFuEv33MYyIlvhEAUTjqACKHgBL5LL5AFy
61ki5WXNtlJQg7CwWU4QOLCBBx86HZWEFSboW3808ynA+y0P/eVbzUk6Pi0tsS/Q91pe2k/jLs7s
X7/8gke4J2fEuOuKwE0hP7jpS6OLF9OWQ0F4QjMUEvHYSJuFbR0Lh7ykSqX7aErFD9SYZ8o22M/b
OqB8L1QixdpImFOgY+FE1yFxlhf0JKckrx/Hh9q+VTRYR3Ai2vtW2QYY6OzUn+05UlHiu3Bm4bZv
/OvI+ZKzcucvTdR7RNdhAHWOpMcDcwz39vs1OUjGlhBrLhAufKILcoWap228IiTBSNP+Z03ByzNX
ssSz8cyutjaHVhPuza16jfg6rI3vd0EMmhPgwdoanHk4wvlSVs4eF7gerawKGuM4COY6A4nlO0S0
ObZGncKZBskm0U9mpB4pJ2v91GQII1WleaGmL8LTEn63QV+ML8SDzheulN93pf3Rww1Aqi4K6BZe
VvPp0GEsxO7ChLoYQlLQhYaZxxRb3Xt9MKz7XtIH3gMDEX2rb4zFsitECt98PNdjrFyeYqBzBh3A
HtLsu7A42/9wRIVfDlW0p2nZdhD2wClJtzYr8Vy8cQopmO/CuDewsWDtPkfbpfJm14paUiBDoOSK
WvuOqEr8PQ0o9PW6WwxvR7QgRU4bqWPbJEY6H0wl4wEitwl0cbSA1y4HWSgjAcsuhKQvXyMXdSOb
WtThz+w68MV+qMiaDzEetaJo7ZlXHsY065jPriyRmUBGxkp/0QXQwe7xvokIMTew5TsemqeZD6IC
CBdP7QETjAmh7Xm9YMu0WAC7pKoohkUppW4S7qYB78v3uATxZVjBAG3l/AG2mdd3b3UIjXuCmQfz
rAbE8VxeE6MQ51e/FYzDb5ca+eh5WwEyk1MC/yEJetKkmDT0aAWgLRi/6wwC20ir7se8E8Bl+pA1
aKqotJl9Bf1VcJvZeGlL463y1qEoCgBTUDF2M+Yf/pD6oWkF067FCdlpqaCCyTBc9rOv/x6uNUQz
GJ9rr2Jw2rKLLNGC6rcA67K1KHE0HYmT+fOjmQD0s3+IQ2MBLPbm577tExbHOY+8ivunP3apYXrs
GGYUM2hZIcoY5yYjYZEyizHPxPUncF0q4Bo+5b+TEva+v07Nte/kMOJ+ZCY1PG8ERCA+WUCKsj/6
YQHHVMGis+8eaXZtWGZc0xa7M+m/s8C6O6vVL4okPXvq0fiVWTjrMGKztjSWhOmLpSH+DmopG324
K6XDo197LmOaxqJ0TXfyrIDEta6BOwclsE4ta5UINuDuo0aISETuIrQewlvggpygMzLopuMDQ/oP
/SsG/BZS+CozsIp1an+bDDzFV73Zhcby0VzhN8EPPdtAhQAQoKjVxQysvPHAr/VQO//WaQtmlLm4
UQX2KMZe1W/rDiOncourx7hTgWV/ijgNoWP6zeWpCR05QNw9mAXlfNC1QmzoSS4EFX670xRx+ryk
QiHLMvoKd2SnjIJVVP6iF7GUSK1CLah9KCNPMhOVRwkZEFMjc/EvDkhu0rBqTq+QdyM7iWKR0QZH
YntaJnU+BCiWg3tvVzzuVjqPVMOrpjEQaUv0M+Ki+zyyvWM2u8QIPIQfuZpyFV8I9gPZvvjvcxD4
XqP+6trPhJoj6HPSMmZdKzYLgTW8oCNoTYSin6+9CqOHq80t7o2tiPwM/UpiWYa+FlRGYJyJNbhK
sr6C3QJeqzxrbkzkZTvJX0/fXW9iIj40n2S6WSHPGscIdywoO+D0sEc/6y8eLYl/34Xy6OIbckIr
pYIk92Fc3RvaHxSVWECuTivW5xQQyRjLARK+Raw+MlEJYz3QoeJI0cMeizX6coQ2PYG2XMDXOLth
dv5X+F0i/ks0Vp2yp3IGNtgSoU/SW2n1Rc4dcaGM2oXn9HWSI/ACH28TPWQWQjpJZE/SQDXayti8
NEety0C4fJsaZ56C6UnI6Wx39O4X+1TIfIuppsOpTv357mN9sQYRrIzW1N3U8NO2YyHBO/m6Z/f3
QxPXhVvuqE8MiNOqjPnKcPvkNbWZG9J217znkSz9x5BIMDi/eNatqHKzepgUjUac1iCP4+bAaJns
uFUYc/uiikhZhdwFaO3cm3EIRd65xr0IfU2KaI0Liq1MuKgR5B9GweJWM3fUtE0gwMFR0RDQRvOW
xvyOOWXJJjU2ps1PINDMpEkawPbmYzgvkjOJFaVrRtOoVkwtHFMVSiRFE/BuAdTwci3YTTG6Ksdo
DmG1i0wwscQubh5jkcuQOjeXce4BRBafYgHjgV8/e+n/RsuWv9dqNSwrrXb+tZCoBBJCiHoSSQJ0
mlbej3G3NjTpidEQ0/fwTfb8Okl1c2lUaoy99W1b4bHkioKgZQs9Cl85WnFJg9h+T9qPrREFBCgH
sMLUD0PJFDlh0zdjAF3TOsy6n1LtPSNLMs0eCLPDNGuoQOYpud4jmuBUxhq/xaC9pXPLpTjHr7RQ
KvdYo596tLtYxUPAOSsKNH5AOt5l9ls/G/I/VT01AN50vcSZSLTvVJKPJN7VeivAddCg0Ycrgor5
p+5VuIB3ZsDoW0a8Jncei0sG9SwiWtEveIzXpMd/dseo4mnfFSf/wAOUgtrt/X92HYWxg6GVaESY
+FwJoq43BQuNb7YqumVVT6jtH/Ex5reAMefolwKywmk63Sng8AT6ph6xCs6LXV6RW0ODefThqmLI
ZziHCpyz5UyWzsHQUFx0cT0THS5NagVDQgK7wH9rvO+wFCGt16mT7kxofV23nZxeKPafos/awqg3
IIBxzPd2MXLQkn3Z6R+oM2nsROZgj9hOM2viOzf6VQe9S0xXOmUOTQ1A/mznviq/nriHkqvSf+Kl
XKTA2d+S1F8UEX0UvTpvlIFEDH9aH1fcL5zf3BJvT9jMV8IOr+sq0cfK+Re5Zbd4bVUIB6B6ZTOq
2Y3E5NliUmOZEO0gwIIcoxvJO+qb1xrU7C9DeIpoknQtbwQgm4O3sHBNjjNevA3DPVEQ47AfdcRk
n4zM7EVuxIWw7JKeLrLEJWHpcqIiysH9Yi4OePI9mSGh31nyQvtL8LmPBb9nseYL2cR+ieFIpG4X
hn+13E6vPEafpg3V61UltiFl8Ja1IUI6GCQu9U7mUakIaH5yc9u6jlIbgUapthg+dwTI2jmAqHkO
0rNbKt7NBUymiVF+AfV66KryTS7lzDk8n4l807a37JV2V5/Mn0HvGcyGnRfNcKrDAsgYLaNaT4MY
jzLIVlfkLy4ePTK/e6av/lhTYVMpSHtcay3PUeGxvWCosDYwMCBf2vb16rHFgL9ptqfGHcdCmOwl
X4TlDzveNjWKM1oPVURAH++1+nPy22GkwU6kUhUpYMWeY493v4cq6hiLkDCRSCYfPYJa/VD2gRdd
RZgjJCq7PdUBtTTueV2EVrpnDbPItATz0ZV57toCNuu23kxAklKDo0q09mSWsSZVTFam8+rSpOfx
PladDlJxanFKlvGCjhqACp/MDGns7UY8mgZaQoLYpHWC6ZxBhmoz8oc00npe+3IgGicZMpB8Iav0
WRq/gxEJZNXHMfEAbKyuqL3XquZunE18Wz/346pPPEGhbQtR3ajCk6gDr9RKbYNcrRNFONN39Qeq
PkJCrLXAt6sJYkRkXzxnTMhJBbmm56FLe5vzPuywQPFU7dThaJkrQgiFqZf6NyMQaDNhnSFVUe14
HE8GpCfvwXu36jWckXPEwTQFyOp+p5isXJbwlLSj9dpu5D9lOmPFa9EP8YYkmsYv4qqU/eY3snKn
BEdnJIFVaYXVXfrFEEXXyxHAaq/mHsXCcX2l5N+9nKhAZMOyaAV2RqJrdWka5M34zG8j0FJKoFTS
juxrIiKp3lmSWHpbHi/gBDgbCjA3cdoJuLvgYJJNoz3pQhScaxSQaiRNOtKlmsOKxum8fpZtkHrO
qCXCULIpoRqWgrkcs8WmWDkPOPFKRK7PdK4MUIeZA+A5S45wwkK6SOnOAUj+6pNyKNFCc7/rlMpE
aEF+fHrGHaF5bu7siJ3unxuIRQTMPvvg0iVEvzb7S1V59F/+H2+RJMNJrc/x1d8dZSlRsDypVcvJ
vYGIx3vyZ5PtMsRYaeHArhruZuJHvu2drAeaIkm+uvoMeQqOuRvTKzQgAHDTAo8ta2Fnp27klFRI
60LeQnBoIUbTOmadm53477olXQGmxrZR81ub73WPKZNxaLjf1cOus7D2bdOQev2/m6rP3k5sB2xA
uDe4lhY8GrOQKdgDOXrJuDExUysB0J1MyEqhizMSkqlVZ7XYw3o3khjsVoHAi1pDyVY0LYP7SbDj
72QMRPIuuEEnDz+8hocPYS8BjFk+13VoQYcJZwEHl3/9DBwuW2oKI5WJ/roEDygTLA5X7D5D8xoI
3JCh8RoIEDwjUM0KzVqnFmO40wj3uK7ySH+TNq6mVXgKqDofIDEKqk1WEYNgnKi0axtSiRUGpH4I
4JL2PSUrvryRz9UNa9SBAHnCg16wF0/BNW9Ubpal2zGkz+glMvBm1Ap8OmqN7KoWhOCX/x1cj/5A
MLHiqu8Zkkc8IOzGKFn8xHkQhVYtm3t3bZsFsI++55lXjmmE0q0m9ZGTbdNcCDiCl4Hd2kS8QVPk
HYyQ9nGAN+gy3wVllQmw4oWGtw8Bqa0NpH9FkrRv0Hop1GWrs50SR+bNZkjHBPPbkTT3DlOCs1i1
h4rMgeSztM5ioPvbkBngqU0r6pYDceV0g5qS9LCC21OrdYeQ4uqj6BGTBV2vJohqnsCbAZFeT7iE
GbMse7amsgL909G8Rzx55G+kAYHAkOGTl8Ehrmh+JUJXBTQZW1QekbZdc0iwJuPrwkyeK+XpFW3X
w2fyXoK0bIsQzz6AEHiz4PUepuo45TquB5uSFaUssNH4Jk7z/tTqyUqs2PGILMgYfozYVCrxJC/c
Ep4sdGOnkFj08+Kl8gkKuaQ6X7vQ6VWqI7zpBZ66QC4liZr0JeI2Aa7FIZ6sMmTjNdrORQlrZtEl
8RXhlWwA8JGf8743qhtsegogT3YykIuFgsQ8cqTBvrXqFsIKh4OBf/wwTdbN3olt9/leh5CocEkd
6WGhRGbPP/QYXmhHhFN9g1IIlXLrDrlbnkd5Ybn09lwa3XnSHEFCs+f2Wphr6yAI8ChSUJZ945Be
dcv+FxZf4tN14UARxgsSNtMoEIspOTwJuwe1K3iosZzlPCA+1glGxad1YzFpe00I5Xwrsp/Q6JZ4
H55eQY2Z9nKU1ysGAIucmrmOTH4xJh5uvFmrY3LGFNBxMMgy5cpUWXJ9C9ZRgLjgTDn8hStqPAh/
jEI/hPuYyya+wCjk8SIrAv92OMmxxARy0IHXypLIClmxa5ku8hbjhoJd6LEQDFL7T+hcgFXVXNjH
MxZyKgieYL3ILbcdznZIvA76CC9rb+xEiycOjYt5CN+tALezMj2rqnFhK0j0z51zWOvRTBLnwt43
rREEBkVhRFV2gr1ttGVGXw/CwiHhrldg+m1Xz4hQ7/a+YVTPYihkG1oy82kt2h7PuOaaAGixIhf3
crTnbiumP/J2hKkDzLA7MVPZ7YbBfMkp8ohwxxM7vqda9VZBc4sjyHDxgbRVHHx4EbPE/hBuLyay
i1OCBx9W+wYyEZptOQsLQHUGj1hqerQI88iELCLzaDs0v8pEsP8OpOAtTQnxVX6EIYUz+AeHVFJI
/qxgr9BY3yBWQcLlJyqAydwE+c4IZJeD/vfdV3osY0BioQGwgsaU+W6Lb8oDfGgc0voQqoENcH7s
m7OusJm/zYxhuQ33R5fo+hZBDZVJHt/NkElIAO1DMVWAGyRkUFVcAyi3IgUTZAqdob9qtzjq7Ffk
bqEnK6+cllPeDdDPY7PcIsJrrG8zDwquh4TfEC5I8ydb9LGCmXKTcrMHs7cHv8FJ4HGs48FNnvKS
sZFtbGHDvLOuYDX4mH+opGerZMEDP2VVfsWc6OD65U79i06zTuoXPZREjnMPnQuonB/9nQ6PhHnJ
rPqK2+/QXevCoRA0i1nn3c1d06lPxi2OkBwsK/umnO5eadxUAtCw3OHZhVqWMQZcAF1FezJZcJEm
NN0PR1l3y9A7LDvbSZZeH0SgLANyl45mVpYYTh5/dvWNK5k+uf/CRAGbFeCmXU43gw/71edyCKyO
0ZmyAK2K3izic4Cp+nxJaj7th42kHayGyG0TUUflwPTCS7X8R4IrUAHqdCxkNfiLan/htUVTTq6s
+Eh1muJd6hNkN+rQi5xMs11uJEC2W/A53aviW6xng7PGocmJ+PPeG9E+Bqi2WDDfQH/Vv6Q8fM1d
Ku3jWoh3cXiUfsoiRa51Zh6ukjnNHeVXjMR8BIJ8kcZhYsULIbj/ct3nE8w7HgOUd+867142Elkm
u5YRfBFY0XEk9a53UqCEdOQHbL4YkFFIBrj7xEQ5rZd08RRDmr/xCTt9URkgMT4sHPYGwGVQPqyq
2AvlnQvw3/EzbO1MOVfLYl5vifhjV5s41DzvnHdHzEdrzEMBJAgYhrEU9fUClKA6hqBhhSX1jvY8
K9sXm4AKSQdItLLbZb9X+86YDkc+NMmMnJVWymoF9UBsQIBy+g1NLWSM+b7c+E2NVRHNQDi7ysfF
NjA5mHjsdvRYj2Rb7C/GWwclMK4vx8iEDTNp3vKL9z2z/MFhbjoBbI+R1CC5zR3uTSAXY8XewUCY
Fi5i2YQ69lwYGxUGcEdFHaVDKx1yS52vf9IAcvfJ9zr22wcH38Ng79okD1qymI/5NmTajFTwITzY
G3OPOiTLeg0Uox/O74wxdWsUhZC0fw+H8anWOSZ9BI5H7aXtrEajP2YFFX3lSeTsEIoJLoP4qa0X
fP11XmSgt6H7RhhrBUE5t/5bHWzkIi+HW7hpv99//MpkjzRtblAjhGvgaUMcn8mU0gCN7FXVBzSM
gEnWNAIkdiuLlesPb2BdeuSPV0Os4aSoev1zogmOm1YAwcxYk87wFbeCQkiPN1YWHp/cLEBEXj5Y
4gs+O+3C7YRAlcH/QE/JAl0kd5YxMIerR48qQFJggGDVMyPMyb4D/qZyahiuCik9r9HsjVW+uTdP
sqGHIDlMKKKWkjwJHdS+tVWum0nG8LjYOMaTw4UyFloXAuAjzub56BMBqF+ST9AVikA3ygEqveEv
E7PaDGehSia2xoZ1tWCRf4kO0sdNvPUAusoEMk7LgKfF1MoLC4rRBH006UOBVIspSyHwd/08ebTq
digc24XsE17mnzdT5WTkgGTwMDae2cFWnGLdkUT/CGzVrTZXDB5Ubk3+z/xu2BBEOQpnp8wrfx2a
1TmUwe952PKR+e5tYAqVrO+DwA5H5mRyw41zRNyCHc/bEpCiFQbJbhPgp9LlBfkcpx2OBoT1bQ6r
xgqZQxEXyFeL3w7+jRdtLtYpaifzDD3FW6llSjMeemnI+k3E7itflzNUlpLIUo1ZsDbkhQk1YrFa
xi4VzgFl8Ii/ZuvoaWpx1GZdmNuDQekKwaXKf1hjpQUlEH5qxwmMG2Q+yVdvEWobqpwa0X1c6hfR
RP6zwToNr78jrRsO6l06yCvO10RGB3H3Qy1HuDOaB3GvY1v5x46GgFw5L3poqYx0rLrwvzLE/fEJ
B41byGEj730GPnZv3euXufzEiWc6szjGaZbfm1C2hqM9kuurXRO2K3wK59q0pIcxmbLxfJN1m0yN
2muCO2GBRMD4KK4TlX0Mn0R2EfpXsl8Elq9nLPeFkwx8XF7JKkki0N1TqnurvnTvSq0rZn6hyT34
LZ5BzroUQ3+K/oXHY2q72LHL/uA7nO91kUFyV3ZSnwdUyMqanBwRBNmiOyFg8C7sUMHpq3x32mUn
miM9D3lRDJpAXhwb8YA8ImlO+Eyn9bwqhRghiPSrZZvMugp+R8g90cpQ3iXtmhmqoFJinbfO25DF
CJu3yGcTdF+Iumv+RDncFJg8RBB9mb2X2BXylsWOpCeoKLw0aMiwo5/BYQ3lihNh8DJ6EeOdcf+j
BB35azse/7xOibEw3AkdjLyUqNbtoPwzlihgJoDy0a9BOrQBq4BmiOyoYt5YtOHZ8JJ0R2L7Jsk2
ngkzbMeLy0kMo220umkW9xEX4Qxmlw3ftZKatFaQX+0ad80Y0m3PmrotL7/Ke5mZbERWJ80u2sFp
x5rEbo8TAuyq/ynuz7Ufox1jT9JXgDu/z5gFJFYr4UFmIeXt2xVvhtXJHfCkhpFgBI13Fs7jgXxf
oZnTcSlyiVi9bWgvj5vhd2NVkrnVLGic3PJp68cq6eM6gnQddmi5VLQZK46vUXRn7lvoA5dA6V1b
44jkZQf/xu/yFLh8nF/dqgImLpajr7U1CIEdEo1OG5R1txys0Lq+A0S8zgsI13HgDZbSeiPYmeGF
Wiqd6hrXhehwjNL5hBHplh4Osohx7bMYoWHTqC7D5F+ameJ5BFRMFwNH2LawIqxa/ioREejwVTJC
Eyp3eURptoQc3jXZlWZUi2dOzfB2zXthA6GeDFRWCjAYOWZ1ePnG32Wy90Hu4JB4GwXi2zEyUvbX
B70zZrDNINQQVZ1L+nPESAK65Xyq20aDy57pjDrOmWZ4CeIZ2da/xzaPIUGSmsBYW2NIBD2pSa8j
kyEAXy/y+2IqfD1JYy4MfOeaJL1/ZOZ4c8ihNChd1F5aArxnmTHkVqMxIGxiVxNsMNzDdkgssDGj
Dr/OTd6z4XN9xItwaTXemD1dyoSj2y2ZQkvY6AvbJU/c85XSCJTz6KeuZQeq6q56RFHA0nJIJxZ9
JzC7PdH1kETxDoHzgEbBWgyImIk/ABPo055QdjF2vlMbLaO53BIPHfIYvCuiuj6kPKDhhfMmSTZr
Qv9E8waomiNG3u84fhlhY/zjSU+slagVuu0NggZ7AdBD2wLMGqXAk3up3hMMhw3Vw7LraveoSw+l
wdo+LUXwBSy432RyRRDIRqq8Ltk56U0Xdun18TvZ3giUDEjl7BPGQ6VQw8FiOwUcg8tpTSQRq1CM
3R4ZgocPd8XiihC4QaPnsyV3BdhxvIT/M/yvUjv+dLOvyFdH5s3Kn31M811raqSUhkYeFMGWySEM
k0rd5jtrqaqvd9GiNgBq2Qf/4S6ccKRoIEYzmXhK/7+LSb58QhWCQ3pvSn+AGch7X46FJ9ERyDRL
pc4tdeyZ1H3YyWmohrdi9fCaIGzpIR/Mqyh0BmxUx+yG1X35pjv2DwfbVLCL+nU9pXsIz8McdPUH
Ao8AzRrnHLBK2GjL385TfZetzTrQ91lxM6xw4+f1YHHrm8hq+BacBIjs+iJfI1N/kSdehR89dWc/
HuDryAZ6HoNPRQAUfX/WYeA6BaZOgShZOdRFRTyrsxZHqzt3l5PvusFFKQ+yPFJ+JVsK2UMNd2iG
qcrR45JoBkFHGHoYg9ZzcqHtW3SniMEepBVRG8cXWUL35P802KLUcuvIMkL2eeBGabvQz2Vb66sP
W1fUA8i23ULyV+/HItoxdmAAlGh4kBFMZGxlGqKy915HKYNh0kf/OaZoSraaYRaN7q/9hIMhzhSg
GoOTLFaEiDv3M+Q8UGci5PvZmMgP0eHTOGso8xXCHNzOCue1xuBBEk6/BA7uIhS0WN7vTZhVK+Q1
o7AlDCWGQH6aHxFQnPuWdnXuVDYvs6Ad/Z05H2QaS9qwnDUYWVjOfDDg/IReDaSrk2Y8Q3+Q9D5z
3k1Y/42iULxdPfPvTH51WbSISJ8jFBqbM8Vi9gpjXs8DpzRAgwdEBTJlC6PW9AddsTZz8mhPDaSz
Rl3XKfwUZGoFZewbQ+tpBhFN2JvfBZTrl47I/jyMOyxCQ81JR+2meAg7YR4K7yENVHTTeLxQkz4J
S4zlRwfhfsMsKfRbKN8HSVgOLd+9xW3u1jg9e9gLPv1b29PCvPGv+Zo+mhxM7oFO7CV7NRX6QD0v
BWxZsuJJMISm26YHLtF7It+ltWQ0rJ5h2E/jWJJ8ZnV0l5Ok73XYNL7Tc9ZNiscgYg6LlyQOxa9K
x4VotgfXPpxKkVunbzdFYo4dnNEcL4JFUxKWe3UVBdYoR1D9AaQd+x0pqfL5GXtx90EbSSgXexRc
yOUIm/z/aySyYejFhcl1viNnENW1uWQdMn6PTlIv26IhJD4DjL/v6xFYU0r5oNbU8si5nK6ht5OF
RBgOVmmlAD7KIPnhP8N92EiMdubUZpJMrZZuiHBjb6QYpBUN5zTmx9n25ZopCBFyCWvR9g0hsUll
MRM89NoaZz72JkyQNODkl7b3rNprEZZLyb/clo67jYVjlQ+Y7czldJmLR8xpNptDp4Lgn8kGpj6S
LbBomovDmymMCjh4HMOCKi6PsuWTwx+s7wGRq6tQAOY7+Sqx5JK43PjBuiTCkN8w6maJhPkBxx3t
4cjFaXDUBIfvVzD3MGLAK1ytXFhoCbb+ps91tUN31XN+SkZ1E7/bAkda8sgnX7ZoMdDP5lR8r/ON
PxKwK6g93jl/+VVcgv6N70yekz46YbeYg4Dxj6HM0AEom0QZBgFEGgvN2i+b/csF9n/g5EkfF9+U
FFVLeF/wcqbkb+Mz57jzngF4+RinyGxETshLMSU7YFIXBT+tfIOKUihW8T4e0/yOAoDijlXRRC2b
kyuyJM5h7hTQo0rextyMqyoeHGhzqQSv4DfW4XYwW5FgBYhAfrDiS05ePwcZScJD7UA4BlhfoIP6
92og59FKaCdjHYEnYd1TYnyi9shF57/kjgwoZD5K2aQvmmEPqUbLhlXrXLRvOPeYqZvIiB/km86t
G5uECV5f6JwV5Knjy5Di+MMvtHkZNKxXAm0HLWk89qW0vuEf+HdrC2HEwzUik87Xowy/0ppSyG+n
4E7iEJumRQKTCYC1cnrSZtvCIuARDOdsLrfGkUbRF3dSahQhKROJBMgtAU8WTrUzAeNpPqBLMmOU
5eEZcp482k2xzaZs7XL4ZOLCsexTtNWuR14i0eOyspSjFmJgjaAeAdMAklGhuhIw5SUrxm5kWX+K
bWO8INqyMRkGw6CMcEqgcxYO6AQeD4SvFaWj4ITjv2gDjm71Lb02RHHavGQnQySVPsnpxUZ8uXIV
iAvLDMMveZsh9F763FBXQhEXg2KwEUMXwwjVcLvNhV2dLNaRk9oqpWC9jRcZ3UWikAGpXleqQAzq
HdcPcfbfPWr3tM/bHo3qskR6jGFDA320vfLSAdaeMyKZjwDVT4lZUuisCfDm0LMG5gbBLbow5IQN
5g7vXNsTw4ZOzbaXlxU6fVrx2/o2ZdGB/kgUsDKGmzstL1UomEwijP/Wl6kBn1mOigRbonAON9yu
lmI8k13Yfmnl3QXxeMPzXLG36VSBfIwIkGp1C22LrZ5O84CWpgSskbB49B5tLvEe3iQ0OmyMz19+
nECfkzb4bivXHEeIllogt/fmri9d0JDk4wCBZO+BDN85DO3I4EQU7zGEmUSTLHOJWiYViqyNLYON
2e+UxYu8fgpgoCmUew6mxZSoinzJ5IBmVIvWIJSscAPiMVfhlGngQMZb7eWNcdKhckEeYQEZBZU7
IBMtlCd0w68oS4LyfAE5x3QqOEitljNSnn6Pe7wN0HU6DlKfsMSEdmOedETfn4JDnB+isfoKH21n
5bwpUPPhWYde+EnGcVGtpyhp80JokFCoeY4/q6g0c8Mxek8tl/qHCh7Bq29HCsewKaVDMYIsLdMs
ZbtO/0OJzpw8oFRy5H5IjO4Olrix9TyQqclPcfaUj7bqLZVzJpcxrA/+iVIXp4okF1Jv9AqcpJ6D
GB2lTMbDY3IKW5w4hVsq1S+OTkrE2TpBIAKCPyPEHBIUvZsQHTEOQrwgcOCbPM7QJlKyIwgDr0OH
Oyo42NZM1GHKD7/rIC05YClji6rW0azoVsSMHfclQRQJtt7RFFDG5bxP+ffq6otdgpfOgmMKpQUV
zpgCn7o3dwUs0qyNZJmIJlioQcPxyTstorNc+pMtVLjudynkrj5sxQ8+mjQU1cmGhEuxjSO5FUPP
3EyREdXxUYvY6Z0ZE9GtIey+XSsWsuM9wfQiG8pkQNnpLHSkeFANldrWxAg2W0CBgDtPqK6Olm1Q
V5yUSnilgIKSlgN5hgAOb+4bfA3DMedG6zJwjztWgEWJpRY1MlfiAgNfCiAeT2SD33+H+ErBI/Dy
ND8G5MOFQaQPJFsHDk4l9cqMz7sK89FmELQ+xvi9TR4jVrfmF8vs9NarlOibYBBgAnq3/OzZDN8C
WXm5JXzAvblej1TxjwUtX61jJ54M+R8EeElrR4E9rPUzzE4uEnCamMQGOkvNsR5nm6soufrrvt90
jnRcVVN9EetdkcpI8tApTUvpxn4HKJOz4QvjnkEgNCmM2AIZCqGTjrtZ8V/EE8OzmRy/65s1cUu2
Vj3IFyCbRZkERINBWzS2dOFLrIFYW9bsquIjsBNo3svcaXk+RTn6JziOXd6zYvj1h30hWEfOWaDP
lBCVntpHyV0ku6Oyv+yrDRcJ70ot5auivApan75IvkjkqUvGeUBuGJjHzdvxhkJ870z+gPjAWIWd
IkEXFXQe6y1lyyTvroMofrD2pc+FeHFEsn6GOEUAx5kvAxdeSmS0Iv3Als0vaRwKEIqbj7VSIKnH
iJzGrh7b8EoVvP1fA8V6pKu25SUcMhMxN4ZzI7xwjO8ZgzJ4GHVVsDkceorUc0LqYl+HCk2zyyFZ
D4gv+R5fykIHYN4Ij/YS1chJVt9j4c9wWKKRUknVmBBY7PkQ2d6/GRCeZsRyPAkjgXV3jvvAVrPN
SBU35Pk8jj1WcTSH1Un/Y5X60q8mW39J/2MsNyRvEchaTOqBYInm+aqN1JTjlQ+v8BimhTZxgQeu
OlgEDTIKMjfTCNp4EiOmHTJ7TbL+nxDueV3Eqal8pwuYk9sB4EkGdlb+aNeuvNatl1Jk2FZfWz1/
65LbXPcUWBsf+mCudJ2wP/7dOHjMeeqET+5FuJgYHVh1SGzzTVss5LZydg2xpi+nxeD3kHbsUrQD
wST3KMfOlJpMMktnqMOvHoFCVQEI6TVPTVlRcbntkZDNyuDSMEzFfX30dI27UiyzUfCe0FPH3URI
c88yJpv4K3Dabqxk0EcwtohPNs7TPzdiV0EQO/42TIc5txPU8rpo4j/xHKS77ySzGUFVEKxa3Xo9
Ku539wkip96fkJD5IK6DyLL+TYskeQYwnMtE13PU/lwSnGejv51SZB9mf5t34VE3OMwXPpeQHmmk
mEnlQUdWQ3Kky1mHk0luDJNWwjtopiDdOiv/HDAmmEsooQIaWOXAUUVXAYbLKc9ph1cNg8Ab3/Wx
q2v5PIOpkTuclp3OtWtTMxXnlVaiVs4+kvhRRloPzcO8gnx75mDWq1bhO0HADtr2z9AEyKz42COB
EJuc6fuBsnU8DmqvOC2k0itIghEM8qmN/7AaJGWl6A9DUSBkmiVLOrNWylDJFyw4vAMWMtQkH4C+
X3QvPo+O5ZRJYr2xSRXPomAIL6NgJybfFF+pXRNObMIX94j9yRKVguBlfCdEZPB5mkLpxoSKyazJ
PusQVKXpGuAd7/43nurhTDjB6sb7mHuIHRhol99Y8G1Jc97QxZ2JTyCM3zByaJHnX5jRvZFsuKG+
fcYtXMwxOCga66QV/VLkGAWIo46bLC/ku7ukE46Dt4uwpL3Jxdr17HM9h6Q0EywL9BkaKXpMhPw8
4iiJ5XKPIkNQ05rt5kc6invVbDm5vOo7A8eVrUwQkZvpqzE1XPKeW2VdEjuM1V3646UQKjgxYsuT
BWNdMFCgO6g26dRy4YO5UEeC2z0hd3ENQ9VDlz6dGCwNMdiH/pqYb6eSbfG2DzWECRSSzoYABf4N
K2vIFxQZ1NpTVsbmqw9pS+eQdBBtDh3yHBFqZFVUDhG/uV+yQ61b6Gu3SMAkQ+XH7nNJ8RMfG8AK
hTuDgdsIF37JXsciAAQZxCyqaEcyRH+aAmhik5dnLiuqBAq75gC+HjAI8s1WmN/mCa3ibrI8LtLz
c2tHyL/2gkZm8TkL4HkgSRwaj3IZsP24NuTBL2mXSFQZwIbGptaBlUlNRGVQQHFfU2/LgaTLRJId
TPUMql1JifQbqppuGRXhj4RLcijkMB/buk6rIvEKPx9UUNwxp3qYG5jTMt+2v/QKG0trXTPMlFzb
DfhpGGy4SNN7JcO6j+Q3nk5vhAI+viJjrvBzDxxgeo/jfaM6ChShqDSfh5hPXT+Ux9+vRSknlYSX
JpL/csvTxQXyWcc1/LsV/XWyHVZZfVgAmeudp40hxAiuZqdh77ATHoe0UfkJSR09NnugIIEJhWYz
8CKABmNujYAMV9vUF/56xgqux0NLiMcHG4X3zQ31RVr0rL4D62WOEVvlSi7xI2Ii1tErQQm+A7fM
drUsMeffGKm5reFNCsDUapLfCjUzKWAzQ+2bCt5Ca4ZJijeNyUOxAktb1ECLAQ42ZV4Hx3fXr7mX
eujrVGIAbeqjfOeIK+Ikwfxs1MKOhgOPqbNmHDdn3oqYG+mYgbPJRP0t87GbceRLVSVNftNc5Sgk
Oj9Ke4gbiCMsg0gJLdo22ZtIDvIfC2FTM1xoweLGUjMELzwd0IOLTuCc76uTjMgxYL8U++ETH1HH
Y/yGIeTHd0aOBWzj2HBDXm695TAY/11OyX8lx8+R9kB/j4NQ/F5/GSw5lvSVQPS1NbNZy0CFkkvi
ozfNFSz6LEsUL1KA3cMa7kS+31cR5vcYh2BFhdMHSG3+FSFlgm6waFYyjJ4eg8qJwT91ZTObsFao
D76EH9fxWGDaFdxCKqG6Vmd1P+Qx4F+ajV/OVM9FDqJTffROn/pi+meP4qsmFHB2PgHkHypu0O9h
xBVVq0yn8A9waByFqiZ0CGpT9Xu9wLieZbkreqi01ejlzi1wcflSZadW328H0F9AkjoBN6BEkndx
F+MbVQARMXWdT8aeJSZqrWlFrBRiWZDJ/uC+jEiam7/MgIIRe0cBByPbKE/jMq/UoaEPXp9MHyXx
X7TsBrJ3ZMVk0QHJr5GI4aE2SZH8LC+xTheHJftv1LokRBZa5A+GOv4nqw7BlMClINqfYBtnC9YV
3Z6JWhzp0lYuu607rZffgfJOxWjNXiPPIBEHm3yKMdzGmZBiODvZ1IGjaUsqGBbfRQrEjZ+Dgm2u
K6EI9qxLitn52MRDZ+MzRosHgA8VpBhLDSflMhmQuiViuNRlvC6NjwoTxbsiWZ3zSSa1rlzpFe2A
JKYQ21vlH3qAEVe07WZFOzypsaivfuDqVpZo4XqRlaoaMBY+31sEJU3fPQlLfwsbfMNtWgNtrL6k
ESeZ1W0UONulWlxzp7QlWNl2CszvsiVDx1X9p0zhaylVJn+lodSjyHZs8vHZIRQ0eBu4ZqFtgv+O
45vBsQ8IWFM/V1cOagLw0w8t+8eiqSTSQP9/8xRktqer/mhTJc2rFZHqvcBmeL7JNKgX9tm3ldzy
NeqhMCq5D5yEP7XraxWy7AghXVUlwyObFNJGNTGDoeKMS+o6GgTuCbCyhHLK+3Ou78FNRzrxcg+3
yb70F18gYwvlJRE0VTzha8fQXuFUh0Pr/8fT6kRUUbujRggLBAXWzzPhvxXVmLk3P1B5M/aiX7YR
8Id+/g4bRZAtdtxwR+71aHn0f6BsWMVmTXENptj/5gCH3q2LyroDnTCpaveaY6vwxAFUldzoIxlx
EyQqd1KH+pDXbWZ8ZwHhqYmIyG2oS7zENlyDh9qcp8Tym0KB4+41NhrpIGkR4bvQdOr81ZHUJg/j
9vfKiZS56KaXFtQRgfKFUYLG8AWdBEbG5Q3wY1HX3p/FnNZA5+9L0SH8LQvWyLlErYoX/zxaVnSs
MIR6KQquyeiJSGBCbOsUSp+Md599jUJeltb7Dm5YxA9ZwGdNvlBdTMaQFtqoW6HcV6faohQW/NMc
Y4rkzh7x9WgC5vPldYQEv1LqWB8se2BPeDSW76qkIZS02/dfzeYeLX9mxxQU3owlsoiZ3QPfHT2J
HYnCD8zs47gme1kq3jIEVOXwmLmIT89KpJq4vYAv8RfFqjXm+h4xHjsGUs4KkInT2mCMPqPQ1Jwz
2Oy6LNa4UZfdSekehm2VhU8AD7QFRHh5BRb+JbXW7o23SgjTgYKihz/h0xZ+NUh/LTKP3KYV9+bf
456Huk7ybIp8ln/dTFYH+6DGSgeWbgwI0unPBa4SjYFRwaQrXAXQ39J4GwMVcpIgZvRg2Pd+eAbg
IN+a5Vol7SXFYYaoHKXy/RhwScdsnIOplQut759DLrmUIe8qBz62zK2dpX1kh/iImcoVgtLID36w
wTplkFolyFQEzMUEpEbp7E5PsxWDFl7Qyw4S8dNZ1fkwCkWbc+xJaeG6RmTYeAKzq7aVsh622RKC
8Uyswrtt0yZ+OUWVnbu0hPjfqinUSYLFr6lDWTN3nOVk3zpbikY8IaVRPYRu34fupZOumlpnW2sn
CmSaOuVIXCMt4U4Zvl9ptjtqCXlqlcKdksHUDk4VK8pjpxmxfxUkVHDBxjoyTbLUTbgragjNqGPB
D0O3h6tr/EqREGObXBF6cMzJiVkSQfdUKx8ybZl8ZyvkzqmxYOJvCsOR7/DYC3GX4NJZwn9GnlMZ
kgTRgakXD7TTTtre99gXxmmFGB/DdQy6BgnJQukml+Uj021S2cfg6KJCxw873st0QDBhr5jnIflR
PfzCKNYU2O3FF8wj+KZ3BIqFs6tS9VLR60RGVEN7JlwkmBOprmIM+FZnQ+MREpzk5dcwd5UUJG4N
i5QPg3nJjZ37Hg12F0hJji8hr8/Bn4II2kA066wN3p2nKU+Jz99UciBQs7iNGePQFMSL5Ruo0u42
zgWG7uuxj2wt+iAOpeiRlhqFloiZl3n6/h4rZwnlFhl3epAquU7rnC/1sXSWo86TlY0PVYJGmaVO
YN3THnfrV9mEsnngN4RcO0YhpKz3OyJ8wcJpmU8gpd2IdBLfeJxxaRNXIuDdI42T5l6Kq+N4l7jM
0qpEdeylJGDbRJi4puok5QIUIP3V97t/kh9CqjZr1wEUQHICY6wYvYC3W5uZWIJROHwIJmWCJGWy
IeOi4YyrY4Uc6KY7/DhhDZYSKyN135NfhFGUpT2aRydUOMizw1hiosmTAlCnFm54u0BdXZYajfzB
HCBVWlH4eTX5UJ15EU73lRRCoonghWPQyYMr7UTYQo9/Yizv6cO62+FvMJw5pd+cemoYG8wxK5+E
ucrtPwLyPRGwmPRtqqt+bl2XT52ybg60tshlieTQBxQTf2xWPIAF1OLVZL7m1NuaPPV8SMCC38aj
wMbnxbqI9tccV3SnZL34o6MyP2XK+bKrC38n0gmiKbXXXYN67G0uen87PHKUsSDgbzyy+TtS5B+9
/5huLJsHdP+ZxU9siKEzYUEILPHkHEP6QOMdy2jY81q2LjAqS95vPHGokkQI8Z4eHQsLFyfpYXIv
6FVOgHImF01B5wZhMySae4OFRjhdoofADu3UylTu6h6zqLiIT2mR4p0WtdMv6k9nkcjk3BqrnKEn
KCu0lm9JAhvBU7D/dvpruyTC6f9lXn6OAPdAykMuEbRVkGAzlh7O7cWcE/8+pftgBTN57zHm51Iz
T27nGJq+meEMoGdlz3SwvyUHt6UWdMOpB5alv3k11e037gpnXM9YOBq0GW9OkQjNG6tnd7k2cx4G
rwt0OJhvEXKanPvGQsaRRBXTsB+AuAhYTEWInkgKhTOMtfY+3NkJsUWujxoTFFMB1QbeVRu5qmw9
uP24bEQRjwsyzeCYBqxXWJL4ylmlo7PvwfMhzR19HxyUaEhFLozvwStry92Gzm8/IXzsStuz+C2B
3mPb0fAouc7WcswtuVqiMdqajMe2bOLYP/Kp05H2yiGDYk3BE9POyZyUI7b6TAsxt0G0lwZB4j+R
ehXUGzjisEDHjlfk/V8/O79S6jNqM5vxwGLAExA4cg/4Y+NdOYSCgM+leKs9l3tTC5Vtv7Mc3JJg
ZF90XPfS8lXlekyBjvVrP4LDbns6g+/uAiUqMpRJ6NmPYQrsZ6oLN9Jbd0hAUydH9mOgp3hVRwn6
8ySruqRiRAPK+KliSSiQ3yAcd4uCYlj6Ytk1pM52d6I5kjo2Q6z0vFYTRzE4aO0GeT9zzeVLsW2k
an/YpTQm117937jpgPzn5pHRPS9Uk+f3aa6NqpXOBixoH1+BKN1PLvg6welsw7qPZYPprYWd0Lv0
Dt9DgBp1Ng8mWdfiEnUYXSc9tYbcX/S1L4zHtw+kgmVkErAdx9Yh9ncvIJyuPB0X1GSrx60Nqy4B
MHSn40o0DWoG8m+dITMWl5crrrTZxtg2nv00vTq/ZxLXCvs5MqzO6jmsocs4ligaYZvCNLRQvUVu
STF7Xm5LUd8H6g8Cepei51kPzsywGtZXdqZF7cn13z5/hjWAfpjtLQ5HDlT1EkXIHkO78h6S2rvS
8shU8keNYq9zLgyOm+2tOv64HHJVshBw++/AVTQ5OpaZov0J4UOCrdoUWiSn/xAoGXoPnyKckFZY
qi8+SGYyuJMcTp1FcFc2NfD9/L3BTAugzmKgxxbKIC3ImHwvyliztCCg6rkVXrJ6ogbgCKwUDloZ
kHcpvhwHWUJumEd6cPqZga4gyqgB++iv8sSzECvNXu7dZk87YIk7aXNKSfpm2TqcFldWF7qwv5Pm
xy38ouGkmdCvcSZsLEQQICG0IWjBGxsIkghF1KIIohCHFpDnY5GZ36uKec9qdsOGlstmh2E8QZHo
kDVFpeok5S+bdNYmYBKcnXVSxxjvz3aI5b8prQupCQACHCOhr/cmK35yLL90Bhpv/vNQhIPqGoB5
25tk8cdZDiF1umHyaNA+fKASAyVLF2lxKEoRZf5DHcRotdBDGthHy9XVBct79dRNw8bZnW4cevmE
GXgLfmL4GtakE/tIyFlpS4Ni0zGjD1Yix0fkcKWyzBRuTDvj1xf6ELo7vGRoThrqwVZpiaPBj3uU
GCbIaJ2D3C34hCbukVIhw751Al0r/My5yPfcIyNmgxQCk6fdaXTH2No9DrVjur1tr24QMLE4iI5c
HpKtKl/Gj/qfU8DZ7Cew2bBzlAGH2HkQ8yNCXdA5Vwj7k9NU0fo2u7XbQ2Ok+gSkQZJhi3ixzAuL
nxZ0iHm6KnDrARgewGsukF9fD3Pa0IqHLNV47bt05iS5p0xeAyP1xOeKaw2RUDUTGUfLwAxcB8Oj
7yUQO/lgRDTsA+22osei1MVERI8KFpW0/gC6826qEM9Qp6hwOrKTnn7HOYgtIPNCh+0K4xTrNfCF
QmDBBjYPZkp1GPpbYrGyy/QGTDBj4XjiOa4Cy80SA3Ea9SZygPF1ToR1xWpfqL2142qweUbxuWY7
LeyAkGgROy8Oj2/7qEFxLU38bizXj7COhRZWJ+94Nt6XU3eSPLRzLfMYb6jyeJVu1Imh6b/B48zj
gTcKCbJe9vW6Nqa35IpA8odeg/d8uQdMBw4DYFU5aVu87AwpP20ohMrHIdZeyGPb2E42YaApa9yd
Pqd1eAMdTNmRaQp/ikjVJpNpwHN+lv18FFlmDQBQiDYDB8HrCtkEASeVVUUBkWJdAeEOfGtRv45d
o2EisoaW9ZzYi3b2fnzX35HD9WCGOOTBk8Z5c1Z0/pbya8RqwBPNZm8ybXmzHkz+QJv0WxytQAOm
eKdHQghodJS/v22nx1RIpbOhMma0a/5L0M7UbIKOTriJABgFffltJh4bn2pjzYuRTe6kjqioNFkS
0iXhQgO6H2GS/xzgGWPsZ+MWd2XOw/skBcI4OAs341NNvohlX2vEBaDJILU7XFzi4cBKm2wC812R
x/OiLt/CzK20ISHht/fQDZKMuKxndn/CQ47neAA7b0SNAdyUE8Q8vXYfzMAjRJDOEaDQmVEELPjk
aj2xPh2LPnSPIJZh2V+Au45FJj/oXHJAo8adGHs+77QV//6c3GnVrBSohuVe2bSFAF4NTIns7FqX
syT057/InFEUDNWXxIz7srAuTI5tcnbJ/mAX5rAOJGkMHtdBRqE755DEvgV2HoSqAfbbKvWDFHvf
WXIWiU951omJFnbsutHIQTWc/oYvVYcyB9wlmElWFmqp+1mcoNSTeXg31XHbm/mDK+b2gmtPT68p
wkzVG6N6X/gZ31v+LHS78ockXt2vWhK3IW0ebuLCinyzolVMLdkLI6m6/qyFtQ126LAhlNs5GKYg
INvRtbwdVZRDokNFRGb05qMlxkL8cV1wlqYJj9Z1UFuX73Zcjxe+hIlwiecFMCJxVBeeSHTjkdr5
JDA45a4N4XO5jVesfoOUSFqzuXExl0KhCuByzcl3YU2SU7DjtqjnanG8ChoVPEVaqTL7Iq3cpcqR
6wk+neoJ+i7O1b2bjqYivN3lHYzmTuoFOzHDP6sgixJukTms7R1UAQNvktRQDwqS7jtCIa+qp/TE
6AckE7w2Pu8w4sEPTz5cmi6nVBPhjzL2wQOCdfLju+bZbnny9t5nSj9JP+VAIKVm9bTVlSrDRktA
LW6feFe7KSBzlAEMlDWsHCq/u1sGZCuK17lSVeVGkPM87crobb2PZn9r3SI6Zm1CFqIINZLzHK32
sh0nN0F5UyZeQh9DVCHwfb1UoaYxZRtyVpYKdfKrh7anWMRcHe61IwkWezxS0wtu+A50TS1cxbUU
FY6FPVMjMHCemV8SkwwkWQZDvYdW/c+vsW8vYZnSlhydqPmN0Nodt42Tvu7B8G58DxFxYbl8grro
/dHgPdUrtbW0ERsjTE8ua1KPDiPwA5LDkJea8E2t8yZQo3fVhM7fc9TghEUPFnXg2ewr5jUU9Wh6
EVXCeynEarBKbE3UrTeE/Wp+UiTBYKD4ZqrJkgNPNSLeMoJr3Rb1VB59JgHbjBhZygP9ZEjnzxfz
FXCLruxGkQ9zqtMxAFJW2LPRgQ+vErpx3rBxR1jbkhr6bu7WLwWL0CQ3hgA/HJKd9nEaoHVmwvTg
Ctj+awWi8/otpCAlueDTzpciGbCQ5DckaaFQV5x1YUYfQshoOaOPD5ydpystnEAcxgXoP0SHH9PR
6Or4vSnEfjKeOxM+tmR/esJftFZakAlCA8g3zlEBIKKP8igzyC/Scj6kJUNVbeV0bSB44I6U6q0r
+LZ1T4Y18MAnWLuHxVu2OBf4B1Z25kH16tpL0YflakzPnbAd5AE/CfMyEWWb510eU/QGbnwxLZEm
/xmaTsBlQwzs6Zm2fMjtcljGln6E7Bp2NfIrNRmdVsz1+EvUhvKqPd38oeSE35T7C7TLXcV/WvXk
Azp+gYnLAI5KA2RN7hRpW9Ev+suYBsk3AYa87VtIa9nedvnCQVsNCPB/BbSF+3BR8RIi+HFqTbWn
6a916T+5i3mB96oBTUki93HE/wbbj4X6TJ45J34GfBEOkUrDqfZ7pcMd3Wt9HMOpD1EjRw/2oudW
sIBLpL9seWGiHUIG9lUcsN+a1PRHMWHt886t4QdPvjNvdftqdbrtyXFvwQ5DUG62r+3muNZlLor/
hs5O84G0imrabtFHw2uLqc/1e98bJfiduVSblbP1IYMTdZLBNonC8JiOyvkiRIhmfWkeZDNd/Lba
Pvkgdv/x1lBzNEiKR6ZfrdiPUGtqagrMSAxn5sPj/ownGtnUJY7bPkmxE+GSymYcyEtQJgpfH5Fl
WqTI4QtAvJ93Yg5MNNy7YShSF2CXzwFTsmqqQWkf80HHbKhOKT90sICVGWbL/fsgYFW+HL7Ibtyg
a27PKp2n52W8q6tUGx6aQbefVuF7S9QkyYjnkeVj3s6iCqRWvVL2bYobUw0zqbRatRIqaz5DjOlP
5yo2gqxYoP0W5YF9MrwnQCquX/tS7IOezXsokE5DVZ5D0g1B7miV2TeGZIoVseR/HGLA6XvyxPJl
NJFLAR9Im+Ty5b21xp890H66mlnAIqBUPwNFp2alDr+0c8Bt+lkVTLs8UGWOWqpMknKS4VxebT3Q
mUtx7avj3HEfc0WILZe4jRujb66rhs1jLiHd+ZGQqdXFuSMRbZggFPf1hvZZuAUKTSuIKh86XZbX
8u+UTnDxeUD4euMqjtmZGfXaEuiP3Nluo/Z+7maBiwsydHg940w33ahkYbPqYMdSt4rvFivWDo0X
nW8A+vZh+pr+3SH0bCqKMjj+L5dCdvJxeG71lhcViVwFuhN9e5lfLaCGhOev5xHVZbnPienyot+j
UBNTAaN4ZL6z5YismCqhN5Aeyw8FHCd1skP1xXQSouG8QU7vZdSC7e2PlErx3fAOUli9fEISADGD
K5nQqw7oRdvYTewTGx2Dkko/S5x7atemt+Ekg4PvmFV1rsUo1xZk8LeMmGL7lVatTV+DelssMMt1
0t4avsYYJx5IU7a5GciITxxAnfWHRN/L7F/valgUUCB0+KpdLW3Zpf9jBTfnp26Bj/AO8a9l8aLi
GF+kGRw7DUCAQPBf6ETDm9oi4bh3HUP7xBBg+LFllb48Xs82c3JU63+XhBKdSRbvAkpTAPS0vBm3
+ql6FlpkT3EBW3xVZoxNamEqRGoRjHolwEchl4ZMpSFk0XTEO1W2fVLoZoFnGTJPFlYHLhlNZ+m0
Sg+/1OpPeYNs1yalB3+XW7qO5pAbRfw1zw2bdZYZ4NnY3VvxsKQNFuAjb5Hw/KrXNyhdpkytwaPD
8A5J3QKf3hlyWevCEObvbVSZrN0XV6nrMoiN4gif5K1uNe7Z4alOmFlM349FS9gyLxdMQLHQz45N
4KD2eubI54hki+TM2fWiFxiQePynqj8HEKi0o5a4V/vv4b6Ofs8wUaeCsuCaUG9X0qjUIUDsYIIN
GvE+I+eZfKhLRzeIrTbJI9zNuyY05yleYVNvyBsgpOcP3sMNy/aIImkAUVq4gks2VSsJznfn3vLa
vBbqqYBfZEcvnR+cvMjIYQRaSko/fFr4rHB4WFBPUlx89c+DDEVHBkHeYbEqz6OvP4oiOjLjstgd
BNxbkU0gB80BiIKBdg9/yl2j8aDP2wX4s1qEu5PzNhdlhWHxVXTz4W90cZkm5deko+iC+cRoMe+2
s2HA5MuzioVcJPUo8OTEYEzh9+ucr+ninL7zDcRivpSF7Ph+ZkFPj1cOIOtLp8aonoJJ2Iy5102r
1jeFt2pGh2m/O8BAfH9GOUP/4V56wqCEMhfCASR+rdXiPTOooVQX94WT4Uesa6UtEtvW7/llU7HQ
HUWzgbhAnFX2m1OCJEBmobKDUlwEhdufZ+hq9r05y/KiWk9oj3fVCdL+pChyJ32KbxTc9dFzWis7
O2R1wJ7WpW7+hrOA8dXLnSATOxpAmXkIVE6CSJG/pXgwFW7ro49ERxsc+jijmtpDfT1XbI2G0Im9
ye/Z45ghQdvgP7PcyPtQAs/92Uk+yCLMI1YXjV+nNCugEw2C1tdgnfptEC1vGOSH8R6hH5ryxzxH
9IgeCX//8IENv07y+cQhG6qh9mZWfq4/9aZmiQURYzVUjoiE/F6acPAHvifKJPGscuGSYconLyqe
HE05Uyff4rKy/fCoSYXinkpQhMjUzUWO3DIM+vpQ0IpKte0sRTawYSH0wEjAF0cGb/iCCYdY0oPG
5/qYu0MJi64f/18kBK2Aon4XRLocFM2uadHSkqY2LTQ6kyluyVgWSE+zF8re5b5qdCEQ2CeknmQN
rB99xfx1zYVRD4EVUG+QYibQ+dxdDCPWo8lz2deL65KiNO12tUMHjfKlajlXY6k/337RTw0w+cSW
rFnw4WVbLS15OoLsiRtV4cYUjYuUnWgPjdkzY3ryENOMjEbCBqOQcUt+ZjNR0bg1m12xADsJ6s6b
ggzNozg59T22ZkOZ1vz5YsVMeD1jV7J772YPoNCIE2CK8lm2v3X6Pw+eh+4JimFcawRwnDXNPFJ0
L+Z92Us6ABJbG2GjRl3kQ/JNW0YOy744FHjudRtYUao0XIb3mzg7vcy1+LD+gKiGANZjKf1hyS8u
gVOcQjZ7P7jCT9GXBVeijS0H3Puuta/9u/Evlx0IWEwpVi9Jx1qqJcxBV4j2Qg+yTCSwTX7Z/Evn
lMYwVISHXmWIRFS5G0H1htXZ071A3+hPh5zAOz+4A2zo/781lCX0BeKO1pX8UYJ6z1Yf72t5+NkL
Ap7aQ34XIkCa/i8inWTi42Mm3OzPghkVN3C6bd1/iilw4RuC9UhjtLlRjs6vt07a53wmOVx03o5k
YeK4ueDRO9Kr8MZX5iA/yo4Iqd8pLhotV1D8gDqm6ircBCQywk7YpJmu9J7HZB9uKbcrm1zL4Aib
i2k9WbK84auzncPU4arL1vWzXCG7NQdAsvGwrjkF57tzLbcZgNl90phmDgJrOzqryg/PE2rHTWRk
CvYa7yFZd1kA1Gm43TCem6m2oek1wpF6VQpeiM6dTYLVhrnVmqbzvW3peun1dCkRsD2cno8Hb2mI
VAb/zFHLrsbrpXBA5gXXsPLV/FiUprvk4j7SE0DQAQzH7vrK2qzpu2rzEKKNV2jeEoDj05aEkYqi
HkWaKWe5EvdDDNe8Lcr5sr/VncCJkn2b5o2xelQMaAJjjMisiQYKfBXm+biEARkGGvCYM2YcjfiI
vIULGEB6IrRxK98YtnS5LrCMn/mxeeNK4rlcIdnbXHI+ciyLqIc2ky7/o/5g2cSvUte76OWz7nAe
KwDo21WZCbFrH8Krut3A4p3V7w3IdEVsX6Kp/t7mHAAFab18pkUZdr4F0zaJUogMo9hJVu9zLYaT
FUpTEQ9f5MeMQm5YiJwb7jUMLHDpYrdQdoW7jq87g8+aBttkph4a/fJwRTLqcqCiGREEbNSJ3nO6
77k/57ph9g4GhHd+hxICZKlOJMo1vm853HzN44zD6PwmrXBnDR2Lzk89mIa+Zem1OMb6Qq03lvgk
oS1t8OfN8W/kw/d8b/SCtAd+AZ3aI48yNAqRIwWOdagXzb6/hiMSeiVRrKnMbjXoVqViynNTO1sK
SkCOdjjPBVps9kRJq0+I/mVruiQKPJzkdAZYZU+9b8nlnk57d73caiKjCN4zMyO7rI3vdVi2Cq3V
dM2TfZI21lM2ypQMGMqO49v8eJgG1vpNtaXRxNA8EqXBK0dQY5XTTr8CCQhmhiD9tQfOaeo4rlHx
IkyRiDxp7oMTBFsDRz+RKlwSgP8+C91lFerzE+MUTXNhyr3dzxldhBpOIOcl0WCUev62EFWDDePB
8mJsCKh1irRcGNx6NSDuo0ugWIjmjrhlHBqjjn2KdvM8+3xddcggGzHqWU0s7Cprs06N2XHQz0Rh
13ifUWP2Sw9IOlEtU6QkGtEGinK9c6944MvDAgOy/tD/we+upFZ1tfBwKT+Dv7PYDB8Ubc9Ij98/
e2x3hQLsZ7BXUsL4WmoujF/BuTQTIgZWl8yXIq1lIFsJMm78zkWxL3g8zVKAqbaqpMfuaQ/hvNjw
BaYwvmCIXidpF/uhgYn4EybNSvJHq6uiKWG6p0a9fpCmOkLBbgpaApp7vRmPzR7g9+2nbqa0jQ/c
k2pxwJ4Q9sezr5kKMgHylc7VFOSOwdw/Sd68Oxg6rKCJwkz1EAo2I1986XNAeOi8B79OVTz4t3k6
CetvU9DIZ6R2SBkhI8Acg2SvX2hNbJbIRo4iUXF/BGraeeJSqJaj7oU9vbobSLpT94oZYLOer7vu
hexiO9h11kialbw+7nUXl7aw8D08qfEO5Mm6QP5kUHaWbm5miwJ7X8/tmHZrkoVzcR1IObAgixGK
wciorOL0MzDLNS23n9Lxw1GtCqgG+xIpBsK4mmdYGmhMwXep6gumw0fy+5TBApaTLUgOeW4cEMsp
evD60kaRrgcwQXeYigN578Nczq4/KN9s57L4s17Ly4aiL/HGo14lwkrUHQABh5AvJhGKe2W97WhX
euoncSuP++Hsht9K4Fm+f2ZCe8b6RGe+jax8IYRgrwAtJpdwGD7uOGYSSkyRmVnea7+ICEB2KrKD
XHAXDufET8CuA+MOQKUM337VABwfFbZwm/EiIcNEYbN2LTMtlu8tAMjUV05eV15K3ty+vaPB/QG9
rPBVEsYfeoRxD5UPsywhMXGumW7gWEm+an0CpLzw4iUAtGiuJAZGzHz7ej+amnew4cktIywETfZP
J3Uyapt02wWP5k1z/VDmF6diD1ggkaaS1Y/e6dMMv7iglXRwtTYTwqw3nIiiXYX/5FRGA3t2Ba4Z
9JqAquUY/D3yXjaArfKEq5jOfgPV2fcPrnNfIY7jl/M6LNrYuD1CXkC0ijYeHkW2PUPkAjZt7xxF
UP6oIBjZKc+Dw1dfxw9W4NBiEbTpuaeXjRV7hL/25gTrZ6taboDADsYwSNONnxMRi5B4IqzoZgv4
eFIkMR65Yx/ZcGrhWeFojUme6hBM5J8/CfyN4xNm2o2ubT5BDGeYMY46Gg3HSv1NGtznNEtg+uHV
5fKlv0FUsDl3duO0sTZFpxZ7FM7JF3tJ9S43CrfQ8pjFJasb4r7cMIyfykzioynqvr9h70OveYsP
GSqNaistMKTAFa0QWLCGXmJi0CHE1wJjIRs3tpWb3PFnM6G9r15CpFwsICv42iAqC/gKRqdoa1dl
CfrAY3nMcCjK6tmIKjlb9xTpkqyhrBRrdbph4sAFwIDkEhl7GfvYPIPi6lvKisX53n57wN6McXy3
ARY3fVVfmtWpypGt7kg8JjQebvRBO2YZLtPBx9xQuv9KVG6zJ2m+RpKQZZjjT9ashU9iB6LdreTX
mdEjRoAEbOFR4JQYbgw5+OvrvIkGphxzmjE8DnhxsqIrPz9t34L0jtRI7teD3g1nwKpGPbMLjc87
AIN+bOMUmqhcbq6bsZNcwl99LenjBBZtA5wUBpcCfRCnXcnH12G0rMW5s3ze5tBD4h1H5syPexw7
JrSXAETSjf8QQ0dPyW82MgtA7w3fPGmNKf/uaAeShi+Ks6a6LogATX+eet/cnrG8JQAKgo6E8XwA
aFSttzBp9Sc3jI5JS6fae3D1wR8/+rwrMEiBlND3JWwOf7V1x/d30LJECu0/2Hpr3XHsH4v9NZHz
HmjnRPwZm9X+D1omzvSg+sfC9upQd8d08eFXFuZyZ8+BLr8eKifK7ldTucUx9/dR1ycTfTGzMN24
vvQMQKfz8G3FmW8aH1OsqXB7ARQtFuPWHPBEzyW8NLENPtYzOnz2tq1gMJJqL7dLJD0CnTHI31lC
PYDOb3sEMSd2bffjzoFv+YO2loOY605wlfewx9rB1kaGFhglPCZaBtGwePgsXBJTawQWscjMcnSQ
03daFhID5LSFXIWlvGPMbonE8hXgLHX00YiGWtNOheOL1PMQf1fLlZE6uaDTJJ8FC6Qk5LA1R9D7
YWQqoKTj6lsx+GgKRyGrVqupQ5PxKqEbIFFvbI8T+1o5N28P4xmFzDyB9TPPCTrg5QWQh2/SLD2q
HDi4+goJCbo7vp/d71R11hxKYJnVc5Uch+fPy0+zEoyTnxtNEJyiOqn4wMxhVhtt4ebKK6zTZrn0
+Ev1EZi36KniykZ3P3Zur/tScNddWh3jPMo0e2IjFNOVuPmuGV8fAMwki2nebmPF5itGnCW+baNC
d/YgeNETB6zSobQk5xlDttHSzpR9lGWV+FBIH0+za/MDIYtSK1h7joiQvTb0dbNZIbDQj2FJD3CZ
3hFAgb4/WGkOAffj28XNqmf6RDhlU5BPiH0TV9x1dgnaroMYhoA4aHjC5oEqBASeoV1vb08VbT2k
6USyQd4l1nxylqLQmolycUxYhnZjm03njEuSUFRKENnd6ZDH8uRGQHpq31kLC9EgLL7BB81NztjC
beJ3rM5ACiPFPfoxV9AesWhCKy/FeeRzVEvS+fsJQQjTxgFJpAeXr0sWvtVWWsEfu9hs6owHabSK
cVH9KeZhxmkzYTLG4/qx2sbvHXt8+8+RjQM8tA3KW+dbRpsE0pWckI21KLqdZ6f7eUUn3uqVmbhT
c4FitVH2E5gvhtDkrRaNAtPpBgUd/OupocQ7Vyq1ZbBqocR8ujZOKZeIUcGbHiTjFfprcY9KLcm8
M736WmOsuaFnEaJdA80LN2YsbkkitjMllWYd20wksN3EKW3lnh8P15mlLXP7HnGcIbAq7dWClEXg
cHPjOVa1XIn6771tPo3OYiNwalnxO0RoErTH9rw29Z5AExa2t8qy2dEokZAbgdu1tKxDR971EdRe
Z0Ozpz7u+AX6wR/9+NJigccNLyb3IudyL56TurZuOJyArudLp5A8EuyPcisJOWRwBxmXUHhkLkmn
voGunW0Of+d20rsxBqr2ilH5Aby82ej3na/k6tpbqPSsbjd3OuMZ7ylBsxD3DzaAC0H/VWKTTxgc
T7OUfOKQzg0Et2JGX3uDkdBMV2qAV/3WnlRGauqPIpUBht7JsScRLLEpgsAny0Sp+fppSWYCEBsj
qJ1J1wCa7QBF/a63kSuoapEeH5SubvnzNNY6L+2J6lZGQmTXNHwbcUG+UnOMv9FSXv/5Fod8Tf9V
K/IJLipMzX6yVVeIoQOcg6aNpSS6eXe4tLE4JyFPYPOexwUp0XqQUXW8uRecqeHReaxECb7iJkUv
2YgTpk3uoNwvaEaQiajvzxRWiX1pX1ony9QNUceKnnWvwviR/uDN3lHEl0i1vcZ9mkbtp7k+6CD0
u2aHF1IEnyXlHIe3i3k10SKZiVtvQOUXfVPuTwVzRYTyteexqJaXsbWjFgSqh1cdl6UjfpLLrALX
M39X9fytZ/0gnu1360pCYZmjsz0VtxhsGmm/CHMXsHHmynOWWAUxoGF5NfDWYMrs7dF9DScHAwQK
BJUGH6+EeVIMmja4pmR7hQ8AIR3EsbHvBMf+Y6mT6NC03S91/VePMZKqti2bf/juE0YB+MzM/pZz
GEzOARPBWBS1BuWyK9qx1XB+mligtqs4NL/R7GI3Ax+3lECRHrEtQ9ZzNzmyC5ug/JNmetORm4Qk
NnuPTB8x/jH7mpge2YzjICCluApfHI4g2pVlzniXnB+AaEW6X9r6yYFl7WVQ9X2hZzXpjY6R0HLr
686qiL+sADY6dRUc21/Owafy9nPkTzZea9uhKrbadetZ4ALWHqI7Ohja1SwAWt8gOc+3f/s6+n3O
0UfkT/r9vy0cETbX261VOMOCitgoUQRfXtqcCOQF+drmGfPNht/Uqggl2FAEcWUU8B/72kbgmYPb
tDQWcprnNOxP11LhtAcLu3mPPIRu1NJQEqxfiaqKcsLmfk7zaZsLkQ+EzBnQM+ZkGOB1pSHJjeFg
XuToTc/V1mvGVqNZTBRKnIZUbpZmRma1sHXc6CuqbSrfSFqkwvFqCefifNWVxfx6eAky54hTKQFw
N7r8510INf/fhnjsB7092R3URURkQg5Ysg6HFF2eqfaR1ktOo5K7oooSR511sW84Lwj6zGozrpld
B8YSpIBfmM2k/A9vh2tATs5hW68vtZ4sCjAjNJSC3nSH7RvnEVJCWSmrSxzGXo/7R4paQMMf3hrH
IRNF5WrjP8tI+WTCniFMUebWMR2hQ2CuDzjudkdxKH/F7O+PlxuVChTWD1tv9XyEyLza66pMI0fM
z1WUcZzdoJnju/LA02yVoh5QsOsONNIDIvGUmKzAO9idlmScCWcJmjIz5/JZY8gi9biWoxQ2aoGH
+V3t4gerkZCHX2qfSen5Mu9CzwZAoumqXlTMcqSDYqTJ/FW3ApQvusLIeXRcPOupdBSmG7AUk4X6
WFinQgB59lSuVL0HO5ECFv5PJlrw74CLcPto0DDaIzbmK9vLaD+V2f2f1Slrx3ZnClNhoD2EdOUC
ahuy/9VJMiGovfz+J4cEg9iSazlA6xcz+FRe7sVxW8nM1VN0rApQcYtxNSNnfAL7/5E7eHUjeM+p
r2kb4uI1/VywWYf0C1Zg9zu7iqWQLUWpwh/ekgslRVrmVOMceVVLeANjP61hpT9LS0dIaCLdOw7I
Ip4fHgKuW0s65UlGsga6DoDFPoYsjAO1+toeQlXdvr4+9haxqgVuFd/i5Rhz1RHovJP8Mh3H+rVQ
MYX/qWU1oy69EbLGk3GkDM3mCmrio2g7try6u3WXO/83kuU/XvanwfHob2zH9FgqQ+VrIsjad0Ei
v+3da/dhAAjYzY0g0tuGrR8YNpGdAayp9SqdOV4dkj1e/krK9JNCrJPW0d4Ud9h+YVTf6ZPZdRWj
ocTN21DcLTyCo1dX7+ejUM3g1mpHMLb1VoPNmjIhU2zqj7FkucjkXvqECnj39Moliciv/RVxpXdp
FWzIElObK0VOwVyifzfQ/A0aHM9JNgmYiJTgDOcY45F0bgRcFNikBNwpDU83wu21j3inpIgpNzSA
jvPttK0e2mZnbNRgVHjfIfx2umh3p/v88KPpQ/SQuxfVZkS7cVpZewe6eWQ5gZ39f/2nSVs0lAxw
g9mprQVHUlseokoWcTTkbiEodDvxRyEZJMiuHSBrnwURyYtR1QD4czJpXIYudKw8MwCYGkPzSbwP
hKshZGwG00N69Fsj94K7qJ0yq75BrKwL1c9sdtBVN2Y/d6o1ZiPLACNNL9+dHVIqsSuHSZzmCR1y
vxubingigPXO4Q5BeOslhIow8SiWbBM5L2HnfWcxlV4ih5WZJEbNuPBnqXE0Wf9Mk/qZg/SrX2Q2
6Y52XFNdIBAioTU0OaDH/2ShpA/oT6WG+IIlvunmmZN1p0z4+OYL7F+rFYxh+9aYI48hJ/CxTTzx
U3Qk29IgA5FdxPD8ysiL1YnlqWeBd+NyEB3qnx6iQVPOlloUxzTFsbeyglGHM95FGGyzuHgNW4J4
zhKCwv/zLMmmk8ofAgGHSvYcxB+V0wFrsjXrFNxg+VRfFEsx+NaStPfSkGKXiXuDvLmxtDagMCPr
nQo3JWxM6yva4kA+4soA++blGp5mehe43JtFn7qQF59XLVYDf6og3Wa62444xrJ3lpDxF8zLVGTr
1iygo+m/47X2Sbt5xq1c0lqSXkQmQS+dfouOmrTRkcRcXYC23oUFhJ1uq2R4+8jHkb05eSZt0N70
Bjojo0BxKLq8IHSYIH1cEiIhCEC9MfapCUDbJn9SuN7R9s36bMFyRUDU9uloEppzaqf1ap2OTkEU
x5y4HrdPoRDZqfrGxBF+bPmt0pOV8/uWlHgrh9wUWUK1MdjOdyshohtolU3OQZKGrC3/FvHkvHUm
79RJ1jVVCk0a9gPnNvX9wSyGWnRwLlP/ruMEOCBkNfK8wzXpjxCGG98PwEizbHbjou2XVAn/NPrf
CziFKkeGxY/EGPDvA8vpL61j+x+oAxJicf1wUQujMiu8WqLmVT+KsDwWGSINhfPyHbR2zfgLKZeO
SP3+Mg1hMXIim/ARvhMUKEsxbxwG5toEZlUbQbkdluGEB0gN7IVO8V5ylGQgHyJ2ELQTXusiL6iV
r8ytsLudvFuFLklOewNi8E6Xnr65V0Zsa2N4beFmlHh4CnalvwQWOa1hxveCfzc7TLimGpPYze2z
mNYdd2rFHNKsQJQKwQVw/dYaQVnHH9cWe33HLZMFKVJkodeWPHMLaVH1TAV2CLpzfRcEC+koO1ue
/MD0//AoeGnZDtAZle1hn+FU0W9EaFWhEz6wgJmif/oSkmzePJHA/C+4zxQKgq2KLyBdhWzdix9W
m8SpwzptGehJG24XBDaWhPLYPX1CTiyiDOUQV7gOSIaWHU0EOOItpg2mfO8k28GXE33lMBOT3XKW
UTiuib9QhtnPHVJ3nIGIaD6rXIotQjEihn6ECIyejxyQZP+I1+CBg2951Cm4kxpqn1cnyqjngiWX
OOyn7NDndvMq3QjlL/b+sO/IwQkLgyTUM2i/UA10LcM+aNhNB3MIMfHGye9EfoCAD9jFNcRugTpQ
GTFmBSC0c6GLjG9UI9zyoKRz27ym6awPm8DqFfZZTX9A4sHunJcRsFZl8AEAO9anqnz9P6Q6SxxG
dggVRc8uLzpfxxLVUslWM4hcp7UAg62q2pHDqAmVdT3XNb59dBvk9hiXN84RzfOodC/Mx4IpZ5zo
D+gSt7g+VVDEaHlpf+jwPGND0kvVKbP0Djr5He31AFc+l5bt0r0o5ZWxTfjOI2yA7tn8PYdET+XY
RA7J2om6znevOaLqVJlCbbfgd7RSRJrdQd1B75NOgQMoSw4C718FCIjKFLja5v6zgOTGD2U/7z4I
KmoCzK8BDynVxzfiblDOga9b0MFKI0CnjZC0hQjoTaa/l1nKAoCgIsrQYY8YJ6zzcQpmjn7LhDb4
h+Lny110mLpmgdcV3dv5FiBPEfWkoqs6GRiLXeCkJDG7eyBIjNJ6X/rrXIy11Co0bpkXXo/DW+lL
rar34PgI2kPH+5f5zN85OJJxvLv0RnUgHfIURC6mzA9ZN5elVRPyP5+9BNkVMYsuL0RodnDfqvOV
wupmfJkzgG8CwFQmd6d9jSpbKzXjNNQgWUIDCxbMgKJBUSm0buHWyHt5MxXgdCST1GeiZNHjssr6
60PiGG6Ias1QxOCSO7VsYdx3GqXhUORLjL7w2Mrqp28KJeXaJBbYwe7kDeoT3NYUzfUW1EFdtXjh
fZK5xsWPR4eq7WeyRoV+vAnbFa1m4RV93PNDNDmCeJ0B4fBZF1w9ASZqU7zc4Ejz1Mw3hDIH0dqr
iCv4I9Xsf9ay+9cHztZHZM0SseJEpjpxRtq0GZCYynhovHuj2Cx1ElfDROSTFN3yNqGbMK377txx
Hr+4wMvvgzv2z8RJdDAGW3qT7fZJ5cmDc0ChGbfv1PersQ6Cb4EJg09aRV3iCPsC4EM0p3q6zQQl
ZGml1WqQuH4w8iWEOhDGNpY6fARP6rY6Hm54a+sbbsf9D2oWhZvl2oJMniwIs7gEtOCBhgbsr1Z0
ucW1OGWNX1E/l9UW5EPopGkHJCnqTUZhLudV7joai+PK34jNl6MbhCgqi0LH+6pvoZA7IA9027w6
dbqbjTf0GyrKRWo68HmdTJ6FvXSHx4JlHB//iZ10IaHU5ucnHhfdVkDrpc4DwmFkyZ3Atvq7v2Nu
cGsPFqtRHKXuIqUZ2xfc9LvuC08ssevME8te9J5ZM1uCPtvhgLuHNRtnk/40CYjqD+djMlvFjGn7
l9XQ4UsgSjBPZoCKDqC+ItF9VoXPaPzvZhjoLfcVmZk6ml5crcLWVMNG52oeBz15vrrpP5ieGwES
5jBRC/n2AhQItfUAFNAS2kEexOD/4wuaxcsOBeGVh/cBadCNDqudABNgoRAb28bZ+EJ52OW2S7ra
mWwNnXAd8PuOpJBLf01Nrkq8lQ+0U4ITEOAchb1vGUcmAJkgLxdF04K4to6x3gZbcIdx2Z9DWQtD
3MBTm2oDXXXk9n45J/pFhi7N2eQZ9Y6R8bn67rwewLxSChbmBh6cLQvEn3X0UB8hzF0YoJEOGWJR
KhLq94vms55f+PXIv7MQO8DPb/v2cp7LKYzNvf4EfNLar4namRl243Mu81RalIhwIo9GcsfdZlkM
5hZrFXfm6BaAAhAGWqyW4HtJASWtk7uy3kONmIDkeMP92fuHt+A0aBR9kvcTc40Nl+kHruFTyz2l
TmZCUq+0pR4maJcBH+7Ojn4mHHQN8T7JT1wxI5ciPNA4itohoaL2Lr98MkgdaxsrVCuSuKM5qAhU
vdopaplMNMWOi/+bI+x6fE5Y65Jf6Zk54HIgg1YruApX05CQRsrz5qPJsP2wsrELNwPuSugt5TH+
Ozb0TqevAfFLdYi99g+Jub3Vdq4zzwGDUjYZkf1YTy9FBc8SC5z1n6DsI6N1EgdCswrxrml7sSLo
2wOErePAhf5NJ6oEmwcmI+mOM1CD7j+fmEP2gsynm0xzLpclf5u8OzVMZWYNdy5G1NWiIvcfZ7Ld
5G9Na0YUGa+Y+jtlIvuIiylnFcwOTbZ9LwD5RVOefQEb8wriE21eqXaeQAg+QxPlLvJZW6QGOSPL
WOuMd+/d8AKyn1Sc57+YDJues18VTTaczuzDtyTK+Zb6ddVqJQXc0FIwsKq0pAKiY5nlwbf0zZ0h
jvn3PNoO01o175SbLRcASCe67vXcLJrhwy6Ulh4YgE8rYKhltmq5fAhVx903wyIcM+nDcj4EqKc/
IuE09Fnid+aDVTjCbNQc0/a2woRVO2H0gNsmuy5qBccjxUV3M9aGaD00KP/BjYCGYjsvuxpO8gjM
/Vj8NEcczkTqpvgxJ8/paMc5+ODoGGryniPz2EMKE59KA9377AoU1uNyKi13DO+z2Yys/mTvWWVO
GU11kK64ab+g67gxB3mHRiHLlFfMZCUurD1b3yObRILzGoXJgugs7gUGykTFwHZZlFqngMuaPSs5
pYSJXEIgDES3XMhea/isZHjw2ps0N6ZUHTKlSmxgoZXMtTQLRAJ55bszEzYBVjLwdJTE9lLUQZDv
yM/Vo2XmXQ5f3vZO450oenouiGNj2ab4TKYpxTPpPd+gA3TqhL6bd/WEAVT9KZEP/4/xa9gdQq9+
/OwdDSl1KxV1ZPFEI7bs8RoxGr/IxRJDecf7oX42W0iUd+AH7WLahaTFbfdpyQ+Z7EV8PQqK+fBI
lKGWPG0b72/o9gMY3c7pQKkZ73vq33cjdMoWo1Bk2GR6xhrjyrdRiqVjSgEoxz49oieqUWMXsTqM
OhJITXyth3MSpvbo/CEplW6fMlfMtSvE4LGeKciWWh/iCiRN9/OEiXZD5XPM729dveO2d60tAh2q
gFqheULjo94bCw4rgCV5XfHhv8GOYoeEtUorQE7PgkY6tGGK3yWbDb6iNuhhQApMX9ckcHhDzrCW
jIlAdv4JUXP4HiHEkwCiRTar7bwMahZ9tjksMbYbPCpX/FWTZ3j+mCoKisWm1hv8WLpORzI/yaB7
hm6Oi8tptf42AqlWDs2xlI6e39xTH1TvggoNJsu6b0MC0bUKuiBvn6fpfU8vivXIEPJwQqQHb2jf
eAqzhYoF/meZqVE8ZbBlbRPP4CbtX/wRo8KHkOpKa56ZIIJGnEOR+UWqpE8pyigsdAP3MCrzUwyY
XeeMYEvN/ujbBaHqqxtCMMp2KvpjqGbLQDlaiHDcPYfwyIcAdHsHRFxh1maCYCgy5DOPkfq5tp1L
l7WtGRkQPVK0FtsleDawRMeSfAo8f0LlwsD02UfYcSqyPdk31AG/GwGBogFg9YhLYdfKN/w/16S6
G269bVMDUZJ4m1RLLDxirJG97464qn63to4YjgjJiQEtMDHSTpZ+uLUJbcrx27GUOFOQmZbGn19c
fYfbsOuz9MUHMIfBKPWaC5xEfDp1eYhZCqSG+gfrhmJiQGradVz+nGfjx7BnWgxPBMHYEFsrRP1l
X+UGl9gprp4XpOSe0M7Q/YXBWSe3EKx1aFQeuCvRymZNvur5XjkpkFoeLoofUSsgn8/KrGAiT3Vz
ugAUlAu8EbSMGsCCRUsmcSluSETL1w9bM4iDLlUyZRS+POUhapgRODFRPJkVsAcHo++NtYUgZVKm
LdZv6Nf5npE2kAIFKaAMXgS5pPHFiODKLkU6tzvQkLoQjtnyl5siw+M8L8vv36wzmrjDLkU5BDvl
072Xx+dZI5jo1gjdM/sqiu+aJjOeNSHYZW0cQ99Cz/zoWLiDkOI5cJ13Y2knaMsrjTQ732+7YTlk
5DRvBy3og1kqBZEjM40gm7QY/7vpP1aMRaMrNr0FVu7k+tIPAIgM0CReliZoawtiO5UAHGI+ONCI
ANV2kl3juNpSlnRnq7ay6+9FXIkB9NbEmE8iDPMb/QoX7i5JLjlqEqyXX+slW3bvI+KW1ShNvutp
Z96nrlOxpNmZDjMlIdSKQYq9NQjsW1xpasRPcfbsTE9m6zcZuO2UsptSRaEnIsjSo5wZpytVZ5Cb
hgtoladZSQkio3+lLe0Boo18jI3ie5z5hwTGR6SHMdhda4JWnE9nZVBZCV+sD7vR9U35fUbvNneZ
mOvJ1qLUMIfJoDNI2LZque7z5gF8RevPq3Q1NcSxZwaYIseXGbXZiBGxsLgMBL4cDtBBrxrcGEQ/
O/3f3SFFEONhVi1V+YF0abmmjnCEX16gZPTRfJf/Fa18UMqG/i10y4wBqtykdEz46e10RQBQosus
eCAdYReRSkAsAvnehcJr/ROM6reDdHt9k9m7ke7cusTo0NBLNO1k5tRNHH5hcY/XCL3BS8kwxpl9
sgAo1zqB/dt+cOaZPElU9ytLQ3mUZ98jblDISrmXozWWsxu4huih1MyRl7AMkQ1U0RDg8Yw1RmuB
Rmprqm3LvKmAoUQapdozSUUEbWODHAH/yNxX1kDjQVSb+FNyMXOlpWHlCJ9sysMwNsRRraGie2n1
lXgAIUbpThwwduiIRlG9cU3bw9jS4GLZQq7vVwMeFS1yVRWyoAO2MGybb9n057u9y+1fWrluP76T
NNM6HpbwWjDgjY+fgj47qaHWHRmpCtKFdGIGJ99mkKKvSl8Ui3D1jKMnroTxyXEhfBny9/5AOthm
0lyCA2FfRSHZJbNGeVUgBJ+HrgTu+C9+ffecaS1JKvG3KCwMl/BC0SZwzNw3dC35GnQF4vZAAXBz
Cq9TlDBqhMv5xyAUEL7p3MH7r9XsVRXP1elIJI52y4AcpqFDy6/GAc+XxJvqUUO2zigYIVAMZBoM
JaLTh792LiyD0y/vptyLq8rqMqb3QV1OnqS8DvLWQd7jC4iIFKwgJsBdfHap5kv/IcSMy4iXC9jD
qKP/cC9J7prLh02rL0DDSE957l2o7kc89P76PfpTYr6JRKXgtIIxy+vAJa9+9f6f1yOtiayuHvpB
ScjDkG5TRA2Vc8vBJmY24+hN0jBl9FlMv6zmM2hZpfKQ5b3Sbt0KVSszBQw9Bf5sq2Et3fo0OMKR
mcFwVT/pu9c8MfHY2nn2ETzL0aTDQ1RY8xyvMRT2TBCV3W7efmro13lNQU6ae17cdEBq5l46NcVx
la2BXtExejCEuQaV83ypCsNI9L0mStmfT5zpAU8m20g6OCF7L0tGqUIccGKzWJ/yz5XAuVaF5cP7
jPAqpnqj9p9+OhFA3kV4FLPfb2dweFoFhUvTZYhGjJo3daWpEGp6XpcBHHX60JrmhasmMhnOCG22
+kpJ4qexF+heBEmAKjHqRm9VGPGb5gQOu1mCc+RkBrfCUYc/od/AA2o6l7waAQr0CemOHPPM+NIj
3LyRYtEIvsHlEqV8ME7dPqdT5OtHom/5nvAem6TXIbrI5oS7n9z3L509VkBf81RzxgwWrceEi2A8
PcbEQFB7MLdBSqj6SITtdxHtoC4XJGstMy73cC4dU5/3DP0q3mWgcBsFFc9Q7C8S2AhOw9q2i9YS
ebIg2D5DXWbx1RpBuZcLJrDcuX5QGPcTguky9qSRuf50WrWAaO2VxJKn5/OQabEBfsXO7c7b3ZIe
SE3iEnYuKCJyemCC65mbDSwNI3Rm2XJuam0mrvF0+AtIZbFmZxzBZzWVloR6nEHtv4uKjDMGde8g
wafryqp7TjvP3v5Db1Ge4fTMTkQjoMjAipzRFtA4E5z6b9+GPQIzR45gHHplnxlbhZBuKaXsmACS
/oH3yeSe5JVdWzzkzZVNVCwHo14Zh2IUZCqFZNi7LAd6aksMt8AjC9TlPleXyQwhn8PwTqsY6Spq
IV2rozApC+AKPXqBs9JseehNaNlphU1tRgnM1yBAGzhtt0E5HULcorcOxYS+QnDwxr4kcimXex+t
7trO3jPc9AlfSAkphQZU9Jpg2D2P8dnwHwgfB5WyAxRfwXOO3vFAMCEAvohl9DrU1lYCtVQ1uVnJ
piubReyUIoBkrQzzw3Poqk+ko9GOA2KP1b4Ivs8KcnXys7XE0QoHcQm5dy7iVqmgI1psQHBMH67N
ydbpvwi9SGbz9Pb6Gofdko8T/u/eg7QoGSOc+RxwwrEZfFnuXppgWJ2sZZji8EcwOI+epBiGgGBT
nvvUsZvm+MsJ50PhW7IWBxNYgXSrV1KHGdW/WvMYLn0weFB+hkfysr8ihGGVx9YkkuSYs+MzWb+t
Q/0FJQ+SNHkrkeAEio25xEy2J+16fTMM4jQY2gpBrwEo+cgptBIwcQop10Vxr6/fqhAuER+16WKR
YxowpIuNGxErdattmJhCJVV6TeZIAMsLNrn7+6npL9QTZP4u/Sn8ELkYO+UPY7AM4tLHXV7lFoX2
J/vy7wVTiZgqzblRH2mEmFQkm7vjAb+A+fVysdfKKBrVzm9+CU+MNP3fIi2NYxRZhUeC4x1h+VjM
J1aKrQDnCdA8PqX7eqUNLZyGbZH3xerZ3cPeCOTe/t7ZCUDbe0UnYNX4HblMGFXN7Xb8EivW/kz/
5eHxXrAASbpWH6Py0hQVPAeO7VKKnLYkp5/+/C4i5TB2lyrAyXg3RBL9gtJgmT3wpDX7int30KrY
syorRaFNbcufVpZNsh7yTcEPjc5pCGA5ONpawYkDhLanm+r8I7gXlmceAgudUCo8iCVYYqRw8Pqh
87vok51N8PGXVxR4dfJbKspraFt/iAjkhp0189+NmhFSOjF/im1kG9AsDmWf06utzw9Mly1B4Tjz
kov8tjs4gnUVxdfpNF72zUy7ZWcLFQfPz1J7MG/BvBw0cF0U+kCcRn8QIxjlJh6DP/MULhForJT2
Pfil90BBALD1zSbY2oBdPB7CZ90Tp6yUyn8g/Lo6m3JLmcZGU1Jy7zElmM8bAcuHx2Z94LEAI3SB
ECJy5Y1/+3ZalHZurBCCHN01NktURKJC00wvk4am+R1LGRDIsW3fyt+dkidqq3kCBgccw8Wuzq8i
7SMQqk0ofQKYmg6H/wkuC66oSNCCjWGmTkbQg/VpMfDD1RQNuWis14oIoL9/Sw279Ubpaz3W4LXI
FO2a8vpBRz8RjMj55vVS5PRYYsA8xZyKLb7Vll7DtZFdSMPKnd5w1CzgenIenVaeT1tDvLHuMFqp
jnIy3XosqXPA9eyIuOdQJYXfyXdVqDl+6s+05EAtmZs43AygtYKGecyUhCg/TtFmBjXkV3NXTnRj
Bkc3yr9SaJDH7sLWASq9XyHfpPuxYPEMLudSdYiGTTfMKSY5E2saHsCIBDMLbjG3MJ/82t1NUryF
xEUxadfepmqJo4Hbt3H8y+cL+lMiG7yVhaaMs5Mn97mnVvsXATMKa1+tntaZIbkvLyLouXZhSahi
s+33dXpn4dcYyyabD3xatUkJR7Ci+j6mB8ZTmde9P8LqPGupCwZRz4NQgtKyM6mB7J3Y97vLDbRk
Jge7p9OuNTC1Rv+Ba1o0+Vc7ehhryRp/rd2/bmbHoxwzLXagZ06FsodsvKqvJDl4YybhNpP6sSTN
bkQBVM8WF/fd/lsrTcPyjGy4NbjVrwK4sdQ4p3nt8cHSUFo4G2sUAI5WW9Qkfg9No5+1dZypZagK
cFeWmYtg3bATx/ukAS6JeWhb0YfWiDqd71b/H8EHMM22a8nb0w7eae6CGTtkewRWZIOm0FE0Vt/8
jRFG5bWH4NTym14lTZpZ5uUj8Kpq2g3qZ2UIrSw2zQ/tbYZjuTZSMGeho9zAerDLQtycFGONUogj
6JllYTOGumDtgpGb4q99P5P2bv8RO8R2JbjywRLb/c2/NYmYNXQeWKnlMw86mN0QUYmhs6BjSKe4
PnwqrgXOv7oHh28Su39H2md3CMAzTv3ZuAW/F6J0peu7zoX5ohWzpCxqbSJo1HSlEEaKMWaHImPx
+F7QOoW1UJa40JqnCp5Gd1/PFIiz5z9TqatdAITisoj8C2HP8tNReDabuGYFPVPk3r6otlgPoX1V
PI24nkHkVzFSS0UfPc2DnvFBJirciv4ah9ouzelgmqC95qWoK/79YL68/+6RVCamhA6Dnww3g+Zy
3s2zMW3FdcgAieqfra1k7uoguiSmfhDO7O/vzcMR9IxpRFVoXEOAe4ippsVv2SsYHuZ48CPAkprl
TcS2YKDlVz9RzjAh1LFlWiayWtyjII0jVVIcyYvgmXy1DzMsxtaVczYHLR2FSEHWcE3GCchrPMlp
cJqBZTV62MpvBNJsNtJbXD/FlLA4Z+Sa8H34LmBeeajw4t+3TTiHMpent94hzuX2r/y9i6ZbP+e/
JGUafP4bvib7D7wMINiYp+GT+e3BsyNpNuuOpEgBvtsjxJwakIHNF0JptknEOs37AgKaBKymcHFr
Big6d4iRnDeznIRaldwF38lAoCzVrjVgqQ5w7EsLFICmy0OpyL3QUGkeEiKuNLqyONrdXW4jrYd9
onz4AC2bSmgyHSPghACm7rvl9w76Zd15NqI4A6Ht81B800PynwfY/8VkL4Va/klo1bmtWg2l3br0
W7pIqjv9t9VwI3Lg9yit5a9/osRd6svnqpuidUz6NRbF9p0KDzmcxSd3Kmx7JBIPe3pEGj9uXpmN
M73dtk8BGCYKhPsWSNDWOwTqivxy2H9hJn44Q64T+w9oL2JtfSQw/hNcQo5JiE9aQFdE5UZ/c6Di
brguqOrqlnFZBK9fKZntxIjZqpKHTuBsCByN+Yq3thhAeHpgZuYI8VRQYA7nbS0GdaILqQPIQyrB
rA828idPxEmyCLDI6EK/E4cXScSQ9MOT3dVDw6K+Rvg8MjpPGsaBFrZXdYsbzhj1d8TYjbIDlHpu
VFODzCgppwHNItiQXiiNSx5NxRzTyz0EZGiG4/VHmwkVJVDo/sYFeIdouKivNI4kmQkqBu9+65cD
pth42cEOMAU088b5e6AEN8fU6VPqjYF8FRsaS7ZlAwktvJlOvatcmMRWkb38/azjgnKapVwiyP+U
mjOC4SYnn3MsP/qOOKI2K+F0e2tkrKsuEsF8PNS3/Z/zIZlM9KwyKjtP4ctv2eYWPh/e57zxMA88
xlaP0eX+H6ne95VdLIqrgmTaa8rMz3+dbXjQXWtUK1yayEXne5FEBenBi92NKuN52uQyPRtdHMK3
fMv2sEgXxfihmg35WhDWgqGvNJJXYM7ngDVa5whztcOUDc1fqoBTJAmvpkPk/1SMcgPWCsBKEfSj
eaJM7aDBYhESEf7eemMppziVxGpHgQYUgrgH9UC4kz3wIePhJJLPyOXRljiOE6qaVWx2qIT0Bw0k
/kAaMmYsmQYKYfvTPZfrYcyVMHkl5MOx5UybHRrltgtQzsQnzRmDIAUG7fKYJgWVFFg2iAm7DXZv
vbM+KwTxLE9+Ow5eTpmsrjOvHjwzP+alHvw5sohASrE4rdisGSd4fQAhUvWwV9u7jQW65oqYnK8R
X69342Suwc0zKNKI5tgrDbZEstM8c414Y9VWueJA9w3eL85jiqPPoZsw4WJ/V88bS6JFcTDiPsxr
OOd3NKCbYEZW/HzO0RnoQ2CzE1haMLq6UbSBN+rdWeQtnEcbPwO3oYAD476MQW4hUm0vfv/JiFAA
PyGg6YFFCvIlxc29+FaOH75Bgw38oaHQP2STj2WsvnpAafAqx/VPuKNzepf3/hTduyJhlWuK3toA
CzBZyfKpBDo8/zR0v0MTCHGupr+R4lKmujn/Mheaj0wezv9muZ+G5ZqsCdcYNgaSYvkZWUFJO/xx
fSSm5dmoNOJl4Wayl2X9/rLSQ1Q5IYgFcURRq1bayhGCaVJkqrSQMBM1QzQt7KSw4lX4wx2x7n/+
swUaL8L+agsabq+VLiM9DxC3r5LCfcyXy9dW1b7UOJnVL5LYirapBUE0zpl3hQ2l8arVeygw7nw+
6L0iVzPh3qodcAtSDN+ft6kXOW8QgTgH+GepDdlXs3RqCMW9XT8r8GU0Kyrj56b2B/UxfFg9O0NL
WhZExAFSONj95mU7/CkZMaEQ3QG1Ljz3gEr3AYQVuh1OE7LoRmJhjGHR029JNhMA5jnt9UjHOLlr
ArEzecP66pdn4Le/b+KOUkIv7RRpHvXqSODTyBHM6sHTwsCkUBVeMMW9Wrht0D/ogtzz18D44PaH
PEMrjM8b69/buuVYk5ynK85NiUznh/g5t+DkGiEvtNB3mAMznVV3ynuhOSYwbk0DGl9ZBQ88Deju
vlkkbeZdeZCPNTlyL5KBn5/Xk71vyFHgb8ZP7XN0j8M0nP4855Hi6UxvIawHJ6PVLMZVzy2SWinf
DmCXwgFRzH9ncGiEcI97i4agax7PxOprCeg45rzYRjdFXHzVfVkP6SwA6DDmcpQzFTfWVLEb9sf+
d8bdEkiLE6xgVnAEmFo3cD6OnIAQmoVVziXZw0ZnNKB6+SoeqBl5PChlothmvfZHWexSyxs2fOIh
kio5v0bIXW/prMNp8kwBBKYUlelm0ED/w/ntmK0R/KDIa5hd/5CJGa0wgeLYRoo1kqahsWBlY2hj
oOUF+uDr5jXsC0mqTMkK2YKrRuwM2i2BArPTo7cYa3CZIEAK9+FgClKIfjoe9zjU+oXaPMxDc1da
bzi/CUUBasr5mFwS9YOMG6Q+a+CcCNmcLdkW+vR93GCKJooTSWCot8iOzVLZ7uLed7dCfUOMhcKo
8Ur/XhMkOjM5k/QNWFcqZVhMBHXoVfC3nHMnnO0oimMV0kCZKHSm/UrNUJaFI78JViMeud9tze7Y
4vAaqG3W29UaC/6x3gfEk/nW0oOKr0WRjdbLs0GDVD/ZYS9BjRxVYZPDwegFESYE9hGWAvdLZNtZ
RNjPvqRb7KjJtUWU1sNX/ZY92aLKbjsJEtKT4qomgCVNSk93EyyVXdLRtPE9rEVuyPxtVHduGtHI
u141Et165Zj95vdkxcoL5nwHJCfJtrGJOPW/CBpTu+wQny2qEY9+yfR7mEQUlI7wmKIel0IgPhAO
0TVWZLvEre9pOTgPQDkMJse0ccdLOU2W8el2ccrFrfGdcl7jUB85vUD/B9eRvuMOOF8dqtMZ4f9K
1yfAL+xd2f4TvLhegckqKICyQVTvYFIzqiAyUmVVu/LjUsmfM/i3o+axVwABKhGbyqhIdQh/FqLA
wXM8/NIFZZskmPD5vMOer3NcJAoFR/HCxWO/1xq53gPhe2sA8tcFnGRAmguywx3lwH1MDn2s0zGO
kYKqt3qf/q748YUtjP8DWWGcPrM/9xqwhq3lvy8T9TuMJHGdWZiVDSWHLl3RDybmtjJFG50OVNq6
/7v3dFyE0syr49eTrV1LXCB84v73n8/C1n35mS1fayJclLmsXmgFkTYEHcTHoc7aqWABMPUMhM9m
xNsgkUfr/U/YDUVqvQbj0dBuA8+8uu9RLbIETW331y5M6ApR4ALH/zNQue8xW9o3aSkE+xJ9MOp5
QaTSBrmA5sgPGtlxRr/RxoRUXl4Af1uj1aOxARpiFJpJ7EO5o2AANxZMcY1hEob9DCRxWM0/aKgf
DNtxMA4BnvtN+qrO35bxMJ7Lry1StWC8AlbPIMOYzpWVsE+a/123O7IHS71wYkh2u1Fk3mYDOOt3
O5QC8RpjAQYDurdmJhthF7PFXCG7KXUVH3U+8Pb7aAicA0CB6Ogn5MxMGljX8+AhbuvkKLyFcyei
qjCvSNH/BLF++zN5s/rBl+VTQA9WjAerIqHezl8QUrV7CxZV97flblVUeOEjiqxwHvcijqDfj5Op
ukIRGPqgmk9MSN+B/mfuZ+NhjDHk93PSHQxu8wZQc5mVznWf7P6CNJcYOB73uR+KLBdU35+XDcWl
nahPb4m6VkCXwTBVrRHBQHhAbdTCp0A9pKeQ7nadhsoOcyPPyNdG8XQ5wsSh5wBSc7PivleL2Sbd
31reRgmEUqX4eTOPUqQ+1SiXPIClbxwQpBEmAZtjLcKaGGCmLJo8QxOIvTIMCzw5Ymebr9dx2gsL
Z+llcIylAkJREhwQe2dkSOuMm/sWit+R4TkxmdTjTU63fjLfn2T+NutPY/fNdLCe5YEuF/cwgQvK
c6DGcjWtjHzweY/anti9xf5WadPmA154SAS1HXlKrKI0vikK7qQLOuJ3+NkoXWdfoiFyOr2hxq3v
tjGaao17WA1OwNqmJ6Mg4F+P1bLyOiS0Gtwui/8529S3Q25F7TsjbSQ3AFpKeV4ty8KB8xOdP9PO
CjLiB/2ei7zgPhSHVjJFHXCBuwvyH4QLD7tVPK0MHPhrhcgM9fhMetd1dZ/WXj0/J2esdrg/0QkU
QvWi/Fwe/8dAkrNcs3RX/4+kKQI6ycAlbQU0HxrtAN6KrHU3VxwCKQkrBOe9wZxBGDxrdyhsT5fF
Cistsp5SoHpDmVJRM0gJ483cSVQhB3/hQQfReZx0YLlXpRlDQlFy55CPdOfYFggOrvqv2K+/OxKq
s6smK+p15ypxX1hHMwWkOiWe8IMB/fI6IT4oszavnXt48WTvccIngjnVf4v+o65vwtS9/DMOJTc1
aKeHH1GAMnkygtMatXC/CP1TmFusV7CVTDWzE/W+JkmgF0MuX3X9UhWqctLFBDH7wtGZRvmtfX4w
8vvtXf2RI5wNSEQlFbSjtNtEA0+V8hBRhB7dUloDtN9EcNZBdnIcasnKwZsmgwEyQ/rfQOch91f0
Z7JgME/8qXK4CSykoNAaC2SSvLKHav7kmSExlNcdpz70CS1oi55zc+UkkoCWBdBYvUG2kbI9I42M
mqTQltE0QOQ9fyPA+r8VQQSL0GswIvERzzRe3E/wh6sSYuzpISjIek7XahZhSkk1XJb1bRG2fCmF
pnN3xAURDW1kidGhrpKDr4pgxXSBcDugRd9g6B0jq5uzRfvRP9XMOgSYFbtuHi1zVhlEgWD7QHZj
Pzbi0KT+lZEHMBoy73KE8IP5Dh9JVvIr33tXJoVcDCuUU2mFR04WIgf+P1OvfyKj/oUDhOG6LePr
GWyD98rJ6WdGeVi8U8DIjGwk/rTsLV1CKWY8pZDNy1f3WSRJK1j3uAUE3tE8t0ALg3/RPhm4CK6i
6DZvlXh1FE6SmQkmFzpGQIKVJ1iangQP6MZZvKUkib1HwNaEra99/zqfEfIx+vDqrjn2anX0BzfJ
az2ZNWVvmpuw+3AtS5xeT15mDg+6BKKMHPqSuuhh/XHymESG2UmpB+9zHVZavDOQUMmWJGutaAgG
1mC1vMZRRN1PBJst/rmMGpHHjhuG3gwCZv1IpBiOqHa47JFKg061ihhJU/exjJ/JY/Jhob/0rwJb
3xvjLo6o93JhapgoTuTd81NQwt1z4y6z0MY5AdX6G+s3xf8JdJyHfnvNYeWUQYIPsjYkzhv3dZYZ
AIInLw7f5pUEqj+qxFI+RXO5FUn/sFTG/BYu2+S4/oWe2wwAMUPP/SbQ879kaM86GVoMSiroJ4TW
g1bv7l2/4mOC9t8DN0L2lgKhyJzb3lsSBRvUVlNfWBvZTz+EUZoD0aUfKSUe4KqeQblSmbAAciUp
pTjCtIJogJZtSFViUooASEOrNP/mT8+AzhJnq1pQDKVuI57AmtaEZXltJxZo/EEmvEEFWUh/5DE/
xc4X/icuNv0cjjeJbSSM5U0SCuJ0jmNEK8nO2MyR/x0p/hrKceqk8qWNbA537ox2WCVr8UIIMRuX
kDkBAC0mT+0IMsk6e6bjdNG5LCptMF1he9HfiVTu/Gn6GpwOUASdKzsIkmU3M3XaUyLsTrunwwIJ
bTktTOyYOHmPcdpkaAKEPhpx9W23sR7DbAYWbbrSd7AbwZf84VH/GSG1LLsidcZ6yQSpDTnNeOaC
Zsdj3NJtWVHrFmC5yhusFb8TC0gJlLIvuv3ER4PTaDXXAkELHaznhfzRAkWny14opEEyhpfpCJCL
yeftGmpEMCAGQAQzve2EnBiXddgGd4S2jaW0AksNgmDpqTxRh2TvC2IU/v+6VLBskC4/e+lPSbX6
wr+80u/QHdsoMYCk8lkLEJ7WwE8//bwhSiAZH5fiOowvpd2piV+EyvFkKOaCHn0zZceqD5dbww7D
9N1KJzrzy46Ysxv9+YeXxSQvR3xzw5RShpbpgtfwC58JbroM9Q9ygcrbNwABq6fSP9iUsIQi/cJA
oRa/yHjwAf3moSnE1HINVfgF2TizKcKLzRBeEwmA+8U+yYseIx82FUG/4whdWvabfjyyBZ+ZFIP0
NscnIAgqh5uTgYU8I49AxrZAFgLMpGSqWbOaKR4njzc+9JlTb4wNlxNsM3EXo8KTmLSkUOYQuiDp
sR1hT8601bq3lwHiPETuJN7dHx2BUPxlgr0zVeapZyMhv8I7aomxk7QCpoEz8+7NbpHpiwJ59JAj
iPpRQ25bHEFxlu9ymqIi3A7ZDm3pVR3cXfFsXKMyYaMvi0Y7647cwgsJVVDpVLHdviSs7VgY1UtX
gFVpPG+DILglyzqKzAy6b0LHO+FCbpUZdMuooTyBUckbn+FK+qifcGNaPN64qfkoj9cyEAALglN6
Pd6isBX/dlf3FKS/M8LlpITmy4BM2LfbzAJ/RnZ2Vq6eEXsJ/TgiVFAphnPtnePPy96AhnVrh9g2
0ZaYr04/b8rHHzO7WLLoft1qG7V+EGoarT6+1k41rA4ZK9z2j+EbJ0dHvByjBPXW+mvMyi65ViAd
+phKAvK9Zv2AY0UBHizTUeB2tjuIowPhmMQdDVCCxuNr2caubdYrE7uCYoXCXLImx4SfEeZo20F+
43LDIrQT2xPmmfy6ppKpVcCWS+X0JWMEc2dMfGcVba94DB53aUj/jufGKNa3IYthOExRQWYTmaBc
4W+rMwYBUj1IGLeFb8RU7PwGB0aUEb8WTyMRrsedEij+gsJOMBJ0v5gwtLHcjPGro0qSNz1NEvEp
i725rSfK1vWu5i9EYDFRln8+jJuvsGb6FeCia6LYcim9VZvjaiP/3GdIwfvcWgcA/6xdDD6XGiKK
m0WQNbm946J4XgJQe2OjUt25ReSoGdI2rHjOi20THJTW6cUMI30ZdzFO/00KuIYcUTsMHPUidVXM
sotXqg5GQwWrZWFojS5scuuG+0WA2EN4Hterj8WRaO/FVQ5AJmWO6t16N0TbcCARxkb2WbDT+G7V
WV3nlYxCoYsdFdbw4sxgHreAzvfQh+DJO8iXZ6UZFt8lZMjtYjHQTuQSamHN1l7uKmVOwBjnMsp4
Iikfb7K1bL6q1u6U/uxqQ3iQE/jHWx8yB5bj76kvW2m5EgNmakvURb77TORQtGvDl/rvSLL95IoE
NEEQb3gHD2tTEmnVoIJrtFtHGub0Ae1SvKiK8TPwBU6MfEDCa9CcuwB8zftTQsyB9Kn0pxRnPsom
x7mXbPdq+h/FMUE71fv8caZFWE+3ALh/5Aw6Xj+BMdv/eVXAsjewDMhVRqrn6fOuovY933AvCN+X
VXRqjAub9S/2t6uwJ/qLr5HYiuLM0ieGJJc5YKaqJYdRPW+57s/NGsyA5mAvFtPVHjbps/QWFoVO
RTn1gdYhWmuO4hCtRQDviC1SSxKtU+neLlH9xCrDhggdXc8dZm0whJGQckC4IDp2ikIhyfCp4Xyv
X5IuFIm5F4MqiwPFbUoTTC4XGNUxmukai7fUrwFM+iQGEVH+NJQ6YHx5Nv/Tiyj8Fzd3Q268yGXj
x0YO+606lGM3+jp5XedvQE9piH1KWTJj7/t8tZMqM1m3IdAU5+XRGUUFG/rAg33/Z//IxcvptnzE
Ze5um+Y0PZKnn0e2BJj+JhFR9D9LmDWv1wUQ3jlsXaRxch26Hk8E6LenSs9owJxIBDN0v2jcFeKb
uMoH1YgxGjBwt9SasxpE0HXVc5N9FhGRmws8cc4kspxkRTrqsTg+MG5HV/IfQ4rJpmJ4dMQfNOvk
5A4zDQ0HQ/NIbJbcdI0MKTWHcK3sUIXKVGak8U/169z1ifZqnqzqrOaV2VURfB6IHhV4NLGOvTWc
PLEAa8+GzAlAoXb6cTUr69kSa8T+DUrI6Rqb2mjru8pn/zqnH5Q7xm9P/W4atG2LcaNF9ENv2sa0
UbPXuSAM8zwUAr9zeDyim+GAzhYROW288lQxk4IDDNgcUSHn2Ih13zmQeeKGHK2Hw3jSpO+pDdVU
C0wcU4MW1guGnOTkssseq9eSH7zHa4lxJrKBS+jakbt9rL4wx+WpPYBK5ou7Eq4zcSf+VmJAJ3q1
J/v/wU5XEOo1avNlMC24MurIXFXm5jcpS7Dpi4oYYqQG5KtoZAbAFkyKeVaRMA2IPC98yQI4Cdi6
4wIp7W3reDyGNgtfS+mv3F06ewRuqGaB6umWVgVC6VbzKmsUCGQi76Z+dXomHd6kK4szJd6v9icV
parPB6kBkz1iTt4bbBENboJQjTUi/V7UhYsc60ZEBVLsSMWvqk0OswUSiO7ruoYBusLgqqYEfgwC
MtIL+r+6tN2tPg19fqVVFeFYqR5aCRjCYoEsFCtZly3OSmo7GjkZC6Q4DsiBLH/aDipaoNYcH/W6
x6tTNtrECRmPkyQrNG1qiAR8wU3F4H1jFadKFuILubmokViKwFdbyeai/LfPxrrRTvgHTFnxkdnL
mfTJZetXASrCNPcMIvzyULTjGKyruhRwPin2g/M2Z/ScO46KNdc/n07mjVfM/qVYy/pvnj0ph+Wj
zNEbEI3+eXCLtxdXqJq6gnKySy41m25llSKU0kxuV8jFbtgEE5Izkp2MZr2xvrfIyyQO3hWUNXrO
L0BoCR+/0xCqrmO18S8pX610A8BSUQK6R1jZc1PRWZNX7EenWUTL2G2HSP9cVgk4vLyVqYvVTQ7E
5KL1QRMTBzzSIlwK2lgyfLiCrMxQcQIUd62MXRl4AuRQiY6I9VZOFvPrJtC9xDKEfK1WowvamcPX
0Wpuf2XCZZvHLDRu/T92ntVunJCAf4jn/HdxwWvIygk4mesI0ldgnXOlu51E66MuhkDqy+eJ66IP
JiObHf5ZaJ6XYtpkvJBrWp3dbDE0DfeprQmEJCPm039AvHhi+ph6Fn0cBWinodD4lAKU6f3+KimH
DREJW+01kIrtHzmQPg99sw4VY8p7aKflPwKmzCrMteWwvFSznlw4qqzhogoG6tKz31Qs/rKbwSXE
8470E88jMBJojrUUVYbwO1nykXwOy1xcYLBrSuLfQLMIrYOSAsIGQjHMqas6kJJs0amSrIgZHF1f
jpQY3XMWA8Ob6cai07yo5u1mrdmBpQ0kZxIXp1p5f23CkxKCEteDMkDcqa8//nbEqJZsB2rGaJls
YH7BR5LWe96GFkP7BAwxc4e96C0BbUHBK7mLGuqqlUAHeCr2UICzDno1qScn6iSU+QX4uROxqFaG
lJ4653ywQ7UHyY5PsCkvDTKcTTcz7lFIi3jty9SP28wE7Fw3LHhj83vfw8xLFlOrwW9wTSEfg5Mq
5Y/h5cM4bY6xnHydRhCwgCml3mmAVyYijNKx5adFaIBAMibFLTI6K4L/9MLbX+spjY/vMCLQAA4+
H3yrAMAzNWAaubhSoXDphF6YyTmuuvx1EKGrb98eopIT3aObbaaDev/LYb39Lt+PJ5GAVkQt/plJ
FBdSz24pq7LpTCVyNBp+rhdLrSW79gAWQnRuFYzFASHpAIK/UVYmp9JmDS2UbRnAXvPcCaJMrlHh
1uLqQdmI/qs7JHdJ9DBIy0VmPrdvMDKSInERnJlTrqLFpCNQuPuc3rWrA5ka0/gg9dacSt2vlio1
qVBoF+FVeyNp277OmMhnkissTJp4VWP105wNLFlCPWxQRRgBO1UbmClks6xKXrIi+3UKXJVSmdT7
+RCkZPrbw6mS9+tA+wSFA/lXr8ZjEd9TcDTUM/QUaB3iUhwnO9elkIr8nH6kyEyqn4mR4GG/q8ym
KlICvo42znTCQmpPm09jfr6YpSmTYHxj+MHadC6Wxz5v88oi+CKu0o5Ia77Gbv7/TOpjgfVKLxOD
8hr2p7qL2aF253vnbvuyBOi4njFIYhJoglSwMwb499lLTW4HuAT+a9mfUS1oHmspPrXEIMsCI71F
MDhUuWuI1o/WC5QKYids9vbIT5BB+gQfoC2Z4aPrfT5E9GSdW7RJ8jJctn+o2Jfy14MmgJVYbgVN
tzPPcmXRSpYp/wLbKy7MZ2pFz3JmyitNmwlKWrfiWXHe3AEqjtbdXyGKXDxlo9B7C968vDXKcDD6
WjQJMMPNk4pFTSfcJkBsB/6MRMoxv+qjb4ZZrJlW9hhsGDxCRR+SYZlBU0z4zzQvfHdyuNtgw2e6
WaTwO/vYQkrZ1/7fESUuTTdMyu14K1eNSJfvkxvwwnSf9dnnTiICmTJgTM9pM4/eb2bGznCC14SK
/hBQi0xRThZwNsNuOimjNSt3KN/Th3yv5eoSRnTys+jzVzfxK4se3yhgx8HFa9HQd71EqA25xjBa
NI6M9gMdrPhuInPrwfBaBp+Xfc5EOcHrXFRyOj6Lwx25sJB9MuaG8chFsH16LqPMqs7lgTrfTP8E
CUGG+JFS8zeXz4COhqg7vmpo7cn7oLueNfWJNB2tm6bD2d1/o2sx1sbVt3RXZ9+WMwTU15WIwSpm
8bBO2e7zHRgLlx2sZ1PJG9E6Tq+oiVW6zNk4E9q/xubHzBtBVR1SBXSmiJsVK0HbknqI1VHZtl1M
7YFWq6U449wFn5BAv1EE3zhbF+UlLY9A06D079QSusvl5LSzC2akhqzNQRvWqu+rjf1VjiCi3zC1
irgvw7tzrhzQiCLczx+uqjmIw02cljnafExOjEg/OJOPzi3qyBh4A3Hcbwz7EKwMZPF2vzyTz5SG
DuD/Qp62R80RZl320UNfGAil9boaKjbi8VqrI9Fz8TChP+m7kF6IaNR6yHfpFtWhcK1DNd2/sN/c
fxU33INSEVAyVQGEB8SCU5Y2ti2zz78Cx1M6iYtHyV5/cfqVaXOI7WA2bpMtl41I4fnVLjHHVOsf
iLG5ULSEMivOYEw5vw1I4ar7YboBZ1vRtU4fyNbvO52YoGUGYikc6KkxKFrQVpOsfTeC+5kRTnTI
U5/8T37Y1370mD4A+wywTl8E5UfOTiYUcwoff6Kfu6JfAgcBWXE6boeWU/oaNq768tWHZzycDI67
qRWXIFY+QnTcS1xZL58+TQd8vuS/N90ns6cT+7wBxNwPX3Z/QPTMFL5jO9V6lwg0H/M41C+PEkX+
a5TQJrDLkmFAMWUiFxVQ4J1R83vZEdIifPzgRGu2MClPQ0nTpCVbHltFG2T4aTAcglCzGnrFhdeW
4KyTC9Ap0OaCojeD9uQbrIPA/XjglwAojw+uQ2EbWkKaWfB6wTGf3RKk1+4eE+OpVZURbDWxb01b
s1xst8jcpzjVyz+LP7slQwKhQ6WR+VkIlSicqIGhdMgfjY9sjAko800/4xoZAKpL2cInt9NcBXlZ
X77EvEwZtLJ1l3NRx7/bNRtBSeHeexByiDkMsrVnrntz1TS+zzB/Rjd8XGRXUJS/HzQzF1CKJRLn
s4Gl0s1gL5ETq9v2Fzc/pR5jHXNrVoMT3dXnGAHD0lHYcsdmxDx3atO+KoJZDqAsvNlI/s1CoQqQ
muixxWFdzWkOy0NHGTn5jccx5xI0jR1+PXEdfHk5wj9nT+u1r25KhOoUfoK5HOU/9bh6JHunsG5e
N9XwjdFfKsi/KC+QU3rI8hVBBTRE52rXkYFS+TvoNlRHNUDmDCguI4JYtHYGWBy2CRAEgQFnQBUg
9lpLs+e+k4eJvB9lxD6Zvemc4kvoOFCMzz2WF54Ke8vT27VmUaEMUJgVgTAZw8+yeZmqqZXfZzS3
ZsszCWAYKNemEo/hKoEO3AbUZ+FrouWgukYNnbKpV0oKHD55f7QHmZlIIA7ZJeEY8s4YtFjILkSS
WQ0bp6qrcdVBO6cl9wKPh2Je3sAv29g+rnR0VtuatEYc2Al9xWsEtOvpLAG5vDdlt29joyKpajlM
xETitgXiPjIRMvoEqNKUNhrzuf3ZsO8hEa/GcPXmOdcxHSz1YaBFZH2GjB8jGZCEWayLhcxBSr59
fg3nBfntVXQ0/3BARWzOQbjSHUUctg4vQRo2+1N9cxR/bendQuPXqL4FDlSR3LYUja3ldv06PUsP
eGyUMenjOR+poFst1IM0G4g0Zbv6m8ejH16/HfMdEjDiQw9bfKaTswtyQ0WZyrmN/WC4uWgvgeUw
IR2d1bOVrf8g6acWkA3p/lB2Jt2y2P4r9GlZVbnPb0ZhQmmLBwZHNuR9gJBuT1ZvswoLqxnabWeq
z24C8ShbGMFu1WjbIv4NLVB1ZkHYC/3n+ZVIX8mDa3iJPNLFwejRbBu4OwLrOgfZdmTsrJIQn6sD
VdZviIMW+NJ74WPVPcKA1E7lRVDBv8HgDyyuIPeONw1Thl1DCOPeWSWs2k1T7RWBDZwAbU+5OFRH
lEcYTb3w2DWoi8iqoce4JvquBgnhA0WZgty+mRzrXA1uNTIpxpL1M1N3OanrRasWF7wVzyI5zIxq
SIgFZ0EsG3xo/NRpA0Tfi7eknZLF7R+pb8Lnm+IkOYYiByveK/UxQRev5BPp8xS4VzKrukPgSxvu
CBgQPq8C9b41PKBGblB4G2nkU/iykHMtrcOKn9CFFV7hxQ1PqvPnRk03nCPQPcPj3LJ+Yl1eb8U+
u0W4I/eACqPB4UAPu/3B9nBz5UpuiK0waUZI0yaodqrzJ8e44ul5FqS2BHCPX7PdXRlppD9Rr3Lg
vtIxHnKf46OjujfC/MctC1+1bioBCELPrAaUCQ4hzmOKPBGH/84/n73t0awBwX7DiXaxnSxzWUlW
S+PTouHd738ZDvJRu3EOGR76Ui7vBrWh/FuvKSQA1krhEWwwU7HikL+SyWYfyt40omtmndj6CRT9
ozBoBUl1rSm4wNPe/4gYYDArJBnbta5wz5T9DbK+8As7UWv0wer6wjUGC67lqGDVzojkc+rXqN+W
ZNO+H+WOt15s2JHSnTLkt3fVUwNoPRztGkVN7zyov4e/0+svo/q9JEZ3Bba4QHv5UYEOMyJnja6G
PHhAc59oVcvsOCf09XONRMZVOcyGLmYiwvQWMfBOyD+wVuP5CWBrBqiThZTobXhmFESX5YzAIIwH
r7H2ITuJM/0gnoauy8yPnJ3w91geZN5CNQ5XtDmvPFUi0+dH+J7qXuymcwLrM+/oM5/H3sQ5Aaya
at0e0o/0l3D86bYkUCDnibNwvX80nC00faInZuaPrH8qBVx2JpftyOP+dAtCUWUKo0xhckwF9COW
QP+UEBVmtUTKwTMSb0HNZ5pDTkhhaFRDn7hlTjE7ZyW8wbYZOup8Mc0ns3zrWGcYBIjL56/NrLtp
DHKnqn+0NfnX7RuoN1QWVdascyZpBFd8Wgn0+R3P8U/kBeK+/u31GQrz5i91d7rz3K3Fl8L96xuP
RT3U/hVfhKmcQ1nnv9++LDzducyb3VdRIo2yc/lJIvdL4AjKmeqj+m2L6NZDTjD1cQQEq1F7R77p
KNffX9FuFA8Q4c+jQgnNAx9zBABXsyFuBdr8EsR9VEd5GcGS8TwfYzFLnhfuaFdYonh2MbTMP8Gn
ETKrtcEetk9s0dxqS0ejDtLtv6S8prtdkE/wXhZ7SslPAbwC5GxdwaLQu3hBs5N57s/hf+g5fWmU
TrBFWRX4+0s0crreuQCU+c2420aplUF/XxHf376NHZw4SZp7E/LVidAItxAHZT+SPIlu6TqDpACo
BJYI0qmZeDIHj+5F693jBDNBYA0Dz7O8D1mQLUvVSr3pipMk5Ji7Y9EtMhh1qSHcZS664f9wPh9k
QO36vlouFRkNaTB3hnYcpsMkg2lLnQxi61zu6BEthALPaFB458TWWLbpfHNg7WVwOGnFDvPr/M67
U48w9XyiY3l6PtDUbq1FmoMmNKlbYXeg2JDc+dUWvCHvr8sjEghMK6PFIlUXpW/DyMLw+sXKalKd
RpjYhuQUaNz2rkWYmuxImUyS2dqVQRb3tnHFB87/ITh+eZqtueVekxEEqEH09tKkO9mpLDl3klQI
6wzE/geLqJH1OS0gAmgoLygz9vrXs9Vi0ItjldIQ+wxJAVekmVbpPncwRgnoEEsNBOhrCJkQsS2O
wsiQ9kyU69FAohLTv14U/WSwwX3nDkOHiC4BdxpVSM5MQai/wEUFXpnN6Jj5tuxvXdFyOLLm9BlV
29nE+hbOk6YbPHQLkYCTaKjaNMhS9VHQ7W4lSsklMlx2Y+9UtA+lV2m47ZwQ1IE772npIoNnlZ6a
OwyV9LT1+OcUwxjH/xDXS3sF0gRFnYy7HbV6nA2dtK3FeEeGwCU/d2FbR4wfPGNUQC188HBe2mwU
lM0KpV+wKDC01oJS1X4wGy3eAbQ7gMK6/5/vYwUkIvzGhvyow7WrDV7zf7bvrjwEqooIS4RsKjtB
SWjokRkteesaZsiCKF5hMWwYRxXpEwpg6NR+5Bdt10ix/f6moqh4bEdzJW6X1Y4RPd1+O2dgp8oJ
WFjG7nWQDVrcR6p23OxutMFfN0t5eF/3IDYMiZzJ+pBVEv5fOqstbTGK7mXIMXOyOL3bpGET/08V
h5b920E/PVxLzIrD/k7x2q3ALcNAth644XqQ1yjAhAD2aG0q04a59X0S9uF0jwc6/68sdoAZA2Iu
VhLOWSNH5SLibHmvw5xvKiEkNRFhBjeIsOOPENTk5zMfkyTTOnTUnCP2MJ9z2VcwSknWy3Y/oLZQ
wNxCwH7ZX3/AG7AFm6o2sPED29BtHy10evRPbgKNBaIHz9FM5vYCaqn2apHQqvPVVKu++XFae+rV
qE4PIKFizmhh/5xfIKhtlEcHMJlRfHdhFUizQcf7UM29SgOXDVCv9/BhlViPDXtnLcQuVBBnw/Yx
AfiiIpYPxxCX3i0eb3yflYrv+fV6W53u7H1iuSodBCi3A2cmd06nnMcEwKldRC3YL7+ZLVxW9nXz
LcPmTUB+xMH6MPpeWfgS9Pn60cQC9zUgDh0tYOqpQcNHFwP1ubY/hW0lNmv8tYOaV7UraEtC1U+9
d+CwtDJpGqmOtNEk/CWmu5aoPYzQPmrah9brV7NZWp/kibgLzcZr6varLM2h/f+uyh+clnckZF69
uEIuyD57r6c1JeZUEY2l0h7nXcxrBdOPSpdCwAuBAtKqZ8bHKKOwNpzOOlYzjcaxLSY5dxpkOxe/
rYUr9oTwFfy31NkxdrWuomHXSPoa8d/F9dDatXhQml/i8bE7xV4qjx+0/oWDva7bj5W8XVludlrq
pJvPcRIv4aqFlb2Jv4IChjmpD3rZvMOTQONGodx7ugoQLmlbDzrsoBAmbzpSVmP8K4ozyNuBm3q8
DOuXt8j+MjutQq4uPYTPhEfZSJh6mUUD6StnDU/5Io2pnqmBAKrfAKY/Lfq1qMhx3812eLjsQlk3
6KwAospzx7c9LdbsmAMJeKXEUY2ZvnClSo78weihVt2d6ZP1SXL4u9WBy2mQm/sWNxxJvE+giYZZ
7b7qMi3g/9SlEBlKvQX7TURmTIpcupJgyWyldkldd833DcRecan8JxLDX+ANY3uQuxleCsy1Gd24
0mho6twLyAGEzAPEYi/5JycjrW3vHCvhVS3e6KOnOOq6Z2n6Bsh4qFq9oz8ejEBsHs0ydk4pxinI
s+lS5nDSBBYHzdtiDGYyRflAq82h5tVm5j/rxIn0MziJJ+s/Qfu4nKTOl2kdvz9akQSXWiwSWiQG
1AlT1eLBRAthC1vsBnC2VYblljshe8KZREZe7kOP1ecoLjbTOeRQ7TGOTDydFSkApKUyh4M8wPtx
DL+XcBv/AcSKERoxe5g6bEcqS3vgbjmiBzb6buS3sfXsvNXPy1HiNsMEv0Cd3xA2D7iaGdWUd8+P
znJp+McdwfamPL/rzjRQ8LtsU5JBFIp7m3S1P4i10fkJXV3v32XRf++V/0xI27s/bmxbALzPC2Jp
mxAxQ0qCxlOo42Uw6ChuF2DEc5LwUoFfYHVi3z68bPH8FzkzcSDbMdxVlKZMSW5Z8Lr2FMi2ZaIr
mBi3Aq9FPZwyaxnYunUsvpim3IKpD2/6YHjw5A9UVMYkq/MoR+IcWh89mD3FcJvvnx4z7SsmW2W5
qfZUUxX5A1tdeYebiW4Ab51J28mcyJ2Bt9UYAiH0q8NlFvoBPV/5ut3H8s2K2BH7vx5Zb5hAuOmE
tmeGqPJXsrMsHd5PaZggoa4yWk2yld62UHXF9Xq6/FUK8liKQaNUu2/mdy/JVutitlfLW0e3/Ex5
mzFw1OE+Z9Lhgg/9BggC5rjtYMXseaYuGTlzfYgV5HZ/zgHyuIBabgS2T78Ya8y7JMe+zb5fPU93
+Gbt01NNjxvIS7dkaoqFsAV6u8KeQIVssCeO2vNfy6LmzdB1r8GmY1fK2OkKbFGo09tQ5D6dDMpo
8nKjmbfxu5CuUeA9fVs8Jh24v8idIWckK6e9tmcKN3vqw+ZYhkf6P5U1tO0hHiGFJQdWXlKGsoDn
UaTwfQitCJbJJkb/oQkIWPyplBtRvEvyo+PZAu+xY5V2J7MPuP5JNWS+VNdz3BEdWVQp6lnh7q56
kKEp2iYhQk48TsUwDZ170L2xuQbfXQB7RXPB0D/rwOSMVxPtSCUNcHKSSALcBbnNxMrEaobe36bx
yK4BEKl+Ylh1g47vgWtEQI8MV8y3Tz3mrwL7yNcnY/4jHSz2wk3KDjHhcBlFzp6563tdoU0Sv1tD
H5XIH0iyXFlMIeccg51CnxRecfDBEb9KkriteCyKW/34VTQjvT0szSKlJ7pRiFKDn5Z6nO0BBt+h
qJ7IQx4p96+BhSaUk8OCojrCTHh9/vk0s1PVdWmiv5A5TIA1xJm20GbNF5GNKNdwDdYEBzNvAq8A
rI4QvmfWe8ohpzZS4Qo1wgkNRxZCisKgigksQ+yO5TrnLFgaNCU0Td+J+UGF/Ok+JYDtpJE1D+vn
w/2Q/WZ4a8vhQimLzRxcVtjtwQpixU9QHbZpZP6mrqlvYb4lTMIIx9QqkDaBBb/QWpwWkO0h2fxF
2mO6yuNZaEU3Al2UZLeD++OnP+mJ9GZK2vBp0nR++duR1sx9/OsW0jrAC/oRly/W20hbg0XRDq7K
B+cBzD65sGhsGbAWAiPAwoq7lzRdQ6d2VXuicK6EuZhl2Hc3R2kLQlcLGCAKzS/HWDKTW5y31huU
AIRYQ8eOd7ke/tB5VwnjWIOoR39zVdPEmn+DS9iSm0i79FCb1KAlqoZnmUpUqdXqt29mMA4p/s+N
5O192m3ByWLEactRmnje/13mdzKu5F0E2qui6hJp+/xxO++BC9f/gEaU5fMAwWrgiisD8ITWx2Pw
3dweVxLVQGnROGPtvCI3S8RG4Ovv+ZpwIsZ2IAmrlEKhG40S9YHtr1WQUlukEVpYKxuQyQajycwn
NjCrlr6fcVOGf4YX+AGKD/nXe6NWq6/+HkD5J5IeuPtYH5FZABilsVyTmPses09l9Cf/0aq+CPjD
D8ZLIBPgjMToYdKkigd7p3n7ni/Pb/b05c9CsFx7U2cqxQXRUVYqN16VL8yF+5jC6lgjozjcQQYK
gRhShAQQVclITaMB3cgfvm9twNoEa5nMHmciKQBe7wg1wYP1yUwhCjSILuMFmkDQzSD+TxYgI6xi
spDAsjGXOfbhq0kOLnnBilTynjSc6wfavlpx/Tm57Ayyb2oVFPM/LC+8C80X5hEGyz79EXqR7kfr
i9VuY7CNxgGJl1X7Q28vOdd42oGX6ToQ3XPBNjjiP/44Pvtd1kZ8ucsKxbiMltUy3OSKSamsRUKC
UL+1qR1FQibgC6ufDvxRB6I0g96pZ6QRJfVTnXy0dHfO+2RyaWqWPTx88FRjIi/NQDvnURarKEXy
60mm7Tqa2b+POuBZd3uxsfe+QoBtPhHW9pDVxF9XulXLhtNm4Sd/wesBgoaVjJHpYogHPRBJB4Cq
pe6lsnTyiUtLWAJjbiTRv3kQeoh2E/mEOCvHY6XuNBT5oJeBPdXq1GDQ73HnVHVDuj6pC1IEtuMO
HueTqh3CoH5mL6jiW15XOuMJ3t97qLGDtLAHhpu/DyEkjorAmEob+ssw6eoyA2OlccHkYSzLSHz+
fAwAwrBF3jDTLUeS9OXHzm0Bg+ROXBJzy2QiF2iqnHo77CJGqNIhKWFkDFBRNJtVtQaI23qbz8lF
19mzZMeLLMKb+Sy7oI0FWr/9qCsDG0cK9kmeL1ueaw+BhrAd1wjXJkz9iJTuUKTQQjfBkR7Ra6KY
5caBdVn4F1HBdDqjWm0AR9epizmMAMJnwEZ9WP2UW1mszHSKkmVX7og4qRCYkl4/Tc0wHd6d4nHV
seM7m97/gNSkpfexI1vld0tHGIZDEBXHuqQJAj4kBd3/MTVI7ByvIVp+pPBqM33BkMbue3XSyhBa
PJ189nXjPtJbtJahMuOFqABNeSSyakJV5LblBRxusZtv8XGEFV975KsI4rwfffzxkmUT0jSjgCLv
QMloEIUy54+GsGy6d7V8rypDlSbLgPubDdRXwdUSurHcL1FKLEaKci1uAJTdQPXtSm+nO8nVsEwZ
rNKnqd2Sk0l7yvoIYTvVs+P2YV2cbdJw2HnppBELwVK/u9KDRcE7MqvCB4xx6k3pYE+TQZfTL/d9
vdi712C2DXQVgemguc1QWdXaLYlBPEyAY07uMU8FrqmR/NCmV4mVlrs+JRl4Zg37k/iMNXlNMUPN
Ad74yth4NRdpLne2/ucuyzW/k8wRJchAwW1u8kfKMtty2Ga2DHda5ol1NV0Q52HyYIwaKiTwopzT
GjJRKU2u0A3Nhcseh6JG7TAtR5DjQGal2WSbR5DXOW+gWW6H4pG4gM11wfOjSimGm2EFQO2jjAlF
+iF+/ajkEwmpz2x3llnPvfAj4kXS0RbeU7t6PbNgTIMsyOS/eiALbSIBcLyt5Qcg+nWAJQm0OFnr
cPbzoeUS/ktl/OSrXez5MwKqW6wfsKrA8cnDRuVaOVK+j19BpaXZBN823EE/Ep4O09p9Q8q5jp6R
g4SlrZwlmkN7VW3CiDb4/ivXGB38LIN7U//Mrf8kLswi6TszdUuak/7/zUtKYUVwELluQE7fvwdR
MUZ+Y8jCcDbKbaqnQgA/46fpjdsm7XxZ8a75kqv+qgg+LnHdLG9bja9izmWmmOVUkmbxWAel89L7
KIbdLZDzZV/MV3JFEDWj97u54zqicEW93Ug254BDPxJOQdHYNxm5xgc0H6evkCmrv0hHdAQDH1Fm
YRhB/0kahuBlNE7pnEzKMWNATDsZX5EhyVPLWTLymUGMIA+xGnaoTR848NuQgEEUxN43GGdScE2h
9I9FQecTp40E5HNEw0EPFWBjApPHU43unzrp9/mXjlhHOBm+YDtZvHSQLEL+ng90caED8bbd+JQV
iWOHqc20Y9ZgdCzindrVkWK5fzU1pjQ9G2Zckeg3/uAgHpXU8h+scbo2PmXvamy9S/L/KShEP8n7
SRAidOXVLBdaE9MpL/m9Qx4y+HXdYeu9z0QrhAxXrA3jrN1eDpiGFLBTRGuxiRRTMZDByDfifqCm
ujeeve9ejZZpbfEdNUs177En1ci5+fCvZbLV4hhUNfCo0C4S4f59J+sq/HQeZn82l7AsYLBeZQCr
XARKZf1yYKzu5X++Pk1VNSLQMy7GIwctTAl0apbxInkS167kyhceXF+ntG1tQA4UBF9pVQaoyE+L
JSslbfOxRy5KjcIv7P6rDZLlqSpzzop6clQUdvo12MjzGgpf3DxMFZ/QF5JgnHe/aa2flm2et5Nz
HlkwtIi2eDBkM/d476tT1zsfeEnR5skyrPHxk+c12Mi6cqvghcp8ux57kgfDzq2NriKDHCcQ6zlZ
wH31Mi9jTaBD2oxrFampk5bL/tF/NslMzO7V0MMAWNecU07lxosSdtJfN7LniNXx4aJeX1D+g2o0
62SZhtCA6z/4cAdQwIf99MWZ9WF2Yyhn5AnRSK9r+rWOjCQ14vbCKqbvY8Kp35kDizvu+xmj4TXA
hrDqMmrfj3k8uP4PobrmNs+lyIaGr7heUEG8tyD5aChbdlcXYl43mDbwqd2L7NRjIKW3ULkrOJob
ZQ5BAthkNSd3M1SZ0q3gMKB6o/EzHWKDbmWw2sDbG5bXQ+tOpS+aY1jgI8smwqz8t+6JFUmE/p8K
PHNFibKUTo/8nnGfQsGwMWgN4tZKroeR8QYHAG+X6XDR0HYHWo//F5WF6QzY4TQIiwvnwJBiFfG4
tDROLG+4fRTTqS6upkO4zyXFYKICi/p2i+MY62qspecN2jYRK+HFJuVC1MrVSAgbg8bD0CSQscek
yUlY5rqbwLg+uR2IcbZ4DJGb+ddIwNhcAsHcngmf3wyHGlFK+imOzBN2opXtAk/+eZ5+CS8Cn2iD
t8TYq8KPS0K0P1z4glUcoWA3ss1t9lGfRTG6ct2Z/KgvI0YlShKKoVDAf3e4Tvi4X1Xq6ibeNpwn
t09jqmswOvvJRNSidgTnPNkI+FuN/UFt9S6J6wz8kKTj3Rt4VVteH3osh+Lwu2IUUIUKZvR7JBRD
xdNlbVRjObRV/GdHItXs3SeZsEvzET8jdy+vzXMyIGSybgjVzdgWQ/npSuht6B1cZlTPJGiv2Rqz
1Ewufb1Bw6Q7oIZfLS1UOeIPJqvnQ71BZ7RadjzCZ+fQo442z0d5F55kSRoTQe+iiM+koCVG6paI
61MKsPBNhhCp7FfPDJOA6wAImzpWdTocXqNJC3HXdGtKuXUNlOfH3N+57MVH+kLTV3/rniDSNjZH
YwVFd2T8YMPYtFYig5vr92dKeMEdF+bxTHPnBvX9bQxewUAA2gEeBbwgS+PCAF109zudo3/bZEGK
6pHP4cY6T/Qo8JbSdGzl0Z1q88xcrq5YS19WnVFjFzh1X13KB/IsPI0XOBp7toyGatg+LNqIvrkP
AXFFc2eyrb+qem5RswxNNx3BlEooh0MkcjcJ4bGydeP5Tl8HINWWsv31GfXpH/k8fSLAwXE5QTaF
p22QoiFkvLHrZLB9kwbE1npT0M0flu7/DNmgftrRA0Iy6Lx5knN+o6IE1/nVtSVH8Bu7daLTA+rI
WzZ1l/ltu6bfMSNQuHINtoB9122PlF6NgN1mwSsbuPNjBjUdc3ruset/S/wHh4d4os0qQVEXHnuh
y8AhCbkYxeq4rk6w/l2ICLRRlPU73vZGyV/AozhdbapxtO+dVzrqyw+LEMm9rI4gKk5M36Fo31Fl
j3ggclCgOc0QsiTMSgpDrJ3oQOOtJhEPZjlIn/7OwNmhw8N6NR07jDjcUJ2tOh8yY5jCilRYWGBT
XxaroiRxps44xUoo14VVi9wa9ybMNSfPoJy2GnU6z4U86B/sNC4yZsOe5+R2x+2ij5rLmot2MVPK
GMojrObWcbJ1kxNfEdh60oMJiCHGcls1rziXeAz+NkyTV/WioHb1ro7mT1stDt+r6qbdjNKFMk8Y
p70EPfeG7T+Ne7MLijlOkHcz7j9ZEL6WKS9pqtB6BBedkr67UX94N0wBt0lNmUAQqwa/Ck6suSmz
iC0AnTgqMtLCxYySal91BXL1XjDjIBQbrf7q90QRND92dmiSOKpnyFbibNrPT++xRNJwJA2bHWJm
6h76IG6lIdSYKgoNrILd8WDyGdppppq3+Sa/IZqbqQVoQjU6gqXLzQO0VsTVBpAIqGUxHnZMHzcs
yd3CtTA3le+ILKZpUWP/jhtLqcPgEBTidE76F0wT5Pk+xtZJH3XRA8vS4qe5auY05mar3Jq/DSWZ
rdJsZKvW9ZAV8c7tHtLfYCZ+nLbgGDIdW3fpWBSKxwaBqRxAYedOhUPU2c2sQ7sDJNb89NY54C9F
SWM9sWZN7ot8wa8p9V2cIczrsSvJ4VrSxKK7uEIcxWUYkv45RO/41ii4UcNczjJK0ABN2kWhckRh
/BVeTnl5baNy+tBzzzjmCEkBFFE61T2Zaf/mhrKe74iN/bdSxPYx4uyE6KqoSKEtSKZ7CNfLzqZE
ZWsHauH2y6TIGmajmc978g41Bg8f8UDIjvDuaR2TrXPCRPM2FR9qdBPQjj3KR5eXJigX3ELJBqmj
WvcQZX2xKdfx+ZgFOKx2EU3wfGXADGrkkw2Gh3wbSeGr8WLM39JYKizIRVdidP/lsV+44vRF/KiP
keFs2py6Cwc4nXnj+v+caJa+UiijadNiLFoyedWR3FDxgWLEF904ubZqTzlJ5GxjrsfN6gCnwLDh
+/KuolDtEm3uJ8weB9hA2zq7AuLzUxBvQfjTs4O7N9rmuu3GBDtP9lS9fR1HjE6ydKWDp38AOpui
g9KkjSjg4GktYv/iUp0HHTplPM/rRMVrxuUxXP2Gzaoc3PJVj+rC85M/XX6A1wiGyFJB7UMljcfW
u9P0O9kWICt1MNTJ5P1E9CYci6DxrjOCfd7kbXT1E4A4WXLTc+8sF0covOYJqsaFrK9v5UNjg7va
KudJ2X/pJIwhEL0nSoBkn0upmJstpFmqWgYMmPDAztYb5WtLFaIrelqV977aJpvX2f8PtBqHDdT9
7srwgk1dAVQuRtdQ0PMkF0Bjvv5JPU6ezYQdyEdDUuu+s03Ao6BeIZAkKZ0QxHlef8O3xeCr3O7M
nO4KWzo/C8H1esYCu+obH15j18RbgqGZinIu6ZA88wED6c8xrFvbn/mZaBDmAeKV5G6y/7lk8lAH
xPuB4ZIgrFNq63UGFJ8VIhmM+efpFRSJ46Bpe3FO10yyLSwpKQEn4u84ysZY2phX6eY8M/OSt+IG
vZ5dPx9ajAozjhMrm+40rqnG4o1jw2ANrJT1GA9D/1eNC+Ys++FbtM0HzPk12BwdOt2dUrU4eJmf
11CmL1g0G4FwGx8D4k5KZqE9B4Py0IRUi2i57jPeLYSmMjILW7rsY5R04L2si7s75W6nMD7J/Opv
GeeQymD36g9mLGZJqlbVxuws9Otn8Y/lzP2AMWfH1BoH5nAcuR4Yzs73WJ299eIBHSeofP2DJWWd
AJ51ENBku9synIN6svAQbFVg48o2rswZ8szfD+ZgJwnWg2iiM9mzqsK4EMTkCQmcLuL8t9B3YjTv
1d82Z+k1LVgVOartnSBVUooXuksBsCDAbpFdW+ASUZ8hSUTmLsdG78S1lVjD93vgTkHsnDLeY42g
LAIgeZrIlYErbWntCHTUFMthXKib7WnRChUnaTZEx7rvOxsN7GzYnqsYCSQggYiBlwS6CAIwoU/j
McaV693UYMYSWqw2gX7UCUVQWA99kLWCSMu9vxsAwelxO92NR0DiEy9Zu4noPP5Z/L2lo/IWIjcG
qgQDvlhfykdyXDA/RoMnbfbwRf3iBT/W6kM3x9uc5KMsmgTCYSHOo2Zwov82Leiz1Pc8BaWmV3EH
OpQK/3SuAmtJsCJcjwsucYi00C+PUexbmx9GHqC+iBO6s+zs9XshYUBrs9c4i3VNigyodlrB/x7H
GXbhPbkyMfwNnjA9VITDskw3uXtaAY0g3uWUWK6S71eMpk2QlRmM/1jzyi7yFCAzQsfxDrdx2SH6
JCjpR0NO6OarKKUsC/uvX8rXrSRjIx+U+wyZ3LGcstQkTngJtcIt9UQYQAzkLCgCHj5qdvNtV+Gg
YfBa9JPNmEzKmgOLRCHZVSN91IdeCIQInd49vt0Ofa2TjhpPoSlIx02XsbPz4oG6VyD0BLQczrwR
VE3KM1a0DcDC38MO53gytfaTauyg4bjxvU/6rx4PCmD/dLA/zrfDYtAyKgtPvv/NqDUC3VXLvP+l
GKYrA2fUsZIiJFElxV543++FkecI7vUG07gNHe/RmPr7hJufoaVcl4mcqqqkZESdOZjSDuiWBJb9
fe11tDavrAemhombMp5ZaoB7+RqyPdfOLtfhRqHL3G9qi2Xljrekrf4HjQOHQPxoMb76qESp+7cw
vOL5/eWgFehd+u8Hy10vGURVOUhdCF1sxemP400WNDdE6vWnO7TBauIUwGR2XeP1ueXHUajfM/pf
qV39I3DQjaF6JguOUMKZAV8rlThazGuw8qQx5BTyEnx9mwZBkIk7nsTuZDzOmk6VOu30LXl5ip7q
wSvmQqdiAg9LhJ3VVnuwZQURPl7MSQNPSfJgYMdhZgp9U49zdVKrUUaE0ummUMhlpER1W7x2l0XL
Ox7CWYD6DQlNQHMgMXQVpAL4QGCzkF4Ll8zaRUbx7DGVWM4BI453TvQBQXN4AOUxAKkrXBfBBi2m
jbXI+cWp3PO7OX/IQfsE7FbMGCbl0hhAMFqcgFrejV+oKtbRUquVNXWaqSmHloZ94Dhz6dt8uMYA
GGGCeZjuJZyVVwsRtoiSwEnwfi/qWupYppGeqZp5MM4SD86EujUUT/SgfAUJsERwpaoK0xWMyoRb
X0KecH00Ga265Wg3mZhWDsIGBioPSwyPkuWcBa8mQLjCLbhdo02IM5ufKo5YgxW7HXV05ZgzkdMz
aLJ2Ho/39Rwtl/AL5vVp8rXoVj3p1IxoHI9PFKSbYESq1jQnATrSR1Zw0mNPymnk4CBVcEnfrl+p
iMXmw3lsmFi2CWjkvYk6pBdr816y5Rk42aAJiI/SF7+78Ql4nF5YoflHNRXhjYU/KgK6drweE47Q
uwmtwGtbi6/a3YdFYG+RQdDXh/+HojN4boXIIbpNNevLpZWR8Sgk1eXbQ36f18s4Rto36NOdfbZm
FX+kC8r+XTZiKBSFv1wRg+jbGV+CndEKivP1EO0iH9KbC6OMLpnUbABN7Lu4D5hBhtCroNXjrUkZ
GwEtfVoFToRaCQFz2KpVVT9hDkB+BrAbXhTOC8fraCosiR0+t3hvkaZHdxVvkPbRWQ/nq/ps1huz
M1xYkqYSm1HMysWhnHMyhSVsEFGN6sNTGzlBYv4mB5koCNKq06aclWR89/lfUfvnFmmt5JEUPLZU
o6XQ+PGBkUzvc9dR8TjvccFAUPSz5e0BFPzhnsIIrlGJ7GXADeLG96yPUwgm2vtSKp9sO2sCT0UP
tiDqIN1o2VbHyKHOGkC6dBV2Sh0T82qT/wbq5zCvdwhbh6Ra00wJ5swzka2P+3ugULjl3gM7SRnq
2EZT9QT48nH2pnLXO3L3BC0lI03jcKLXFrEBUS9Pb3Q/N3/HBaDGVFu0k9QgfF/hCl7rxN1wmFsS
kYTa2VZgHPh3+MO+qHlDXqfFN1GkSHFF3Mewj2rHk3LLHyfe/5f33IQskvla8sWzNq/I5XFGP8SZ
V8lC1CRljOmRoDP65S2xAX9fONKYqfQ9l94atZtWVTGyBdtIK4WR91oASAnmWZtUpo1rA4acxzyn
fmKsHV+7KUjj9nFYN9ny+Oafa/JTiS5FHH/GQphnd/opmuNZwSEdo024qG92QnUR29nuKoCZqioJ
iRjUMQndZy7Ij489mGg4xUBBpsR8QxenM3OZr2nCfY3sd6VJSPkXh0rMX5lf/pr0RYd6x8MvtHuo
nPVg9xfdFink2HmYEkvT0wgHvIDiKWG2idDJ17l6l9zfN/CZd2jjyXJF52Au8rb5iMU6Bkwd4HPH
haCkfuIV/tj0wlz/Hc2BXyZkjscfkRrqJgl26AXLpZQgTTnjBgazEjHcbd4EuTjZcibhTqTY5xJW
CuqhNBH6wNOGSxyldzoAM+IpEOcJyxO37IxuUVLIcLZMo/rBJCW1GX9+w0pK9I1HqB0fxtvudtmP
2+p5AevhFnMgeIu37QeCbBpThXiytnirTOgE5/6lgyhaVtsEAKTiI4ODj24Y9J5JadyI9x4CPVWO
/aUfjNRrQH/ZQEWj84HKtup5HWoObDteSKWPoDlrJvoVMca4VaVtsHjs7dWi56VbKuiPW4kGQsHV
X0eguM4P4ne95ijvCZRFS5CNJ3fxTVyp6G7Yk9/kVYWYolZ2UEOAYKc3sf4P285V63pZNX+AhAgG
67vU7aIMT6Op2KUHnhdxoAx03ELSRQNzkXneo8K8A1s6JERRy91rm4MpJ+DX/nD4+mFbrWqhxrg/
bNuU1ogL+NTdTx5avgq6QBgxyA7kVxj4WuJicl6YQ2h+M1y9qgIOS+BP1Tul8dIOLbhf0werHQpS
OQEBuk1RmqO2fsTO9ZB9TPzv/VT8ZHgPR6W31I5rUDSrvUcSjcRMPmac7sRR/gocUxokcMVzZEUN
KxutjbphWjD2JrVu4kuaeOXCCuKUSyfnSuQ9D76RPsdAWE32Ma89r16WvssprkSE54geuJoAkrqo
fesU8p941GnAa92ecqWcHgP/GGnPigbiLJz3sICTzs8oHHJdymdGaDPRekm/1lwXPOncLSIpnlNY
Pvox7UXkJDJKTXT6wIIM1dbHTOKQC4BOPvNpZWqQUb1dNdwJb+DxDL0MrRMGS3Nvy/M7aieFHcT1
tJWw6vaj/kGrvswrpkarcEHMb7x6+CKY/jed+RQ5fhLkxVNqHDKe2FFk4S/67WghUmm08/UPBFJh
xaNdXJgqDQit38SRID0NcHY1tQFQ0PNHUgDWOKt6Y/jnSOJaE73ea+c5IEAKbH0ESsrfqmhg2mNd
FZfdQd+zoksr3Sh+UtOrmCNuH2tj8vvPvAfL4h3t+eKU17GTPRrOsaZFBbk2GfQ/af/g693schYc
zzKyo+5ndKf/7ue16F5JAFiyPpy3N5TTy7+DWFxmZwNAzvQM6z5ixVvtWdmM4plL5yREOkoRp6QW
y5y+hC2RVCqDwsvMOULWoI7r6CMNATY/vSf5SHgSPN+1bek2I2WEDExodtMrQkdypxD9NdroWAkg
mMEvD+dhVYerdYUzymdsPcutAP//Pv4qUdrzN3x9Q/E0GztFOUFa66NbKoWfBkVSldD5+On0oVR3
YHIHjenTSqknDp1AhYOhhIIqXDJ6zx2CjqZWkjIxcV7EKnocz5/wtIa1ErXMSPMglLAY65MED7MB
0u8b0UP/CIW2mTQGgj6sem8DdnldYxc90Z+/e/4QocP5VJEujN5EGUbtWv1wIFZ3jzFi9jOEBhg8
99b7l+9vFL3Si+nt3Yl5Idak7YrEo4cSUD54ZpLL3xvsowB/abyJAlVLeTYqvRvB4SH16TVBamaE
unNBuZhuMwPy2h9b/R9tUFTB28z12iYJJCwR0IJNx7SxnAemyPZOjS6umuXnSv5PiqxjicWRBBik
A0bh1cigeCwA6JoI13ME1+/plkmAjwCHkaeCIF+b1kaQVrx0XydsQYllh4lO3fUNZ4nCXihWQm1N
0E9nEYlMw3qgV939MgfYf2hQrdDtEEtbkUof40BgOZtGtZuIFFlBXVyai1a7wJZ+yGgChAbQmhxY
wfHml+M6MS7CMGQdVFNBegJdRwLWnPkVAxFSLekrlEOBDVB/7fkG0z93QxYKNtY025PZMzx8mu6g
nhAz7G6Ak0RXBeW6tJhQXo4eZiJE9XohOigjC78XRM4dM1wjJuOOiu++OlOjUB192XwgMUgiWkEx
gFEA2yQbFG1apv11kSbMUYwwbSqwq/qMC3zG3TBnBfpirkDZJMGe5i/6oauR7pwL+Cvlec5MoSfB
hsMkMV5r2PEkbdguFKyrSpg8hDZa7XkXF2nnd4ZXxCF5k6kn9jhVm1ur9JtNQJh8m6OkTFcgXLCe
YhrC04WykhPFG2Vzs5CnLJEDYlXEq3Wy6GsrFN3WhGrojzKbpUzXfJbAV3mMWaqDcQ+Yb1JnyrZa
0bvnzRzC6Zgn1Ulvthj8TZORebugRSNk3/tG8TGqTQ6+nxyTwrvJA+0QqBuhOE0q/nz8avoj1GkY
3xYH3rllfjq35kKjZ09kJtxbByUGbrcBsR+n15uUvENppV2zEgcq7cV+Mj238RjfjvyWpfVfHX8l
ZNOuIvCc1EshfQI2SrGdy2mxsxfOF46U2WaHmj8ACx9f1ODrlyIId313O5NkmE2kwX4QAD6eAEyw
QovqbYl3gSVQDwVW0OlvEoJV17ymImpUxt5ghbUAraRifVfw8Stpo5KcA5IAdrJg49c7sicRRmIR
3k4hyOt3/6MME8bfXRTgB8lIgkMycsgX8VG6yI4kz3yLJnyTZ3O12wgkYMuj9/AQ2WHTci1UByHc
7lzNzhdtL1++jKIZsJfGI9jZJDQuGoKClVPKh/7ip/FAdj9bXcVJ9ufhgMMA7hf5P4PrNK4vIeRw
Kf/9hR94ryYnJRpmq01wQ3+HIaupvMpa+nivOl7vmKRtIIsPmqjOSHX+bxaCxRAl3kQPklLysYXa
KKLz8LdPfQgJQqwBjAos0Z9BZVArwch9jdFirEQHxII7E0XxaRpMSwSfoUvd6AhfCa6cMS/2O/E4
d2i4/Tqv6RCZ39Q2MZFYyuW04lamrlGxXRsfZ7ryK4lbUF8ZH4I98uk6VxX4nxdCWc7GE0kMx2Hx
iTDq1QMD6kGDgdLyF5z3yAKdn0Y5t1IZuToyMPsJrDEFU6Rk5PC4tAKhejsG6CJAb1jpZFEKsNJi
1FFT7RJ94BpLmvKXpub6QP3xXmlNsiONDmD9wvuxvSNC9yAGobYks1zHkDBq/3ijB6xMxQZPNNaD
fa1Sa8yYQuAgQOqwDdhgmt9lMsd2n7wpsRGuwzKYeHYBskQhjPhILrLYEjD0NwlSi0L/TRBV/qmi
VVWGDYCpYRQQXVfpkI7ugburH8DfHjqt1h5rKmCuzU8uOoDk9FPHgIqf6b19WO/jaZYkIb8tmnZi
4RjRArToidls7iE6QrddkNHtFpsiUXha08DpfLfA/g/SE0vsym0wcKY7RlSi0NPdw5qNcxmBfLEJ
sSfHHyD24RYJ0pOuh5rTeQN/2ohNqUmGeNBmavlYkGxt4+DPMmA0sBsaGEMsVqDm5xXfuNU1RSKq
+KgWMOQnGaEVV0qfPOEiTclVeum8bnP8JKUeHcqxnSQ1v+NUl0MTzvU5uv9+PQJRO7I813Bz/Ud0
ItkGo4FDxaJ4VbfWXOmKrSKvCPou0g18Ld2eNl3/OKX3+5+crpUsFWrhy02YqAGIrrOXdinABX21
+JDuLwuPXVu6othmomsmp0Bme4CbxRxbfJjl4ZWQOvzJPRNGNDzMs8YRUchlJWdISE+a3InF9ny5
YEi6POM9Dj20hYDWVymJRZouqKldtNOQaQzcFfp2d1jt7aB4mdjHBgJZ9Ccl0C0qfXZVr4Cb/3ML
zkpKeFUYNGhQPnL4SIdg/hIqm4iDeK5TBdURLqmvEAfl+brJ3VvFxBwiEDqk49Y+Im8bUy4k7zb4
BSdcXIKOju56fbNrQxFOfQ5gFl3Xb9K6pJn0jLz7kSsvhHWve1bLFyXb4JCTQDaDm97qHr4d/7ni
0dFfqihoe6aGVU0nvsQ6njScUuITWfYQxSfuvxk/uEi8UYUar161goRoin/yeXHYog1LsvGnbj3N
S5w5J1k5fwfXeb9BXwoeCNrApS2Qey3vUCUDPu2ka0Y6ckRoOvPYkUwpUPvtyTX0FrNI9im2hHBJ
O+4dqrVkXjSGA9E+O/Ip71AxqeVIVAHs0Wnjk2P7kI7XondWV9TIIMagcePdn1kQCC+Y4Ge0HZwr
EESAaqQY4ENKrMQeA3nkR3C13DuuyUt6cKjmNU08XiEh9I/LNybaIkyQ98cMy0+AidG7kgSvzETk
uZvzs41qxv0wNsc2P9ZdfnAsdaSijs7wKfSmMAHjO9YxG+BuEru4d8ek/ABQg8ylH90sXpv55HxX
J92x9LWX1aIGuCocV3OXYUddhitxnDhA5Ay5l+bhDq4mgfY4f8gK8pj6mdsYVQ4vziFTYG+baywM
rk4lys2nbErPVkgCKga4rlywM9s0qczLMJu+WwgyGfm42ke0qKveRg0yv+E81Tcr3eKqb9k0KDrk
H8FZ6yY6RtaK6m8MQnlkjhDe2MBidUr1IklrY1GbzIBfgDVfE+/7lQwqaSJCwzZYNcOGQ/bMQWm9
NhakX9HFWcCf47/+FdHcJmuIRJDdA9Ph92qFFW6WjjSGuHXwWStXIw81u59DIEqURnkxkuW4ghaV
GLEVXE2u4mjZl4+EwEtp2Rn2QsGnhwYPKqyHYgTOqilbG2Cbqzga1C6cQW4rNTKG6TopkftInEyo
ITO8PQAKuztYWuYeckO3eSSPj+V4NrbSUrKgzxbP0ctoL96tsDaPLAzJ6olqyPHBpD526KSSPU0w
Ozy6zLnGPCor91pjnlwyIjcwOfhw8lGRLRXg11irqQphDW4yHCz5undFgD3KzwJxR9OfBBFxntEm
5Wjal6S7YM2EQm8NiltVE3PSq+fixn9GJND7gg5m80BuS7rhaf21wC/4fD95jRvH7u3Ola/+9Xsk
dUzKmEQA51wQLZfFSVnPzdSEnBxAHyLEfsyVJDCN0AfX+m2U9zveiHxOU0R2FD7h/BjMJkIOjrxn
4x8t7Wh3X1BIAWaBvZAFOlGHfF3IPG5ARo1P/+pXXaB3N1d8INbZVpiUESArwset0HgxiK0w69fZ
ifmx0rSUgM51f5+xrH4CN96XuYSsKST6+jT1Zpv4TTzizVIbJ1O81SY1t2ZDRy+feCgmAeQkcdl+
H6ebrn8zU2R3IvU6xb5y/fryzY3D1Wkg67rVt5N3J/6ciTNSik4chYTfuJRSafshd7VBcU8y4rfg
BWi2TDB1OOvfiA3g/iYVwEwnrfwTCxKduG9FVkcc9cwd9+Bh4RTd3GaGH/WwLgfCW3ZFJRKkx6u6
7mkeII4EDTYTyl5GhEX+Nef8m9uCfmbmfPpLU5kLvA7AnY/xSDtGP5osAc3CavQf0h3JVFYRkNdW
4LTHv6lTl+jUc0i4Hx9Xa5pEAi8/7SasZ5FETJojRw648wQ1tkOnaxCmZU7khJrBMCio44QOfabs
WdxXfYkLUO7pYLvIx+ywpFKkHMNDEUBxBi6zSzizKhLPylCxF59f605qlT4P3P87O9S9z7zEz0yT
tcIWEoiZZWu5VHGKMbq9YSSSFro6Sx9UypLZx0Eu76WmjyGjJbIoi3q/r9ClSKpGQqdOLFu/pvxK
OFZKeIEGwqt7Xatzaij41Ww8jGKkuhVxW13cdjfgGL9oj8sdrNmlrxC9jw/w1U1U/DT8jpHSctEO
5aRDXyx5knekKas3O74g9PkvCqO2kO+891tJgEM6rdHxj9zPZ27SNRo8yCNjhG4/Ow9j3Irnk+Xx
3L7dBsg9tQyV4Jyrov2JxyTwO/mCRpQ/cDkdxGPilhTaU8wOiB945dLG3EzRzKJZfZyc476RL93Q
dj2++bEk5WHO366drfiM74NcJTyBnjiDN0KiZiZqmpOjBsTLQeb9ZpmZq0KRtn0AZm3mSsDbris0
HqxqFvgu6XELCVxOsJLSD00hALq7BZU1/TLCxzN9iENHpES6y26lMhBRDpJyni9/8aZdWN9pXEV8
i84TLTBECKsBkA6w6hqE9UCZuiLXvrZNzVRanM8VSOnxt1D8mmoB/qOeoQWuCYP0yiKb3lEizu2u
ZUZdxgXvtoD5/YompV1K7ZTymLbZxmor27VeChNxUFQXfX7EvU6p5aiMRKXw03g+/DiGVYIZSiGs
vBm+TDuGqRn50x0HcIhcFfXRznItf3rYBUngq/OKAcawum13H7RvNQ1gJ+XMhwGubjtbCyWy9GjG
5TPHcMp6LiSyP3UJopAkJ6hdmb8XHWjUeIEQDtJVBgJKKgW89CoirWWfYvvqiwGNmzPE6UyASQuM
HzcJYYZPeXMQtMh8VoTJzlOeRjlY6TAgdRVZFVZKF1dUQijI4UmoFojyryW5o+KevvQ0PbhYd0vY
ulgh5cIs+wdtjwXuwKXsFrCAMkaTg8Xt621YPl+q/PqOUjmoXAbS5sKnonh0oVBTE0GwOsOoB7BY
ENiiJbDbV8sEJuiqSWOeGVFKtyxdmm03TEniJWQ9oOQUjmcl7jd6n3hJf+5xDD0bd4+b3hJ0p08V
zL2G1/RGLHCb56nMZrnMPAJukMoQPahJ2yCc9sHKob10JH5NdIR3wmVIGFPaxhRwqHZWsftTgMnW
P6OgxjAlqDT0qZIlpK+7d269lkBcE4lMyQXkOcZfGr1ycPZElrUVtC+dMrfkOV+OaqnORHdq6SL9
GfEAJRJEo+DsPZZYHeZuhbZ2dngoNogj3WBQnja/+Bcv9P89cCsrqOVW0eC0xLfFBgCkEwhs0X3G
gc+Bt+pvuFJ2JgdiEqgZPyXvEDGm/krCbCei238OZLP4/6Xr4Wy+vKqJgbLgar2iTRKob1vPIAhJ
udiRbgUryhHqaAB9tPVj8ZFeBZGGJA3BZkOqwS2PlcwkIoT5jKKKgCnaKUpQXRWJV7Xkvz+gVX8S
1WMgL63LrDu8Kq3RSm3P0+yTXYu6fX7kJGQLfl52qVnKix04jPLq2TkkZFVJpXoV1hZINvtPOg+V
u/QAgAr354VHDt+oe2pVlFl82DmCoMh0mkRl+6dSAxA42jtTFrx4QfX9mVuKY4lkiXVQf59BUcSM
4gNJB1KX+MxD6cyS+hi2ouAYuW+Y/ENVMB1RdKGcnoSjlzz46oqDiNQ7wPuiuNaP7D2oZGgJEptn
+27z2eZ8XXO3yqAnyycKux6gugUBeMoWk53J/ztU7Jraj+azYvqJHB29Yt+QGspeydl0g0L6OiVO
Fa+kCfc3jHeQoIG7GiT3nelpEdH2Ea3s99chSGAwehaLWj6fDavPT1IgbFeq2cVCGaSx9ZaoJx5N
nq9JAVYhC4L+NvaSbMkCMQkl5LeORicGTwx0d6TYTB23MTtngibgie6/4m590LebxTDF32E1t2KK
xlnKpGxysXvfud6ILhKy8w732PyF+kFYkfWOT861u4EZPd+EZG7MNGIZGG1zolVY40dpxp5ms3uK
+sCxu2vRMbhDUNbj7RpuAnSiqAEgMnNcRzy1jMu/S6w09PHuAii1MqR1XIVBs8+T0wqO8GPZ3Ioe
xI4CUzzQDAzBbvCG66i4N7xQiwdp8+KB2hYcZAb+6WuFqbbHKFwbo4wGE7qZ0Aw0PmUsZeNmLZVV
7D9jq1qCuC1sFYi9DHruj4bM+68UmfAdbcn7hgWl/lrcOjDWjZUukLDZvC8jDBPQ8+s/f5t3+M0z
0x12Yme7GczZwH3l66jfSgwJYe0NbPGW63x3t2TJUjGCd6Yi7IDlQ7s3H3mW7NAocmGTqHriA8t7
LDBRk3LE0fUpCujLjb+rNgszNF4ybIkJ/TOAmy4dm0Zkcdb3PQB/uOiwKVQTbRhV7Ukd/vkw5fn5
29PuPh5JN/X+fyY6JQaqMFtvVB/HVGl1rhBrjwRf6yCZ1j492jYTrHH0ifOTOZ63cxF9MdwoDeER
jfSVg2sGly5IoqYXeGm5GhybafSh5ynyLIbGC2vFZfMdeC6qSMblR6wj/W3z8orSisDPwwzeJOAd
Np6q4yYG8AnudIfg+AuuaOSmNyposQosDXEFmMs/4SM7LjX6xudR7IF2wx/HkB7TSJfFp++HfBqP
us6xdIjChRlfMLeK12ZFmJWwWU/vL4lnWZoijX8RPRp47Q24BtUyBA4DfnEpGvCNraxZ1i8fJloG
SmFps36ZJoI+Tk1mRAVYfw6txcKRFXWgA14ivfXOd7J3MAetKbJhZ3ySve1r9i4yUryh1SmmrCa4
pnkLyOj385Ew4E9Wf2UqPOwCn1gIWurRZPYCo/QXyyDwnaIdVos8tBW97lkTyp/MRbS4/idkNr+6
0N2eLDTegIi/pMeeAwtpxf8VoFM0JVuzt2u+J6kkQQMWYBsx3Yfg7VQP2b03QDh8egRdMcqUK4Y7
I8XtJS5g9udKj7J2ebpabbbewSHZ9A4OUjCxz6MoxamnSZjrsK9cRLRWoFdxoMR53SSKTSKLj+cA
gTvhyihYY8Mj9jGZCWUTFKPU8g6xe5quogw3j6x/4k3OZf5agI0WfkVRGKyn11pJumzNnrnC1wGg
janCKCIinduluEomFwJtV7CxcLyiLHvm5v4o0XRrA9XR6WaxNa5UKERG9uR/uQR37e3QpISjK23W
gkJxpj03BbX7I5U/gpGty56riqpeKkMR+2TBh2t7cHPZ0pCmMATiN+eTlbnnbE/nWtXuXBTkY655
v2JlxH142Va5jZsMyJ4Nx6E8u9TZ/L2m4acG5BcLmZTpblLMr6HP92BI+fn2IN8h65j3b61UDp31
UlEtQpEqC8/A53yNWlxBUyBMj6m7Y2u8ZLeltLHXUFcWDmxiQtu0+93/cgVghd59qKrCXOTaMg8K
7eFD4UELhqVk945MWgsR3qi+NNcRLWjZqHRSmsUfRS+h3BmqczpfQFSvg+P9n0TtJ1UM/oA0kBxG
BWKlMxLPUVmlByL4NA+R2YZ/reBqMjroIxydDIrCF1khrO6BAUEDYCJNyrgij3yWDMhKdzVK7e9i
qymfSZ1rpbDH2zTwKfqBhSUVq2qN42+Gt7fA/iAIlN/1dJjLLarcWfE92Z+/nBdXBDsxD6IRYBeQ
6+ldCeXul0jiIapq41gspAqvxdY28ZWIgCFtXUzWyJ/akXz0fSrYQWqpIRR4P2oekbtw/44mzE3p
K63lKsHzwS9nzzdEw0rHSz3JY2VpBPxoj7N4whl3IsfDg/+4dRgS6kvH72uhL50sBxm5QkRbQec6
rIj4zOko1mn2BX73mK6SEfytjX1+XTQSj1pP78sP6pXzND6kct7TLy7KUlTWHeRGHns4ZYhIZT2S
AxUfTFILU72cfgUn/0cU05Awr9il86ifljXH8UVs/dBfNcwPA/2YjDqOZdzP3CP69DCUk466sFNk
htY8bktWMAEM4VnGOH09POTeSX7ZhyHvSLXFtIRp7BBVgF2fz2YtHIQ2P/BVnD0evebvXIm9R2KM
s+rlr4ARki6sfuUwlIEQ3JMD/1OOaIAy6m5d0H71N/GX4Mi2fAqaxbpnrso/ljyIp3iCnTwUYM4D
fpojtjtTEJ89ZY8pDviBO6BtePdFrQxpsAm0MhGclfLs0+EG0XZwFjVCNiCYrcEyJVd5ccWta6ON
FewqbjQ0HcJ4day25JxLC8SApHkPDMXUBjblJveq7cMwzxLWCsUwKHfVRU8uGElztoVKWGTWtX7v
KtNE6AER+ihiRcRJK5Jt5mhkjSYjJlRy+fLKhiIXUqqlotnxKUPxIG/+f1qCv8NyDEZT5HzEEZzG
CT1d2/HAcXaINEvQ7HTMaEXJVGNjwi7CtZd6aV+YZX/im4e/k6RREGfAPTuYPXwRNAR7nHCw3Rfp
AYUzYaqPL3ZgztAOKHyBQkOKP2DoPttmE67gjNDc8Lb81SFvmdeQaT/EC3Z1wB6JeetBOlrkOFvL
PV+m/+SvBABFunaZbvR6xI42R7jD9BCJ6l6Piu4znixnsUhw+GsqfFx5wIQppYCz6jkMKvd3OtFE
OxDLzHV/BKvhDJVtB4u7m6tnWa5ashZnWMD1JxMv9mwitp1A3bXYFWshGauR+R6j1koKTVofoCx0
xS7zW7SUDdA47nuCsxN/lVn1xFde07d59ldTcO5HzdK8wBrgdzGOQ10feHIVIRTbLYWLTCb0YFQB
jqabuvbZkjNWvk+Svh7r28WwC3c6Q6v9PHAZgn0PIi69+K745pBQi7Lx1d9/ynJspafEu6v8sWbG
HqCy8MtHiGmOdFVMVoTNkQWzJzqOT1JEnS+TkeUf6BvQJ6Inu1JURTh2bvo1wnvEdRpfY44EUtP8
pVtfwJEKxSFM0D5GtAG6vctTOxoQ8IWuK6Bus6rtG3vT26428EuaenZEZ8weq/VWnXhV6AcC2ctv
tsW7DATMizAKUtj9NRQiEJJIE04Au45YZXrOCEAP41oLHN2kbyE6zje47zmzl0kUky8JzTaiVlVG
+AtOjf3ttToiditBFUdGzWnRqgj33zf9Hzaoj9nHo7xUxHj3eMvqpGTH7o8GcdlbPuSyuqRcwC2Z
iuYkFqOSrBBbyJfZUBfhXCCVmQtdSQwQYcA3+GTc83e6MkyFqmTne2Ngt4F9gj1Q4+30pWBgqgYL
rzTPJ48Zq3cg5tv4Fu5P/rC04raaeWTTUZwvmcD3AYH3sbGaouysf4+GIIzjB2W2KWAesJr3CVq/
ii8SqtAyV3N2vx1J9D1j3RSoQI4+9YxrpZmuWXZAqGSy6alHg68Npw1PS0BKg0w6S9XgmzXrz5xf
O+pXa6GRdKYFyU5W4n6Mjxtb7lyHlW/fvu25fdq/h2sa6rul0d17rkpQ2G8D6nkgVBDPAOBrqwk1
tH2rIXEjdHUXhu7gQKqEIHur3cSDPHZYWr/rQXFLDzGOMU0QYM3RaKIblike9aCQFY8ecQhyYXu0
LQVp5q3QZAjgZ/V+hG3FTlrRSeQHpfvPViSd2ph/bWLdBoGVDcPTG5cCZ+S5RslIcDB4kAD6jUf9
iIVPsenjqyeV645vQpRMmC/ssXWACxSGyczzS8t6YmZb2RJiGzXd1luB8LGlwm1BCtmXhN5drmiX
hu9QpYv4QT/div/QeYIgX0gVpKsquFzoRJdwBMjjwpLZCkgPocJO79GUYwGd5Y98EePqytnY6os5
wMPJPWj5UVUyTB7OQ4+Ch731Gja897ZBbPDduuXKPmqKqrOFCLZOOe1LytnJtTq9+I/Xacy+s+rb
vfIlXkKe8gj8tnuxqyL4dxlykeafJsuX+lGvqrdNQdz6ZP/sRCkSquOeaFbQl7MC13u1TCJctDN8
iotJcz04Fr4Aw6cX4JSYith9pdUn9coVzEg4zCYqtG0UQvoSwiSqEP6BKzz3xlQSkXHudw9TixFx
BgpWh9zmqmvmJFWXF0Yg2pHVTga8ImJAW7c9dKCO+yzxo5EQ2gQzwKrgfyqfBcj0sQ2C2VzlNfQL
BoyUktWpZzfUV9k6Mf1IiVmMDVCoWvc9RNnE229CHMwK8qeZS1Jv5UOUCI6kZ0Ggp+eLuMKCYTAC
lwVRTfewpTGdn3a8RZ/m6xKC0btfLRzfH5xj7DYuUcYnedyn2VPrUEIM4uJqaUJmQSsKQwW8IDL9
o+HX7N26+gRz/p52DrxivV/ro5mwkxERM2zGb1icfWLPF32M5aZRB9Ca9G009tYT09dUNNSFiZsP
9yQJckxyFFYdjWi17VvjrMX/3J7WSWldu36yg2riZ+lxrFb4EmZuMWNcL7l2j0TBoIPbOugZ0MTX
mOOoQZzHu69wfqZQ55xPzXsWT85gUGt+4OEEfGtgQHC8q1jYAsawPT+Ok1f8Vlpdo6vDJxB0+2sK
/xNmjvGYpAkNUuRgpfO6Tv8qPRLBy2Jkjv0U0gDaGcck4rYxVTzDj41xBM61hVhW60FZiKl2sY5K
VFg2rbWVbtppAYZHwpSBht3hlJLwavIrEYgmmrqReEtRt7MEMFNd7jAhQe4aTAr7ewRXxqEp056w
z17sLXV1fd+MJ0wYOrkP1pKNc5bxU+VoErwRkAqTAKSG7GAvLOdEh+isFs+q7ssKlKK/CJTXU/i6
4klmVdazIu0Y71KCW2BbZ5EJe5Lii+ft5ComewlYvmQMBhPMPpaXhVL33jE17ZySXnP/3Pb0+WzB
9LrdJSx8XSN/i2TGaV1mePelOx9Jri+eIXy1dN5c93cTbiMg8SrGWcxIeGTJ1dmgKZ11QUDk/5yz
FMZZbRHjScolL5x1Hs4rk5xFXe1+yttzOKwNQLYC7Ryp3M6x21GKOAhFqckOcHE8a/rTdlus51E7
b0CkPtbZg55OS94Dxdar9B+DQiTFbok1odwijsM+hI3i+ngrpuAg+RHxQXISVFnF0s0b4NJarbb9
YOV7xZJ/E4ZtJbZX11ehxOZi41J7+DfX9H1xwx+AowYApK+qxj0V3Ydl/5T864A/XhstdBG8SgOB
VBT8SIvOltBDwZtenKynWvvM6R5bNwYtKg0u2PMiWOKiVrldhrhSuJYVYAj1H79SclvZK6/vYCed
FQC7DufA0ebooY55n7Of5K7/mcIrM5A6w+BCiSY6+49Z0Snu3jHmLqJrk1mF19KjnsuQK3iqH0Pf
rOhRVBGInUirDAB7EGC6vM++TeuQRegBfKeIW/y4tBrgXEJZ+jH3U8i81pNXIk9ZDw11/nqMLPc0
JpoSx7ajF6wsw215wQpFAnG8vEwRSCB617PGrFAlEIWe0jO0ippuh2FWZPUH/76NEw5MYU8ic6gt
AiscG76EqrM2ca6rpJ2QOmwdtbfhzqdw5+BiYediFtvK1IFSf4IEW0pvcRy/M7Z5/iIqWzWXCSbc
C176463wfsYqvRTF3zf+ULlHvU38sWcQUU6Xu13I46rG33XhSXc7xUEZXj8FM94Cmz65o7MGOFbg
BX1QnlORUgggeUvuwBFqTgDR3xZMkUGrO1I9NrzJ4ol/JA4eCtgTJFF7NikknH+0aFbcr+6xTxKm
ooiUfmv1aXG6gtBfZhd3mUbnPAk7hhJ9fL6AS/j+PqPVuqkdKoze+OuNo6yzGzuqjgc4DiYGTSuG
R9r+WSIqOPT3g+Zf5KmgBm0MjUnr9rB9Y8u3/IEkJypjeZyCoyMXB2PO7XEGIAzTEcOqWJpa3iDD
M/cIX4R8Az821hpo/B1BMqYhhWOW+L9e+9cDctK8p8Bbdxk2YsPGEqADwtuJqjEtuWctQ77bjdWY
0+9bzAYb3zvrnzECo/uYHql3SM4KQbqyEpAhEGeeYEtn8i6UAbB7SkYCD1/9ewNsWSIKLfupXLOW
xv/3JuXbwc9926fU991fHAX4vwSRMMecUNmwwX2F7wKnoZTF9po+dNNBz7/rZYblhtao7MvCGOZH
bXrSvq+c8S7w88lw6AbtdcYRdYNLsnltRN8Bn4Z1XJTdao/Cj4IgaZMmmlyx7fjwJmG4pUxuPXff
LT14aVZGLb/Q5I9PPFTXWr9KCgDw04Du0sd1b7xm2W0x0vgzFI+TA2lOI2X830S5ByMg0gL12tp7
FXSI5PkxN3Z4Bf94gAcdTo7WS3oftl4GWWA0mpcUKAF1Vucx8GBw2LLMp5NY8VBW/4wtFcYdx8OP
RuwTmy/NXrr1memYh6OKhFY/vDmRt7wcIK9xlnjDIBeO+VBpG2GEWOh3KobGMmUjQ6y9HTNnPIrc
mMbysqyHyit8KEtS74LogPdE/DAkPef/+cnJ6vZIGoQ4eGvspl0J26AiaFwZOV15OCl9twkpwGyv
B6xXKwU33GxZqjt34zEIMiBsyOq2wFjKdWgn+OWX5XvD7xKnBmy1aUl/vlQ4slx0HiUX16hYOPs5
m3TIQ0+ei0rRvr7nWPjF7p1Se4L5e8TaA5F8iIWw2cG6Xo7oJLJI1BwNQMTaHzAzoKw5f2ATswMH
igHna1Q6HRM/97jI308nodKYcfrd8Ljluv9TmwBjFaIWrA+Ct68GPZWjBFH2cm72beLxOTw0X7Bi
WUVcXBjAad03YkMkQythidzV3S8gs5jIbxqakQI2m7yr9zilrRAKwmXenccdVdvTd2mfW6xykiVW
v5ksx5xnGW4b4poLd9i//+FBfLl2ff6S0vx0mdgVzllI8I82xCR2FepX7zXgWQshbaWXC46HNCTl
Z2Z4nvFtEyFoyvuH6NgBq1UHm2ZFpjmxkQbjSutBGEl8BG0sgP5reH4qysdncQLoKnaA24hsascN
fD0O/CpoAx7PkWY53Io8lgiYUOtX5J0sxghvV4DubTETY5eYgQjYDUCmme4isPwGDKiInx9/YFL5
lCkeiQ7NthHlHaioct1P+hGdx/6KSaI4djYNm84j0IUI9PgZqz8le5ZUTZJ9POGw7GudL3OEfVo7
GU5ZQwbOZzG//pjqaDe2DmMP5PFXCemvdYqeeddijCtexy7O6DNIggeAIaA+ilOLWUp17yCjkEl4
R9timiv+/lPmg3PzAMErnS9O91XC02T5DpTVizzkGKm+ne6wwkFOu+W0RtE+secTobWQqLDkwbcg
b5cdtfnzWacCgdi0gBr/uaWU5puy8oTDa4zddNmNv3pq8eHQHg90Yhh68wHvNYBpsbl/SLdhWQNg
vIqtvMyu2ReWsX7ZrGMsCHD29lUfkL2vyTi4wmSEzs23+qBmqvanSuLUiYQOlcMzZZrs0eMW6Loy
QIwiBvMI0jo8+VxEWvZcEU0kBc1kTWzOhrSJkQWBh4vVVykhnsr9xZHKo16qpPeZol1ufDFwWuRk
t2OgJy89tzYgMJiJvrELUk4LWT4EAeyaKg3dKDBfvQORfU/wBj4HlvK9HPtXJFWgy/FkMq9JGapj
KxSZDGXP1nfcpO83+emopl5/ibb00h/y5DAE1D2C8iYUMsAfH069ngsW6qyDzOVSlJpY8NMAw12p
+r+d3nyF8WXQ+GGjwoODaBG7ZgtQhgxsaWgMdSwtx08F9Fule8dhWmBJ+Lk38s0lJlUJdFr3mcOf
n3CtmnM7GU7OPKcxYvg/N9qo3P0kUj6oVi1rZsbGEvorFxtmivATq8kU/3srE4+I3xeZLSDUfjG6
vi8rEp9ZNRsPdrzySAKpSjRBdwfl5b32+qET3DcleTmAy94BEHrGogzjcsCYSjlwLozRVmrJoZy+
qLmm1x5jhHiBHMLylcQ+eyIKSgahMCLDSXoZy+1dpheDF7bW9la+Xe7g4YFhc0uvX1zITZwTF+4x
M3ooJ9Y2VDgSevUbOGrK9QUNA6sQYDl8u92PDlEVZ1mqbyd0NYwsOizDd7tXgoXHCRDB5La0V8gL
Bp6bXUHeqMK0tii5aEp/pdxfQ3Ha3ZScR1w5H3HqCF89o/IcVu8IaW0kEGy1jnCCaZCmXIn8sB0z
8WPhjbMJYi5w4K9zvjeL7inqwZhk5zbn3yHz2oYGeWpTmFZdJnEnwYXzYyItz8s0bP2xTWVNgMh5
VBpByXXPlaPoFsufjMD8yN1VrU2b3FwluNl+ANOB015v9n/FOLad6G0gEiVtetqX6ZOOfNNV4S1l
oulYn/mM6IOdOEmMgSB6RVxkzdLXQlLW9r0UvWKWDNiB3L3uJq9sMLl/mWnNhX/RIzrA5bwDn+a/
bajO1JKRgo2HSEtjOWbMhiuY+u2SCoRSl6VryGdmI6W4K8Bg4dfrcB2UPVqExztU06Qbty7CA8VS
uh9/Ia8RETixRZmVOcKWt66W+I2dPcvExcNfUkHeFABOKAABTl+e9Q10hf/LdLs8NQ4Kc85kwkEY
RjnXiMqLxHqaiEUcy+VMBz4HPazVGijbs/R+ZOWFlDl0jr1IDrl04MA2uOH3r4qwdB5GL4X78G/7
mTP0JG519zFCnLPVxSE+CXgokA3s1ht8blphW+fcv3ym+s8WlFHGo7rnsTbcj9TiMAfpWyukln5e
8yGIgQBQC/OFt/OhL4adHU+JXfuLDTStmtla1Jk98BnCoqcl+5Cs0LoMtH+xVz5QONhThUtzWEtC
4VT1dPAIdr3CDQhl6Boap16HM+cftRyjrFja16btwu2wkqAYqd3dFbIPPDaK/8D4Q6s3z1bqqhCx
PUaczUiIoS4AKsvDyA4nGy1+h/B3hlkwa1iJR5pGJ5k5a3QHLKZikbrNMe5wZ22uc1Yt3ozuGPiO
DsVqRBKY20fNblKixZUrv8+oDygn8kVmJmSMxnT+rp7M/yee7tLJbGEcPPBR3LxiVUFPCgFqxPWF
1Vvu+V9X3lQ2K/k8h1/xHc6jiOYep5t13YZp9LJDut4trJrrgWn1i+6EXbOOLQg9CGbWDlmz3bdJ
lOTGAJFXU7Wf1YVQUnIUPSH63kho0+e8bYskeKasNHMG0igjT3Eid9OmcVl5CMrryHwLdS1TPOFI
zV0SDpBbewkgeXp0gHRLhBk4PIAb16FlaL1fOPFY9Qf7M1rfej9HbIQiT+oEQBeXa3zmCnV3miTD
w1dAkGi1+lTMGCc2XWJy1NTHjA8vBnLKfplB8MOWaCEIxWh9EeR6zNqXjBn0wh1MSoP5VUvzNk/8
LzaIE2EozoasNxXbudGp0hDCTFNKhDEKLyP5PxQY9seokST28HYBw3qfvHcqwfimg+p0M0qSMdwN
wkg4loS9RUI3aKWnzOP5xSldULhutPzs6Updhh2AI0zNc4TJTqsCh+dHsmH6/DA3R9qDnhEYIxnc
Pb0xZY3ksfhhoeqIfLiTtSkiIwwhc81RmSCZe1CR7VWdkzyKpjbx8XanUppOEZhaOo3bg7zX6W31
eXaAw+J9cuVgP9keAjwlY4ACTumIKxrZJzFud1ZSH8sGseJB/MRhrLu3ei4Yw/zH2d0hMaNvmT18
J/ZuWJvwl12QzcFnMuwuGIA9LsP9ngBAFSqcM4TjibmHaTcVfwUSh3fmuyhCACi6EjAEDcayVnNv
5RaspYgSj7sF8ND7ddv0vFIJTb439bDA8CWvMAK1RzQ0UdKMYIOTeHMBomWCHUO2Iscai0l1zJ5p
58uq75DjVtOxeCzD5RSEvGEnrrNh5NfD30a4SshfIRKxg73/Dhrx71ZtxKdJE2tMGipXddIBZ+6R
Q2IPa//tEWVTAfWL9O/fPvoSTyvaTRYhvSgcl6oRzUlXQOOTnLIjqMad8CausxK1supPznSUcAFb
hlJayEgesv5EDa/KRVM+zHZKEgy1zNkZG1u/66BVlyfCebJYCjiotDz2Jue0OYbHAmlteRUUBxt6
vDZRoUYxjJymJWT5NAN4WKGJNqdqbKl0Z3rYVjJgX+EgmB9gIGbZ3v9IQomaH1is7R16dy5OcinD
Vqtl7jjaqWqAffs5CB5tx1n5gasRAjYahoaOsD9JihUI+QCeTelipxsc1AKWOMRYa53ZLTqDNMnr
Uth28MfRw8wp1F/ZkiJil8JZuHxZAmGHMwW1rIecJNZSwW8JS7pusLNg+yyfRsoOsrBl+XPTkzHX
PZyfVEo69ci5zNTOTCrGF6PZ8yQZr9eEOrvxqKDBsM8liP+KzPw+k+uN4l96rnb9USEyvdxh+2Tu
W4XBkYeKTNDdpuB+jN5GwKJKowNQXGA2Gfo9avDkQfp/XYJrN1g7+PS+hRAhUot8YILKtjysteOj
5FlWF8mnKk+NKURact0zvaek1fDxE5t+3TqNdZwl8D+tP44JUnijQtjdJZ9+gmBmFtqnhQCBqNns
9WN55gdP7yIqOE2zFA0zQOl4OI1qZU+lwIzBkLJuksWpDphu+zmTEuBMVyogjeS5haMw1EKdlCz5
7yXb70yKy4QYV9+qmiz/u+goOaHogMHmoekJNJFbZaYHwuXXBnA4tBeUWEOSJB3+objHpb0s8w46
E58N3jEDdc32lul2HKhpnI8UF73BEmqu4uvAHnIgQLGp8YEXA4So5vW8qwPmCNpZ0NTvAN63ka+j
uxyOEQP39nOykRsgx/5mFCRW7dn5Y0J81yuL1P0bOP1o3PIvbyrpePl0+gscAP549dIUNb4ugRQC
fngmdl7dCZYXdf+wh34NdtIe90o23NTwJ9f9CPy584UmaZ9xXRzZf0KCGdRbu+BPiGkEQo9F8kTz
82k0cc5n8NiyhdXV73BV/ru9EuRkRvv7Ex85B8aXHBaGnT3rOKXQZPAs3nMpkd2DCtYgJUnzxzYz
+bAtU5sR+m6iIAxoEm8UdGYo8JpPjk2FAfCwqFPyQUnLEAxS0RUnpqgmbbBfK2/CNe1YEsRU6fxv
mbaFioi5+nQhgcqozRjNpzh0zbiVahPETgvvweikF+zJ8iNE6sKeyGxXt3mh/XTFMXKuQlLPWPsy
LgXtz9wKffudUdsR+vSltDBxnpUQsJaCCo4qgm2hxvCd/ojb0Iyv+vdRQS/6Fz1UAg6GCn1v8bnP
9yyhA+7fDhODJQ3mBS0++tlngbAXeWhJWuhEWT7WBqWsOPZ1fhnLvnEB5wDU/p3TSe2N/v9cfcuV
S1qZKhu5DgKkykuyX//vRNtwVMB7ra5RTEmCJ9J+ZYHYMpN1TPQ4RROOvR4V2YGxS3vC1x7/dQke
iqyN2/Kn7oyuoSKfQ/W9uIW1T69qh2UO5Ej4+c8Ia+lxCh/R7N+2s8lWMA/LkHxa7tkQOXTwDn68
peC4kF1vaLVxDphCV8mJECry5mWL1AZlOMkcmN3imdCutqvmm5Cu1+Qx7W8Ewz4udqr3cVnevty4
cBdt9D+m68YftTbged04XX3r9VxTC0EEPol37f+U7tel+XknhRsKZp0q33QRIWZkJbPfm+kV2Vog
Kw4/bobwrG5ujwiZRlO/hpPuElhJzONDxXh2FVsmk5uE+rbY0jBob9JGiIiQQnOCarOMdsCvvftc
reW3XUIs3LJjYwPY6WHx2bTbZ/PZ0SXJpVv+zaXakeH6YcvEETmS9GUal6ohL5zaFfeNAcYykB+C
TyQ/oVQ1xNK0cr41wHupEgg3fFWnOY2tFSorYzlG1tUL2dz3WeQY/vruFKSsOdqf7hR0Y3xCt0HA
FCxgfrixxq+nclf+a17XOQFHQlxXvcXtYMjlu5dvCKtj1nRQLV8jpapjZ6y45ix7kpRI46qb1BH1
RbpPWW6YZWaDzvcGX/bQKQYcxPkMsO1Ef3A6n35zE6WBh2vBjJGBs8VW3n3nsWPCgEr28flhBVlh
R9yRja2qPHTSockjwx0vKUGAfq/ub1qlAbzg/WU7FDW0VaezCEkfGqROlsylG2QqhB/X68Ij9Eg4
BPMKGTobeocsnBhBQU1kvdrbNdq2U/XjF1IDAnYyIPEgj2HeNbNVuBStAS/ijbjwpEUfSdOc2Dm+
6f8AIvt9WONuQpeczPzraWoCDthMT7fOIlZ3cHn4D4x9QFHoDbxW2upFRkZRdsmtm/LuckaOo4i6
MnY3l9yNtmeYchgUbpi3tOAknh774TeBp54jZde7QbcuQpuJ6wJ+eAWtyw9qCkCXFcjNwGRUlaP5
hmIwAwbdpwq/vSjyPetdtkaaPuLsGEexvbC1GM0g6nVlyPoT+TeMIyKhBAHhXRbXCTw8e9YpsT+o
aEoLAOAJcP6LWkQD6Qi+I6HK2s1OdYqn5LDVfe8cIyQcU3xoHEzJTPVMIuQC5YnsI/Ce+fyhMopC
mNMgNtZQaPjqQFVeStaWlLPySgTqUb4Hr6LuUcnEehNqpPIuO5l/N0kLoWJTylawpmhi9ob6Gsfb
YQ+0FleN83jBd/OFOBvLQwn5cUrsBV7NRgxQGfKh4Pdos0HbMY1XSyioSOtCzB4B2CgthgdqSYdu
QPJcWEuZt+4G9oRtl7/k1TonBXxtlbvuGv3XbOjAQ2N3sA6cLWt5wp6s5wTf3iQCXcFOCwkKWKtC
VvD8VphbYkqOJtZ1iE+P/KZx6p8YNDltgsHq0JmapIkG5qJK/lXJFsMi1Pf6STihQi3IJQDTkCBx
4hWmXYnrHQexaVjfNa4XhKgyiaZqvrwKSWbsn52Aa6o2qV1i0HESIKZ6+ENWMDba/r6hA0EhoYS9
yYWjrkejoNg3YPEjkvHQDuynylV7msw4aSIjHuLVMzTPHbGm6Nx5X0pZ+FDP74SMb7BWohUjABxn
FqIrjq4Xn6beFb0Ktekn6R6pw3aCRdCgKOk2osmYd5T7tHAxP1gc+4rsqOPbuqQhiU6f0QpVnCs/
0DyT4UJm/zuY1EJO5KYLhWrdn0nLLN6SKv6CWdl3pwDpxHyLbuaZidMHm/fr7LZ/4AmFxge2C8PO
+QoWriWci8r3TLg2cfoAbc4p9O/ICIJmpxYatl0Z0Wm+ZyIjZf5ql2jFbE468+BzSVGNRkdpE7Kd
OCccgQla93cTPW68Nh2+zv+R4wJlRlaGloVe1j+1RuMW294mjQq6+VhITA2zH5xxL/Z0dulB360b
WeSuBHH0VPySaPiDp+42XiB7o8CMhv+k5wveVJw3AMIpT5wjTCeQhnwRXzPBlHqQAWFAkDneG+ZN
E2bsuTlzH98NBTFT58bNL/6JWrVKFJCfCiie+U7edjaOlUrlQ+9b8gcMFIxeejtBZVelDtiLxran
HP7WyYik4RCoO7/fC06zBhHwQqD2kVIvE3QYIPXtokku9RHJDccz33pfJdo+/nHs1RLr2XBmlef1
p2qLQfjjIoRzhjOG+56RpBx7iFDPYAKvE03I4iXjjvfZAkN1HSHGU/K6kn6HIt/WXgEj++1KuSgG
dv74qeiPr62UvU2AKimh2img4XswY9GdrgzrZV6oPBpZku3Y+LF9woGmncD7Ng6Cb765MtAFetwh
Fl/9/Q8e/bNmEkPMutJgmRy/1yCzNHzzs451YI2ZwaESsD+24kauxuaCzlixBfnPSo/U+n5UsuI2
zX5N10nF/d2t2SGMPWGRMdIItkXnivNldx1DqJ6Y7hDjer9JjwCddzuw7e47ezNHwWymiFcLEB3a
5iCKtthatS0hSStwG9xpRUXFsVRnUWpaGgsU+S1Rfo5CG1cnMZlHF2ZP9GFdTaO3qRCtSPLVMmi0
d2ub/0qW9rIc8WmBeEAuabRQWLIaE7VKC1qfII9WTT4POmv/q78JT7yh27Awpxou3F/yGLzSfHSh
mRe6dHNjtQuK/1+4oDZW4cV9b75SgAASQch4WcYRgjBZBuON2We1wT0IsPmTZuyvgEGCHx7Xti3t
MujpLKTn9iucBSWbRPlNJ9RxL0WAziI/GJRYNTktGzMU5UY1RHu75Wl4uGIVLNJaSGr8HrCie1E1
aLWgWbQhpTsUxksOjdjeALsTHd7G6KuZpksCzdlCwhgHMqEx/P9IyOLxsCI58I9CU+xyxSdp4bpR
biFQCVByXLiMjs5NG4D+QBjaLf+Dr3aZLdJDvodM7dHHfWCpLo2XQvMgiCTFn/wMQDCECIoxJ/sI
PVcnHbxpxTaxAXYDx4ftX0n3Id5ioupyor30xgDWz7qaNHhJY+woojm1rs+gXO/y/3n93tPWZKJY
ctJGP4Kg7e5s7ZE7wuO4YgjfxIlNsjQoG0ep7/3tjz/PqYiL2zZy7STT1fdzYcL1AH/vTaEIPD4m
pnmdtq4yCRtqXBeBtJVPPxXdb03G6bxpHTaYINcEhlmbaU17IZtyA0M1D/AvkXhVDU32ItjWPAED
d69wBcXtz8A7s4Bwp/Ao6TWPIi1KAWCQg/jGZgWBFVnBDJZC0UwGezkk5TY/P8D/7vjEDVao6+ai
hJfj8LH+YXy+W5j27mQUlhtiSKOIq62QmA2eqAQlIgncH1zvnJzwxiIORUmvt/ZuNoL9dt9ZoFD1
Xy4gDMKfhh71KDWE6p+YaG8VoWT2mIHwukiWL2z/oqsMEBHlVy7ayvg6DxIVnLX2O4r9+2cMrG6V
2uJ3bh1RckdLWvmGSsU45Og2aSSLB2utLLUrWZ4+sb0sLx+O61r9TrS/Gnmzom27yfMuZ2MgIsBP
qZJbKSxhHsGALTeWbuoO/CqFXSZV9kpaCLyghPvuZJouyzJilSYLaF029uN64CNHaf6tHWY2NHDY
uHGPExOgDhkWmagdhthLQ5vyIEqTv+9RIxjdL2DMOSroOW3XNxPQPoua7di3WMtB6tHogXx9Mrdg
DtXCcZIQu315VX/zt7YblnsPMrpKzq65gguNLsshG880WnNWg0zlgO7gbq+rjX3W7tiy3KVlz7Ge
P7xej+9Aq1T7ccw3b0tUNDQ4e+QN0tHSClNdtmDTSLxtuRngKE3+CY80bK99qoei38/UkWsXRB3O
9k32DV6MRy+J3pvtqHoRUtmKq8j8NvldG69ftE40gXuD0QGnnJJyddVqRO7KWcxp1TrwWXyc8S07
TSUBygsEEA7Fe3aPn9aBAE1c7PWYJnbhBbzEBH4I3VS5jHOQhDFNBvFpJQYGOTUSJlFuAsnPUcH0
R8A5ySXleJaBBOL2QTYerhYOuF2L1Bo+qqr6GYoUK9ynPR76uGmrHBY0x7ejxswH10vsSNLeM8Qs
6j4VoonSk5lv9kK+I/Jjp5VF/MnEAWlFDAfiJAR9ZG6UAfEkyguLnwDKVQhgw5S6BXovQfQ9GEOJ
2PFhgDsXyReHBc7y8qFp2ErZ5V07qATQN9UE1OPL8XlW4+dSF/hH03y69mv+TNOFYQRe7jVJIgMT
pGOcx/0PWdocRvWcEVv0QwX++mmSa15VS8SReoBYh4X+moqmxhU5Zj6TKwCBYqJUn1DwWdm7egjV
byyoB9r818YIm8fFhRNSJ9A0UEmj4t5LOXeyjU870vHMKJUA1u0dc2+C4/VM46PbpOK/2K/qQUYv
U+/Z6J8mbUpUtRPgWecjcVz93zbtqvCPLGnlA7YBsx6T4TIQS7xDzM4SMYCuZc0fv7sVbQuL3Xpm
QhxOCSX3AUjAcAnBZQX7S/K93O6tjlyd985q4VeIe2SwbwPtpgQykcTlOc3MWtyARLNx1W8h0Lkt
DkLUF0KecGpdfzdxE6LOY3BfIYtUhR59yjZy1iEQl0g2CdlxzZyim++Haw3ZOl2sADJlXGaoa2tm
X2SddH4YYtrBU10j27C5N6Ckb/LoKwQqKPiEkqLVzfbUlInZwNom9qkQu1auHmV+z3mQkDe2kQPB
sD0kn8nqud1ObwK3Wx7Ia62UvEwq6aPDQWRpVuKxuz0fJDyYLNSOvaESauAgJlAJgKUNuhSnbnCj
pgDYOEMgTL3pwJ4oRdlunWypkxIeiWGyDt5LyWrWBJAI+Hmk4g9jAVW8Ebdo2ej5fSUuks/Kx3P/
7fpFnnsz60mcW5DVsOM581aYV1hr6DauYwdafcbETRkKaTJWSr9SSItE1a0qafVtOGKaG4Lblt3b
6h659suzZo3hBQzR8HEThc6iDIdhTSaTRRYASjoy1QHT51ZtDl2g3y8t7X9c8vxRru/l/ZbdZe3W
zboq2R9sxTZJpbreQvx0r4MxvjfpiRffgmoHMI0Mcvs+3yrYaz7H0f7K6VJ/fRlHXPVXO7AKoucq
x9jhQiMK7IvsS9KICrJXWjHX0kUIhDs2pzy8jOTiWy6l/7YfYOSz7Ijihx3cpb9FujZcm+a2ftlU
BO4nnOsIbTlGDerey40sozp9OyqK+uO9BUv+5POUoRcDeEumrPAqhYxYbgQoMPQDa3NrJy8CIH8v
+UDqxGufz1A4fTuv3mIm+ASOw77nZ/ghozvCRuzaETP4TnbjMHwkpq3FuH1h8KhkwNWM3vEPWLK3
ijdji0FXoMTJMUJtQlu7NrLLRgNutNVSqRgE0Hf00c9/YcAU5Tjgkm0R0e7PKl7eIXAVGn15UB6Q
cTA++9vf/qa4Evga8i3f08JuWgX5Th/og036ZzNNKsZDSDFfryKyWxU5SiO28jkKx0ErTc37aE89
0VL0tjMcd5l0ghCnQ+UaOVSChAI/WzrSfd8XnY62tAKOJ+74/JQUpb5MseEfJQb9PTd9ww3beYP3
j5on7CvNRq5HwPB3oyUKkyD9pFizeRnyMa585zVnd88UomRwbm1BIgMlvcjjpJfUmmDG2NUMRyMp
BsYD+XFq0ey2EaK5bJlWP5wXMMYHWnnP1Tw3xDubhmze64he3Mpf6+vEq6bQKYaRDwl+aHd82Io2
Yeca1efLMra7x0UrpXKV0TOVCs3VV7kC1tv6bjojBViRZ7urGFVZspL+9G+MH9ZY3tryMqNyAls5
Orc5e7HzqTu0VWx8N0tGEdvUygOuJtl7d5IpR0BsQ7HyTGdPjqcc8CgsJH6GnncyxXSzwCHTmLxI
zFtxvu+yL2+xMUH0BJS/9FlZnLO1rdDK7ffZCeO7UpzeSF7KjEg9hgLdXjSg5emkuRZJp6gvCYGd
imOlRIvi2CtJ7deJUwd2lOYK14m5PxqRT3YLdA8r9uuP+v9ZGVAsnRCBrEzawkhQU42+QXujtmwf
M/6H8SHJrS8Bbry5Z91fmjf030BHbjsk+y5DBv78w8Ax6YDVekduyYx9DRkAjJ4X8aqdNkpFxCWn
bOAy8K3oVdcGLewZocwc6uk172Xik6+rAq+Z3cD3O9+8lHkoriS39+1gL1kktGPrrKQRS//o8NDs
t2JcmMBi4Aj2xveHDLCd4DE4kaBuFMtcL0V5HR/9a1+pIzSaEHjwg1DEU14ERfy1WXfh8FAkW0cf
K6ts6I6JMNMkpXm7N2WfE82Iupzo5FSpLldntytKc4S+coCO9HStn0cNoORRXVRpapa46j9ol5cI
xvpMtRlvvqhygkEz0RROQbKKXfNV82UDPxGU1ztgNklAEPd6hmrpsL5lENYHWf9iGerW0M2jVmt3
yE7/AiQRjlwTpKRYreZZbT+1zbiI1yGxBONmdy7rgmDLGXavAjLap8+C06DZ3/TSXTr9+XaP7B6T
0/liLXAZjOjpP6RRpUx0KCFm2hBjLwljFE9PPhsCfSEyvJRDGtZSLFEjOA8MVHqdsCrBUV/t5VQ+
SC8QkL1MJKeggFXYU2Sy6/AMLfBRcsHB2XnjPmkt8N8RYmKV1yBZTjAqRiBacq/Fp8bySFcaVrjm
BguD+0oIXsZs7kyyInxalDwucfDrqoYQggG0n5YepKEpxFHqmQk8J8ib9lUXeefPkQtDA7dII1qO
oyipflFM5gbJY/DXGzwZPDYmpnxM/IWJA+PiEjlcPHBvABGCYak/8qS1tEVO/bixv6W4uAT/fyRI
fPUDqfTS61pcCT4AOolbKaI1YsfxFkHQa6rj2GOv97Bjim5Cxym3Vh/scv8MsVCDcBdpbgbCiwfw
xdHWYR/aXlljsn5Ne8QE09tQpgOmQxKLmVSGJkoxMTA17fJvXs1nVzoacP3MQaYhv3malkLOs8sl
KvJhDrRPaqwYG97WWt7Yy+NA2c9JbEk97567f4ZT2PH1nj7uC8hBal0lOK3irSdDQDvUOrhfDqK/
KEJ6lFR08Xv39pbP8gEaqylrAhI0z1SrajnBuK0/zRkJC2YVvaAdrQh0sp0FjeX53l/wlKJqkpHz
y4/95NH9EKfPiLA/xdTnVgTH6zI+H2pu40kqHEwpguZD4t1U2yvoCBD0troW1eed4Ka2zZvJH/V2
CEmP9LfGpFA3Ap6vjiaD9ClbUWaKHYpNZOyERelLsA7Qd6LC+0/qe4evjsta6Jh08FYv5nHqcbjY
ADv4yR9bGsRuvBUnOe9y9PaqPlUqdSUEzQDrcQ47b33G1EuiBlRoKxhLDn3FultlQDoxAn9UUGfD
HQ+fFuE3+OmH3UHCGO/vD3gxQIduu5e1xCMwNmsgNb0OqLXYQind7VDUB7Cn3VXJPcfQ4tps0J50
8Lw1WzQrLJoX42gN+K28HIJbejQeHgDkyLIbyhrlgPP8xAHdTHhACiih4MayitH1Jh3pXvSbw1ra
M4Prj7jVmcV9S2vxJ7JWMXvyKhmP+R1IJPCe8CrgXZCR4BsbFWfvZlhr85KP1b6+g1To+RnRazd0
sofdm3MItnjwd7qXtNixsoixYUK5BRM3xXtToUdPVDp/9Uqi5TKhiyf3bkNFh5SUyocib13HXSd1
SaWpzrWpAVjtJqxajOxz/EXgC7FzBdtwCJRscR6R7avqGVU/HPXBFM7844R68VMsbKHwlMFsbMUa
IRmHvIxYN6EvSj0RDwB+9s5PeNyN94fIg4Ad1EUtXvfX116Mu5lrA+HfJsTMvVHIf4RGqW8IlrnA
zXjU8Jff8aZwnynOpKqNKll69QTvk87dytunWow/wsCAr9/G1zexG5c5G/ErwM3M2PUkDV+WJoPU
opNHUb1QOSgh8OsmSZpyWvGbGvSSmWT8Gv7x+mzlGDB3zbdfTspF4xXYDPhYCF6MteioZjMuwpZV
os5j2xoizavLdEEkHOlVTOgKHb1tjNC9DIW9jqbp6N+CTyrzj7IoEkgPPmJnSspNeSM7ZI1a/U9S
AqRQY9kA3iTnAsFTAla6sTIBVAW3TNq/mZvoOlb2B5awhq73UPkSEMcHDCq8yHu28iKohiOo5VdP
HAfyktgivxeT73gDHB7LXAMQKl4XheMmWnKe8U/qwbjkYAGnpzTaDr2ygccKoeGZVUA/ON6O8x9e
URhS6UM0DCtpb29G2MPfb95YiqEdn4vLyPLHuw4cr+r5Abk5S8ZucPvGYhrt+XNjUeWuXdVBMZsY
OERnJlTehbpeZNwj5Rfud3C0biICzPM79TPgO+0VD7H5W3o8C5nGlj0bAkOW0j1WAHiaJWT7gaN/
vq2OsjAboYjPXZwbx5Uv4ngXE5r6oYcxt9NmT6JWt9gFrOEzG5NuJrFSRWw1X640zWiHZvypDCup
rj+2Zq2J4ZP7THq+7MdWxfznCTc+ZhjicL3ch2yLli1kDFhfKY3iWwL3cgpYEKfKLtItQXQfepUB
lKBWP0EEV1lujZdULP8P8PPyf1e5nndW1Ja/fARs/7yb39yKSMmBR60lv1SEIj1sa3nT79sRyzhw
oXuVXZcSq0skor58KTO4W0shrWMrFGVFxNMkaRdCu4jfYaWrzpNDhvpX9PAaT4WHytD+aZpmyt1w
GvFzPnnRb4lRHLfYcQ0LLrVOCEwmFlwVWZYNQfM8V9dvw1+amSoblDlpscrAvE0lzrX9VxKml4NA
m9nygI5YRAoYFMjjMj4Dwa+3pRRqf/KHWC38lAhRtZckGajGWlh4BWQtPEi5FqVADu9uxmbEX+Zk
DcnCJPv5slqhdHzOh6ypJH4XnXkxNcZgO77fZ+XWe7zGejMDQys4Q4YcwuuxzL/bC5/4kHsGxZaa
rOFMBfOCRXxkk6ab85jI7uhl8OWm1BNA7aGjejQEWeJbgV24JcqpFyScjRU1DSR8tJyouzl6aKkO
Y8eM7mKb7SrVjw6HWWBjxlDoUkggw38ThhG0yxa/Hi59iGs3vbfNRt1+s2FKOO1cA3baEhQQWZ5x
2KrCeA7gGwOWG5c7cLiDyhF0rHgHRtLWEeIrLb5p7+aEBFpgnQWXNicCt6iRR1JatQ70Pgzx+Fh2
FI2dJ6Lccu0wnjVNDW/V9WZBa/tE54ou0qurksOATVatS1xpjbBoJZdR6uxTCxRAYDQc8RL5WDaf
3vSRB5K9hrmMe9cady4KW9ZXysTMeqkTdu1AVkz0mM6TCbFTarry4HtgYeIQd8X1DdqxJiKHPvI1
3KxXsqdIvYQpMbvpBGDER/XvpHZZUbDvjBClJ6bz8r974hAy0m2CZ+FxVqweTNvR6W3EmbEJKtw3
uESirvJyA2os7a8+dfTgcmv4ssgYWkJ+CnkFooCjwgdkotAVh6I2I0aVqMYylvQ/d7XWtiF9t8Pv
pO5yDMrc0H+vGNokbhw61lBuElqGplSzs0th8PcN4jWAh1tLd+9kd6dQyxYlMgzMSAbEYGoXoEl9
pPKb794RmRhJ49NS43YjRuzpju/d4Ulzbyf4mfeo23IJIyTUflyIS05NMu2bTqMcheYNFH4jJv2/
+vdrsz3nHnRqFG+OEXlLvXIjElQIs+Z1dlLnHTCBbQ0ZLBTKVRuxkiv/xKMoyNruG6yMAzjLQtZJ
PmVmAXu84hqGU8sq5T8nRKzcFtk/Z9GS8PB4EQXnurhTyEUaLe3Laldd8YzfAg/JW9WhrJaOsscg
ZsqoC3lcJyAAsV+MS1aKkg/YWWC0+txZznCMCsZkq2UnYuZgODzgni4I3vWmP4loADjLZ2nkwcYW
zaNUTMr6XjeOXlGetSBiL0L2HC5rgd5gdFqxgDlNs9IIWUJeyawQMp61OrMRTGa5Rh14DkurCiQJ
iajrY2kKSgpndey32OMn0jHWHuXw1fpvyUL57n6z1CXFIO9OQu6TOgblyo2OJqdnwKlcqWpSeSc0
p3wba5kl4dfqq2dmaz+ESbul9ecsS6PUfU2s6X6zwnnLmD9BcaM2RtbkCYyNxhGiq9u74RiBnUVR
OHIl9KYI2nlKhKt4Xb25uOyKy4KfOPd/fH1oLGPnJz/YViCJiUK7qj7WFOEi8so/wWl18NDsXTsW
C7kAhy82QembL6XMum+BBFNtqx1PI4CS+d18qmkUrfdZEOCOxHLtyQkT6xmdkeC7BeZX9yr8txV6
4zpv39XBIV+FxIYc3VpPwXXCNi0kwUZoUjohpKmJ8hmcUlLj65nNdUuV8F7Eycyc+ggrlAXOAaPg
NBtTK9mrh1rkFJ5hHMI9V8VAEmkzFLs0LchWY7IHofuPDXOcAuG6IC/vgBso12vlNHn5A0x9oWJ2
3pIMTODlnAQnQnK+jlpt/eypGIuJUSPNVHJbaPLnrjJ3hDvFbEfqTSpLq/o5pzcdWxLj9X3pQK0y
FY/FnT3zo2go6KKOKyrFHNP1pUuAodYjkwVI0uLLlm3t0P6PSF4LWDx0j4oR3eAixNvAEz+pX2h0
DiBthXz1Ca7UGMyt1Vh38LVdF0U4AYbxySmrHRwcT9qsMy3y/p/UI1duE+BI69lI4Tzqz33wAeuz
gC5T5rnCiWD7wNcZvZwDZ6roRk8cTNGTo+p2cIcQshOBppgWBG6oCkmFF+y/blcEkUE73rjJb+d6
eBSxg13h5/GIg2IwGj+yVOT/KXm6J39kjr1yd5SfHXUxeK7XxZnQd9Fgj3Qc2aSwk6r6Z5kW+iO1
EdSgX86p4wFfrREcZGugY5x5N9frK6Okkf7yWLRtxOBQVkUHOIU8XQVtO8kiY1VPeVvtQ45Tuf8k
xJDnAPj7GojGZL+IY495sgI2NmeCM9WZvy7bfOKHX9CkKmOAFDYljsTJd+pQ/NmHRkYDLCc/+w/8
Fv/NvWMlayX0Gh1Cxgg1AvGC5GuhtRWf2YA8kuq8FzANHq5Yf7KTVsXbcc5QqP4NdnwCdCEN129H
AcGwmmYW29G1ZCRonC6p9QnssBzQ9I5slSfPUuq7yaBTQDXzgDKbpOi4OafPUAumnlyp/gGE19VF
PqIyOXU8tFhCIcyvJFl7vFpWWFb34mGDCgUuaztPBjtVcSmgJhBBD6G4VIAXo5+AuhpGKwNsP95Q
SAY22GW454CkoXiHv5m+7TlLXig/H6BQenc2bhODivBpTn4Z2BWDAZ43pP+5zqL+s0+qM69daeKs
D1GxgPosq2hpsp3XnlLVpd4VatXFUshASBiZGUDi0JSYAjK80Alle/dKOwwZJryll7LkVxnI28id
9/ZoNiIhLbjeZKfponmR6qX3lbAW0waKdjQ+DPu+waL9NUkdBCcBUAxutMw7tWAndi+XiqKjc/Dm
Teqhgw4djSk9EM7UfZvqoRA4y/sPrssGlMO2slYO9FIRKAEGTNrhlk5EzWqpqC4BMMhYTjrHgm7i
ZndenQLQtzoCv1X8qq5iLXrcjrwdqHpNDZCsvt8NBjVNmqETaf+MJSzRyL6S/WreAlN9Qs+i5ni5
h46q97/rDnd1SUwgMHkaMeI1X5AsbtiNpDtH+fmF0FiGGwTwLGjSsCImkiK/aZl9A/9PgcYi0TY9
eQ1pfqfbBOkrvTwnzI6VW9dcto2YULLosms6zKD+ZfsMkuK0bTGB4jZvCvSJBp/d130dwLDEKk6d
JgTgKLafDXELYH0+KaV/F7sS+pgYqAYs5fRkxCc9jpw1xwgFtLX9LAFzrTUH5VOIDR4GK6ln6t6R
15K086dMtryhPRhiz7awyOsAiMcEU66DSskbyd1gf8wtLf9fhcdi1TtvT9NrLIgWZR5B6x81YQcu
UaY1/fHselAxPsdSu0B7GaotSqlmm71uwiKm0UQh4SE69gUGD+h2s+hgqCl115EV34z7F18oydJJ
MxgjLYEb4e35RIhvq5Yo0eZwSHRnmE9y8H7YNfc1FUTbkiyyCq+Mn5hOmBCpDMppA5m7QBJ7lcJZ
yscbqpYveD8FjwnSicUt1WNHO+DTA0bC++C1OxKRJSxv1gpdtIonX0g6PHExFehpBdKlmLR3tGyl
b0QnFKvyJeUZNcUpmiJ1iABVoQqlvZ9Oa8xyca9pCQsVNxdxl7mSEAZyTX9VZlTW3JwA8djO7bEg
xnlL/kg5bvZDKXKAOyFUAWMGu//zG2a/bfTjdWI5rlAoEW6frtpZKhJeLKshRSUd4kbUAsGYlPzD
sEKc39NYnL0rzMBhhf+B1NF9X1SvBaty5p96kGUtt1jwi2KfqBWTb8v+h89HofLwdQugM0QhYkXI
KrUpueUu4mFHmzj/BtWJObnUt6h/O//JJIgBP3QIvNMVyCXBWCxXVvnicghYAmqoL9vW0CB02NUS
qrn10b/dcX5b6JYGKCz0ShPk464lqLWM4aJ3bMUy3rSs6gCkzN3oeOVy+ST6HnGqp56rgGlT40RD
OrIvSZlhixQa7NuH6v5gooRnQtpGU4DFsj1RgLJkcu16aivczXbipe839b9wLNCMO3c4BiSF2An2
yt+Han5LEBnKBkq7Xu1k/GF7ShTdmpjr1wjxJATVdqCkK7w8SnAsqFleEbwJUdce7D+1C/hHjSYo
scHGP6wSF1mtU+OpffI1FVYMpSMWWx8tx+C8e0xt4iKNA7QfNT+OX3l9G8PSTXj072GO9qUxVlWM
EoYbW+dI1mZReqMONwvgt4rDpMhXcaBAcK+f/0rDWyNM8l4SIWACrEUhxy+mBvvZoESk4mMBxr9A
v1y/Doz4f7j+UHqL0PjXPTYtgoNhDOpfqQh5Lm37JK5owoRkn7s4bt0lOzZD13Aj/WkhjiEJUvcp
CTi4W1BlB+JQlMIJw7pw6s6Cm3y+5O/EWQ0j8y+4/fh1Kd5iHwYaM/CDSXH/rBzF+kSh74LU0v0X
36pcFmGerV9HivtbiYN3SBBNk7b4NQPTuF7qz+D1rcRgNxxwDahhOXxSFLMwF1pYMj5KtTvMs7Et
RQlgcc0UeseT0kMahd7KAbbVywNcaIOjI0/hMLQmIOortbDsCW3FZqaVVZ8tI66kAClvlQF3fFid
lv3J17td2HNFR2yAklvJqrwQlTLjBI9yEeED0lTnK34Ya01+xLJAiGT2sujqZxjQCHcgnbihWEHh
FNgrGYC2e0bwFze1lhk2ZtuHyBOqUq5/IiulaHGk/qSBUDGIwBI8VHAOrPTPmaCx1VYXXBQ+vh6N
gDw+hrxiLNZ+P02GGZ/LFuLgqdOJQha/9RvI/EK4a0WvYyg+H30uvStY4xuFgaLnT+QCP7EfNsXx
VSiX3r9c3iv8a7QUM1leN/59QF4/Oai5jTOUFvcafOkTpGAMzybjNzk6onmrcH3q9vBSrrcLwJQm
EVR2QKEUETcfqNrfS5raBQKffziH70KNaiiunAEn9G3RuX/tPViHwh1Wx4QK5+LXLvI+LrDHQInh
YEmxKx5/cfSSXOTRfFCEXAKcfhAR6sr5lhi6V9F2KGdnDcE9p1mopjZR17+qnm/vJStMFQHzIMsl
E6IcIkJMLlPVTmvFE5HzLu3OsodNDQ5rluRkQDIkmHEVDD3EmbazIuS+R73Y9KUltiZAYi4ySX35
v9t1uwMZYgTkl+6oIAho3/gqZZHcGA2CMJfUPt7zqE5L0ftuWN9XP2r55k0rbuJyVdfXCn1KegDc
drTGrnPjxJYhR0yerbUVXWWzJvLYQH7UiHUJW5uhm0E1xIev3Bh25HIYIVH4Eai2CMloH0oE5bwY
Go0Y+e3Nh124tFd+82/P6b1AwwFq42P+LQTy2Bkf4ZMvfW+an7wIjHg1w9dnYUOMY02jlZlcD2jU
ReHIJFJTcyEF1xf8ASEbJelKGyUzGqu3AHTF95Kh4fox+FPCjSZ8fY6WKHkm0Audk7KcRxCOaBbO
VtWjc4TsSCQkOrzWWeOijQrjwJ8zoWiOCoYnzVd8ENPiXxkU0phm4yYu9jC7PI4QlHSwbcfGnUik
D9/ty6cxILOFFO/Gb2BUygbRF0pOXxuesqEhq6879WTVIVYuZYsl9fuoQ9ACktflG5xJd5FlrinI
ncOPxFHoFjxSiunyktq197/yuNuFNQKh762r0DHuGet33U0ThzeZkUQ2WwD/cZhicxd9gSW0yQMP
tH9EP1Bkt42PPvXXBNGNwF/wMCrAAGyinydT8hraIIrRIKswIKH9SbZAMHOLrKUu/upfe1Uz2fy6
WZYKpfCDOCZIKEHYjRvcy2EY7wma2DqN8vBqfJTuqGQwUBKDNuCth6mEZqg6421lQaeywGA8pEvT
yNRQH8xqfOXEdwI6LMARQdK6/S68toX2av/jLiJ+PKHIAMnHQ9Yk8dfnxTSk2nAxWXOskxBtr6z/
RPgYo2P7gThBArHddU5pem451iLU9WyxxEWmMHOSbF3zCxlknAsTWRoLtn46s9yI+bF53USrp2iW
V5T7xVJVi8rjOk0SlQYFcIkO8VQYtCyiWmpGK+54go7PDb6+qORtS3vgpJkRhcgwDTvbX11Myn/T
HXZUnYs3zeegyBoQpmeFQaDP41EV6BityEpJplr9koR7t9TTKUqqcliF14nNPszIdB3+7gHn+AaI
BOKvAeEBpKYopn+KY7pKmGZE6IuYmSJ7DZZzDQWVIta/okalRleoi+zPJ5nI99fmDvKF01hVoq11
vgnkQwzCzT+ghX3BhZRhHEcUkribF+0D2TG40agIwoG3wzD5A97iIpp4X3ElajhuN22su2+bcB8S
Vh/z1iK63g0+a39u41kSkdhOCogYtWzeKF3/mWtEMxfsXQjG1iTehbjAwhOqhqwxYTB36u3UrXA+
iABgDKJWVZbSuKmgfAdGfp2XWYculkkbDQZqY9I8wyCXW0Ads57X1RqYwHuu6nTdXqLIE5149wCl
jZAAalaseBK0tWnqCCpz/atqwJpIBL1+GnAIm7BfLPePBsyeIuqs4rx+0XmWPutRyT2ojczUBmEe
vUEFTG2PjphJqPNxXfv8le2HZ8sFDAB/BISkF+LP3D8Ej7K8LljU9sHQpuda2wdjTqFkdivdRyOi
edxCjlH9SlADwLebzR+DaozALnnm2c0AWiuslC/9AK/TyOVFigrdIGDjaRjE1V5Bj6nGNy/lisT1
kG9ozrfKfgqtAGoVxyIaR+8rdHG+Exl5pwRXo6ofb2duOtyV13PqT6T7YmmNrdj0wpOuUqEdxqxY
65wS8b5FO48l8nnJK1Fk6P72m6pr3bTlY03Won46ChPGYu/JGLRz0oSj2BxMpsYlAxEEJgymwNHO
q6JeWlOl3rAJr7etyKRnjAcczYNpk/CD24/VnjcstwHxJ/9RDpSGts11vKNNnRirDFJ00cObCbQJ
qzGatSDyv9pW0AP4UsM1YQUTFEPOM8hzkjMd4ZH4z7SbinpsgcLKSb+vv9bo5Yd6zbGopO5uLr9Z
joSH42VY60YUgFQmsJaMcqKwdqK/4qkQVf83siUtx2Lc+pl0zHVFJNZJ5j/Qy0H3ppOo0CVuKn5b
W4d0MxPoDtmzNot7Gx7Myfwr4DMD9kHr0OUa7Kk1byYGlFJLiTrFSeUnOkIEt9v22VLPIaYS9U4r
pGSGYztOoirLSIJrFYQtq0mcSFaLEKrwrmb2ZQc0VfgLC+vaXnP0IhcM3bCvV/gGZMxm4++jEQt7
v0UwxF1Yho/Ms0cdx5omFO0SvNtm5d6yQJEY4TpT/5omtZlpPmx/p3IIwz7yCWFXbDieiY2VI8NL
6Oh+yCR3cdPGehcJ1ucGHaJG1iUzdhBQsSDO2TQ58rwzKbsN1dx3flT6+kZ6EW13fiXrh6yGtX/4
QS4A2SOd6R6UliFV5CGfSezwz//Dc29UAXv1at/owvoK6mjy+e3Qw2FuIsKxh45mrbViG7a7j10k
MKOOUz7rn6xWyZ9WSL0E3oDnWgMxm8npTqxofaljkSgZwznbVkK8WSqvDMouh45eDvj6YB0sfcCb
9bW878eUfPfAylq/Brq2BFoc0CvEetPYZ8j8H2Z4wTvod3AZ4S/95jaYTm82TpT5Xq8VypXTA3v2
niJWeapinpq5mOLQo5ycNrFJjuEj32t2RT6l0powlZaAefNsVuwMuLUSZZXnSHK6XcV6cSiX12E5
SNxWKz5P48PB/ZJMHEaF7yx2SbYLjjk8wcVm98e4LzrLbyoL8Esefql8ZkJq0bqlLQjxEBShamm2
VXy7ysY01kKvgnHJeN8Lmsl5J1QR/rCtBvhNVX1mll11/8zvAKB9E6/5s5gBw7+yvrSF9Fs6UpI6
y8W0hi3BFsbr8iqygV1tC+M45++0VsfBwDxtxXLTftHDIFPjzEKsckupRmCnLLrMgmSe8Z6kGWpL
SDhF5+LAqozrleBjK7Pi2UMWjcFFJsBvqPz2rgAoiTiG64ZXt1RgosCP5+WwqGPXCTihngnRjWDp
GZ95UqeAPgqciA2Hqqq31L5/4G/l3xf7UPDg5SITXmXX4fdZ+plvS79m3y4baYfEHjcxLvGfcx+f
+jtKAWLPx10U0y6zisIBCHSZiXKHYwIkZ93KrBfBFgpL06FiddeSMXg1LlyeMpiQ38hzBDlA0G2h
FW6KXhJVnQ5TplfXC6JpTTViWtH2bQ1P/tWj2y3LwpGAEtrcobPMh0gdWs+tbVZQu5ziPzLL++eS
91EoYm9VALpookIXWiNA6E6+OZWd3FxOHAPgZdgJlUfqiS5La9UGYflII3ijeU1VPXJr+8LNxmQ/
4M3J6A+nsjoDX+pSMljBPu/GchG4RBUPZFgmUo9JrKD47286u0W2pOZxiUE7bFsd3xFrfjKzV7TX
QBntIUGgBY5ROsGRgJOMb4dnvcUcNIvVwqVVF7W+JtYo9D8SkewfwthR4WoGbZVpDk8RGK0WDPIa
zwsFS+bZj1ZLcVc5Ws95fMlhGJ6cDq3tU3nuMTFqCcqsNhNquQTC7ryvIORywCrI/xw3CMttFf5Y
UizYEFUSkTM/xUCx/7PUAEpkMakTWbtEQnyzslQHOjkNvw3X8kqcMKIUIV5uLoItsdQajjdG2yXx
ClSGIiZXw++WQm7Pi4ZYTDvQ8l6sygX5aExg0wy1UlUsaaNFbM/YWhQwJfqfu0N0SOfzbltdrOSQ
jAbzWzRmqcJYV9HEbD/Fpu7w204mBWoy1wTSR6pysteZRoKfEQ7pfXnx/7WxqEIohrmOo3ofR1GF
leXCKH/crbnRoOGPCL9VG9LzRHSoVMHWM096Xtmkion5H/a0XCMjfOwF72dRzSuV11J1pRk7zJFD
rf17HzUHhoq8qJPNC83nCyzsporSLhciaT1d+Tb6FFv//R3Pw19n19ULQKhyVglxoY5T8GO1shkp
R2alsAYlhj/cRjSDMInh5WwYODTb0ft8ePEkuvIZUdHoazgO1UewLFVWlT/Ukn6pqzFBoRyHVUnm
8yauLHzMi8m+5yYL9wXhqNkEkgQGzpgJ2QfjUFVhRXqcb13e2zBkDp7Rjf8GIrH8kbkeilseXEPl
cp7GNuaJK3KM0KUdXAE1z04NuLFWO9kTPs3dESYoCdYSx6mkgoiF2hmFaLccXn3QFbZXkeBZtsg2
Y2VqtMnxA5v3LXkezxxqFaev4Q+FQs7+j4lxAP/HWQCQG5EPUKY/dSg3vYIVstmSq6KKT6aL9wKJ
t2CG8H07xZXR4i0sAbuwyPMCmVm98Hymb/JU0gugbLnpyrXplyOvn1r7gNO4YNmhI3PIYbXmisWw
N3kO7aj0TwfHOIVk847UjPKEXd4pmEZbDhEcEGaqa9AlaqBkexshv2hVIM5MuX8pwE5qi27l99Nh
Awq+tysZiAAszGB9TbelcBOEvQvDfElgB4M7rzrVx2xm1dq79vBLlTaPhgvMOyv15+8yEJ7zNYQ/
eojnG7QdkMzYjsMEaqpLgpmDSzY++IFNdadp8gcH7uxMgfK+5ZkQAs7sB1wdIapxZ9Y/0NKDWxW1
zg382TETKUG9bX0gRWTxj2gBn38J2q2SGsbqKIQmrp9OH+x2nwAvW3cDp8OTc1ynUwt0uJZuNQdP
VwvwSAlWiaRfEjH1MtlepY5gBW2miLOOHnvdSOn/9MzdIdjPkaHYK+BKlV6tEYIoN54xqfJnFQKH
xwQvTczw0eUExdjvstHFD12baO3OHD/jINUsGMNpZvl2OYUUmuLUMMUQCXOWRBwUVgml4yCoGa6N
Hsn08pNd4v+pqJfDeanVQCcWy17EdunQiK2OsfOhdyVy0Nju4QbZP330d+lOJVi+2apiQ4Wg5153
LhXpbxrFC8KCY9VQFL40C38osJnE9XmbIIoNvrkMy3DvHsDMDRkcX0rceTiEQCvACgwvx8uyrIP+
iA96dLUE41m2tFY8FfoCReUtrZbhJkNAfZ1T6yBpia554vNE7neTaeQFWkTso7Jd6307R43Sm2RO
s0Njsdn8si8hgH9qiKQq4QMctjm/o2FwFYoTsQ3qj1QiWga0JOtTCeR/WllgQ6YJ3lSZ5TNg7YQz
q1+rIv2bh7C9DPSgSoa5RVn0lx/3mbWMF+uweF5zJ2xUWc3zDUoGpRn4A8YT1pykjoA1GyjoMnRQ
QB1JvKKkQCCQyHBLTL6gIcqKVKGVn5hGUzF1zy/Iah1mJcY5C5FZJqhoea4JYVJ/sdq2GYNJK0KB
wDvA+iOFVox7MfTEbUgdhRbGjYGsudjd8eI2pGarzQyzUN8OT1OGrEii/rrUkI5WjrNSRKD3YRZi
f4a8DHpRoNzwEZYiTLPN4Oa9bS76jwYgGVfmGI6F+Tb3Eqcela3LtpqHN7QbtCpvUm0JatKZWE8Z
WdrLBOn5o35jMxkQqDpeRLx8c8E+mD8OoPnxgjp+vWQyZjtFKu+Z1fjQdhd1S99NxtPhPsKpJTtY
rEzxnCQhtt9YRWoVMpMopc22RkEKRL+ZrT06M6qbgm6jVgsCtJDD1rssifNqlljTgRbdxORGtxlV
T0+RBj4NdOKBij1mMl0ZdMpHu1cGEAtdQ2JMrsP2sRuXkgQhzKo5VZ94NFgvOWnJbB0N0hdio67Q
50IvO+zR/ZeN0rPsRVyFn1ePNwwvJqgSzJ0kUmtPQnnIn+NolbHAVvp03FkSXCfNrgfWhw9p92xw
/QLrQhXqnumq3DE+iuZqspfZJb0ihdYEqr43SxQZBiHCa/GkdERbbD1EeO0W59UB1cO+CYiP7PB9
7Ae6z+hB18aB35dO8XYR0IK4n5OuM0MO2ZD0/i1+8o12Wsy2nloJhHVbCZAmjOIB2fM8xMENerEz
XdZtVfe1kGvw+Z40SnRF+WozjbaOgM5fbWLgodkiKy6kd2PVuo2D658U2eQZ3obNzvRBxpHmlV7u
E6BWiD2SOQkNqRsHZTRVQ04U5yg4k/Gqxs3QPALvyu9sQZoqKI1KNEcLElrodKQVMwj+dyo48srO
/dCfbHYlHyaabEhdo0J9APhje+uY6fGpCKFD2j+jJQ582bn5cbnj7J2SEbbOCkJR7T5c+CRa5i7e
PDr/sDrmKD/kopk2MT4hKdLNRvEpsZH+2elXMVXf+cTFWTWiiCRaqHoJtnd0plR31NGNLgmYqqBA
fCtqdmiY4rcy836lxEfp2RwIq6598Sr2GjWK5COu9hMnqttxtaZAWIWR+kMwcVMuLBYstjxsCoMe
nG9It4fWUk4DnpR7AeXYmvMiJU/PcffJf3EVmpU7lEAmhh+udgaxhfzrtNTHUl3T+BNePjomf0gA
7aEPVkh+dTpNYH+GawusuCbE410tH2Qb/J085l7iDLHXBYhntyPhxr5t/To4W7tYOQvp19CwKq7l
LFSEYq6A6+Fu40tpk6ZZyCuS8td561rw12co3cXM4+PwP/lwk9An8K78WlLFea55WMSGLKypcQ4p
c8eeWXbqjtMvqhi1VVErG5KNAmU9c6BgGhg/10PX76UZiPwhVrRiTKvPu7wjH2qcgWLms3OCxkT2
ZrQb1eDbVafxEV1GwLD/FqkGigf+3ZFnb+GEroubjTMAfkJxpzCGrXBeiZy3DbXm4a8lmUD0t8qe
/+bnGOSPAKM50aYN8rJZWiZ/lSycpXHz0sMm4W5ZphPmM4b3+wIwfD3LmSWverN+pnl1U++fEmzl
X5DUQaxoFXNSLry15MC2EeXQ38/qtQ+Owosh4n4MsHnexVXYv8E7vu90CsoekgQyUet3WUJN/PiH
RimRfq3Y1m6Hq51yPtYjQ6PdOC6CSRV+zIOAP3vZhxm1/Ad+/phP/LDpfrjLJDhSMnrpt6gtcQtk
BiBcKhv1p1Jt1m8gijYtTXoiDvSexc6qBxSP1hp58AXiHa/Y3W1fcH231g6EfQg4s05ur1GC1ZQr
qbyX4pF7Dd3ape1ntbV5n/2bkQbTUfJr5isAhU2q1w2Abq+AFOtiwSGzSIqd+1D8f7MRuIe2nysv
kB7kf9ZFAWPnzu62g+Xzs/cIyUSyK8bXx5qZMKAg7C8p+/N7fLCDt+ZzKdzrl8KLc7OlfiZt87fZ
ZZ42/0sAxqjvo4BI5uV1t4wCh3u5+Vr6YTnv3DVuLOG9cmN0DfQoEk9/4PgZTmejTQ9ejGtC/Cbu
tcEOi6QtVcWEqzgQgPXOS8Df4xXPV50fYzN1no6N3F5jZFfxaqfjEOxJP9zWoDdrItkeBfrNZ6gH
u6tcbcM3iG6k4lzlbXKVXk2rGLpJK7oQByWkRAIgZUuj62iuEdc6XMQ4Nf3GQFIyYf+Mex3DzcKS
QwU3KlRP0kbExXsbZo/odUzhA4hgUK3le2HXKRJKA07/krBEIkBoAVUlzkbqC+AxbgMy82zPZMow
irFSUPGDu+ZLDeYpUIOIFFiMl+zqx3bwa2cPCy5CaKqzBABfetpspKQGr3P+F0FHG7jBtBdWYgDy
xqgB4wRURAvSV/0oqVEDgZYheWWTpDjsvHpO1QARzXXIcniDdoyyLZWK/nf2zglqT688ongcBe2d
fRI5694uZ/ec6H3S76u3xGPs7C8EFtczt/qqUGD8Ka1loQurLM+pGKA9vMMxxiMQ1eqwgsZQVp6Q
0MuU+ZqaZP/f6Mz39hnsgEMNsAclHTRj7xG7/Q3ETfipwlWsf7wkrfCtd/AVL4Ae/MR8uPzocZ61
PBcEmgc5D2UeDgZyXOH91eZQvQDlLexeD2L7MnzRyJH4ikfee6ezFs3dePY51D/Q9PABzW9+THuj
W+ebwBt+4OsTccrqCwPCGaa6RCM3mZzK7i+G0dLHse1ghIO9nL50UyUwQDF9Qd+N4ikKlD+N8MWA
c2qdLCU4pQYkZyTqXeVYvnLVoT15Akf67GUGRC2sbQ0OgnIvvBMrTz5otx56jtXTGK/QjGrl8Qnc
rs+WBchXpWCAmwmUmDWXobyn7/KE1zUg0pjvoxKdcY/Ls3IfjaLC+CQGviZYC/wPo6fRhRzLOBIC
FlWpvf43T5V4Y3aJYAjeyt4D+pJZjG1RbP4Q15dVdLmCvzvSWX14lupoG7VkkIk7RIrSHrPN/hwm
tHUBjBFH3HeTrWh9m0ULWIayr3goMB0tSR9xcBJWDCQlRFjy/Z1Y+vvRiVcoz9aPsH6PhIFjNBrN
RyCT/6HLp0RSfHlKf7NlPuIqjw1el1T8deCwzgWFWTuE+woub15kbL0284kP4aEh6AfH8Mh+39Di
dRdPFx3I+ITFnF9neL5i7CDOUjzAeF6GAg0zDCxYn/Q8DTxNw/fSGyy41KdzRhofLsdLOTzQZAq/
W8K40zUTiI6iR1gMqrsTWfBwMYsr6x+azApurqmxZCNymVj05EvIPrr71eNtmLNAlNaVxWRW/pNA
tkIEivdKwfEtaP17T7Zt8SsuP/e/Q4wmhZDcWtkTmpo+jizovHAaEhHgJwS9kAW6xL+QEqzA6oQ/
wr233dlJr3gde04a7JGHX/ASA6Kp3fb/A+qcO21MZSPkLCVckywowTYYwxOkZSGEac7TLYRzG1C3
itmkyK6OJ+8YU5lBOlU4e46fmhgL4/7QqyN2ID3E3qYc4aXsU4SvA71WcsCK3zfH1bYLcIdEoeUP
1hVvUSFRTiYzZ/maAoX4Q4eGeTh0AYDkyS1PCiDjmxWUpcCH/G5D8voYB38Kq45i2F9at52k7TDq
bpYmZKAiqdgXwfm0plTd5d1ihX3ivXtnj7ONYCKjrKQc3azlAOkOy5GKvCfDJXrFW7KvENw8l8bX
Q6lOdKOZ9dQbZjmDyoscBJar1CQD3YYMAveOUOwh5Jf2666T8l4aQYFFi8LQmDW/2ZQKXU3aZly5
G1z+SjUEd9mEC2n77v6rMXfwkOAXv8LWHCMsgX0EXGVoEihZru56fnNgrw8DilXw6lILoDXkQDKw
Y5bD0Czd7AFt1ccDMj434lDlyRgiCNHk2lYKVLKVFbsJt+0CXsaBMATeokFm1rC9bO5btPIQffI+
6LabMd1tZMpymTUQz0u8GKjI0ohHhgIB5taLru+hbWrxXxVXKNDXzPVnzYp0goHYHERHqZOzCh98
q9WVrbftc7DTQkA48TEBBwK21pGqCq7pRdlDj5wYsTy2JHVT07PW1ZcHzgRKWlxb/3tJ94AQqOni
3WrHFnX7C7h1+9+Q5hENstQfMBFcQhw20rU+Lq6gPph/8ojYbkbY0K4CXBpX/7chUUGXggQ0lQpO
sgOokmHHgSkaRu30UQnV1djoBl9rPAw1f8hrQJX904wJ/1ouofiK1YXAEVl1Yo/MyAPyQyqPjkuM
/BbR/NebCiZi4QLWGoUmxtwmtOXKhnnppiyee9KpDGJtVQ+Yw7D8QZbWGkhvUmOShRYhl1Pyv0ui
OgBuXyATlJBX5JmRua9aSzfr0qTY+G1uWlPxPa7TsrwNwojRqfVAhtmYus+P5u2R1NsPdGS9/P47
ODpPqfO/VuOMcLfRr9AO2GU/l4hXYRZSospvM78rK+mh6tn7sU89MtjlRYYR0Dj0e9GEJeKy8hNw
KlsFizFKAk0+iGeE5jmzIBxJrpEIKHbg4B8QzT5iPqj3egwPxmE2MI8BId2EV44qAXl8/c/rkqEB
j+ueETGeesz/YhOojc3rVNMDjSnXd+7BTgTXj0cOvCVGbjybPPy46oy0GwER1YpmNPDNW7aykfz4
yTlCTmTj3zqNyjm3dk7gW2+2wxEv+8repmfqU5sK5PTbN1QKEMAQsg1sZ/RC6PB2GY3rDEcRHYD+
z4s+Y6SKgUBoktHoEVeWGdXulA+x+VvAV260XxV+Xpco973rzmKy6oyF7Eai2gBXgEfnuotHCFtP
YdWH2w9R/QdiFwNQVXQ8u4mWxDjQSDgPVB+pHnqmHYhum9WUSKyPslkgCpa0JnSn/X/uY1/2evVI
g5p6hrU9pXHjexf97lNJ2j9wHU2kc2g46DY63lRwuj5g/SYwztLkAYISlmg4BaPKOf7tBUfqBrzZ
62C3MCDAJBPsQRUCRP6Oj7VFJDKECLJGSu3HbG5ZzLXKed/HeFz2nDmkwDg/KWMHvPGIfO4XXrQH
LBBEzrkwAvjXWScxxtVEUf8l1VEL5elMNJwZ2JPEv4wo+WFvaiA4rnoE7gXdQxp6teruJrRa748i
zzj+XQWJMoKiuO8OMj//QHyMhINkJGiyzJO2WUbdyifqzi/KVerikUvyqOr60bfYSV8ZbBL0ZVAP
1kEHqG5eEBFjWONsVNJ5k0vIU9licKyHvLtTHDe1zNEcaqe3SQh7cOCr/IZjLRgDkjLsehDyCCVQ
fgP7uigXRqGrimmTq521GVWTpBef4UMjWfUIJEWwOZ2zETIVE4VutLKyiVieUYTCSnsTBRparF1l
CWdNmYz3vJvPAa1qEINhg7MrhINITdbSrgyVBSaZGiV/c0ysJiYCq6cN41a/zeyNXPh8OYXPrNsq
hRX5mfGnZyCLChdtaAD8bqdSzYA1wuxty+z2L5+GNOtQRg9qh2QW8AAvz0gbg/7BbQutMbE/30sC
3O4lCUn2dqrj+yBEXe+wXLlQihACVwQULHaX7Y85K3zrieBWAbjJnkKZYkg/rBgijOJIUbhWDjO2
pi/Wixha8jXty+wC6qBRc97Usscelp0jMU3pzKFhjkYm1uyNHB7wEUgQyYuMrpkuwagLxtCY5Ofi
/Dqn8+eTHsIwCh61+VUlLwNvHPAZ7BYcdk/1WNCyVfmD2aNkfVKp5/1fTXXv71q4IMl+jRNy5fTL
xLzibW+9SllNktF4UsMMhvFqkgcy4g7IObEFOfmnbNDqbQkh9/PLrip04ok7/hxzFjbAXK++PVBu
cM1VWA0W8znqsi+zG6+w/3qOTaA9dgRnpztBXMq9uUaDjFk9lSdSrNpiuk4cru+kMEJLrA0MHB7l
Kxp0oCPfnvwjL3ZcDQjLfWVHUqumUBhB7dEIsG/LOXvwq6SDiTnIsgBKCVZvPg0ogVyW2Ki9ySFw
nyy1949/MXvRUyIhkSzTLajO0NRkWJ7/MnkgAHArHwXfG+UnZoZILPz3t57lsYSecelZYsjGcbf2
GyI9scXmyMhABhSgadYdbpsd1PTmgYVmjNGEmZcE5IKxdo8AlDeeXDVRSNq3NIoXRinJXhZJ0NAQ
XkHllCNSFs1A7UYUupz3meju2qqLi40no9GN8U165sgTi8FJekBMTKy8IVJeQXMXlMKDGJ1a9q4P
+tAOUPsMwlnNYiESS7T8hjWkGSfBLazItqz6SeCiTFWkPauFmubFS8MlqTBDLHalgrxbEbn9bI0R
pLMG5wu70VhYslnkMeMSTzKqfAwUbUCWmI8/T/GBowGOPY0zkEhB3Dsa66MlgfVuHKFNof15QNl6
4XLv0lkahyU0i/rJcY6qd9QYfqvk1T3dqGSS7j1p527MWoy/qZAH6/b8QNa8gu/g7QWMLc0zGRV3
2lzlfNDK8U0QZI29Got/MMt3zJtPVFhlVdqS9VXtTtAIXf6rfUgBs83fb6zACRCVeQ6rLPFazm+T
i4ZESZydVBbeRt9sr+yIvYIDmrdrKoYx+jEmd0OjGOPFaPkvUpIzw3qAYWzbDmgo4hhr7NmEEgPV
K4gNI22ti6XNinR4JQflNfvw0ZyozA7OnyT3+KcgrHBlfSIRe9QFtQLG33PudnSGSoIB3I500T6k
OfmkIvDBVJg/NU6O9nKXybZlcW58f/STSgLZ+6G9E5PU+0MZwyzNJMIucZtJbJLeBAkAGxs/b+N+
Ow+aVTWTRPY1zJixT52VjXpbzLCGje61Y8Pr9NeYSC8shTZ8G00oJAQ49/0EqcUMq8RxsClwe/iD
olSUNmWfDJOxSx8ZUviMH4AxBD0CfiAJAnOSHxu6Yuu4ZxJMOLR7i0hA/X2ESfk6Qaby4Z6/lOi9
3RKouAMLN0DGThV+8LpVByojzoiLIq2cH2IQPfnodH/CTo/Qt6CQ7fKgdqUqvWM/GNj5vBOAiBpD
gByILwRzILT+JlWqYx7XpArUW0mPATFw+cG9BjOCTlP4xRFzjnkkFtFmM5czECs6SDKx5bvHd0aB
C0atEXchtgU3i6vXUz51rup2p+kECJHtOGBH6uatfkVem7VMdduxprS8a1KiM0NGaAPVLC3riYzj
CuJf5VwYZk/b8cWuFJ6eIVySJAJUs1j4BKKKOwKdzruRndjoDXXnQ6820cGS6/EpcCbtFaRVIus7
uS3gmMJEF0qcBRrWJl4Oh6UZef07k4C1HqjPRf7f6RMG5z1IlPnNkIa4AA+WqKY5gUi00xqvylQi
Ljk3Ic6E+HeVyjVItlsFN2KnM/hU95hUplM3fVPHzSOcHAUSZgrP6YpjeBlH3BJB8GgWSYoUTktV
2NTtQmnte6A87jSUjC4oQPslIDAPc7UW2UKpOb48CrOdb9/6aMDi0O7xybNHJFF+uZNNmHz/YPGQ
ufgia9SsQ0pxgHEblM/aWGuWYnBhwTDv5CNGte0som9FZNdSX3hfHBcNfbfa04xvxJowrc6V3EBI
8Kgq3K0guu8+vgoxiCEk2pCMTSrnMX6oISlMhVU9vHExkCHvk4fcOaPIjlsygOIIMcgkM3zLu+8u
ZJRmtgyeWBmOh4LesgqXpYUF1yYiKdc2AG1nb13ErtUSoLI65WMAtAhDKQpoEYX/sYWiHn6Z7rLf
iYZRTy/RaiEie38oYzzCIBmAUOi79KNHZgK9+gf5L98fZ8zHSHMd6WkiL74uNK4q7MqL29b7F7mU
UPoLh0rCmMAwzJlAuCICRTNjSHYX1mPGpmfWmvnzOUC5RntdRkniO6NO2uo0PpC5x9hrYBeB0/ad
xjaYqLO5W6HCOiESExSUWdBLimYRwP2GGhW0DuUudv8Xi5FybGiarIRRh4yUl4kCFcynVGPJt/MB
OFIdjA/QYqO8sTGWA5t6JKhufsP/HkxQ3VK7nXior2MY0xUE7dr3Pn5rFTZpfmFaHh+IWnMY+sxM
h+TRw/mO21ZA7e7MuKr7lcJb1/ikXIjVvlHG+4p3ZGhTbkgi97ti/e60V0n2Vszw8EOdxOwrH6vo
BzWBubjaG05dz/YtHAtWlDrOzdzXvOBySfe1TyneFNMq54YhCqL/LNH94t+thyceMYcuxRDQqfZ4
wa6/7y5y0cumc2NCZk4IgWl6IinPeE3dBx+7NDhrFgH2xtraCv953RSTJbCjJ2uMmsBZX00whXHp
cvAjGhZauKrh2GJXzDx/DZSSkl6RxYS7z9uJ8uJCu0CekvlHSCN7n1VGMlmTXw8dcylk95hlsRae
qu1cLp4FtgLEXhotp1mPVxUqZGsckxsTupi9CKz5e+eZzZjlxwOtlJfhlMGWVPoCiou+HpfI0nK/
aA9+8DnScWjbiR6+7mPnufBCNp1/m0MTjvRyaSQUCPxNUxPQKklNlHC90SqIqacbafme4mNf7UlY
gmL26+rtBSW/eSbK6YS+XHNblh4PXeQhgWNvrDjevTmRn5N2w1zEcUyeUveGl0OFTjLZ3KAXDstT
Rt3z2n3cYNJt+1IAeIOQzSV3ga/oLU76PX3SFJrm+pTdAjWhR4aJ1BzZf7NuRlg9DuIWnRJorQ9t
ZA+1mE74DfRGyCC5x4ZuLPl3kd3lY3cZO8EuarMuForHHAMJqOMLJy452i/H934czBcLRmCgjSBk
mBTo68WHEeVXambVG4+VXJtdaOuMTk38YaF3fKntsj1KIrzoC2fEZ5tKiawXOVCAopytYIwD0UFa
CFVdqC017Mz5eKBtwnKB9rTONCyBOSSdEpKgL1gIWI0oWi3Z+gsQ7Gf648BQz0J+bEuZLzTqadsJ
LFfqwEq2sdVZRnfihznaTZ3G9g/qkR56Me6ImwN4gzPx1oENUGJUbin0NJuKHFAPvJ2/XG1n070W
9YHnuVplCLi5ffp2JxGDku80hLQ2IcMcMbazsy3E+z6lzo0BcLvNusqDOeZhT2dLtFZiAi/nUtil
+HPWCFp1ZLQTw+bqx/Ku8uFdsRb6d21M7ie7VWihpeBwGGy5RhnnaR9VHKxJeorHcwyW/DdiUf+0
0Dyhpgwg96R5EX/gDo1NzW8EZMmBBuO7NWQQIIIRM0SNd5/XOQAAtEgELtUAwQlj/J4YGCh2EKDd
7R6Hugz2qzQA5pJRGeFVR55BUZVNWhX6gnHxOaXKP7yW9vcStMc1FxtwHrKA2qpX70MszIOMTwl/
K8vqKJDApm1eS0jIsENk5S1RFOpcXYSyDwZ9xmbRDdZunQCQBw0YZdw8rSidKzaR7S8+i8TBn8L+
Om9QuimapZRmfNZ1c+Jr7vrQJ4Ej/H4dJFjkr7ZaWctVtxjuRrdKWye8q/vSiye98SA9yJVlP1ks
RzCbdfzSCLNLs9Mv2lQq+XAOgGEbjudcSO05r74OQammqf4IlRLEUdFV/bY7+jeZT1P+zXx7jVv+
jTRD9ZNRF1nx9jwxVlRoGPA6wtfdoCeDIaYT+G4j5aSj+zpf2Yo4+0kOo0T3h5Ek9D9tV5cyhbay
n5A/lSscMBjwfwXFUOx4qgDovc76RWVSbj+PinPeysVlpqX2WYutBHBVVjy4IOdgirKKqJV7BmWF
LsNKuHdPBoCam9SoGWQeXMn7RFvuHpMuL4+jov6evSKSrwqfxbLm1FX5l6xBO3VUOVscV+BwAtop
jdMqEVduXQk1fiSODT+9yOypgn39in6zpDQVdmk4/cTQf1zh+e9aJ17F8y22yTxvrGFTgydYvrpG
EZaD8HloAGLJmEdOhub8CGg9DcHrw7Tye2s+5eL0gr/TIF+ynukRkMiA5GDcxV+1SHEp6XZ9fzwO
AS1TmJAdkrwuOPkL2zKqziqJ1et1+4vHzO5+A64v6n73XUWiesjYNjm8YH+nVmv0PCMR70ysyKjk
qc3NU8ev1eRxd8+pnVvk0K1rY4+phPAY38lOeR+6lSQ0IkdGy985G2YTefEAfXBNfYGhyGT0aqBX
qJrhxGwG88sYXfaGsnl7R2VChwkMtbkvXZl9MXY9/xcvb7Q++VpzUvqc2eFnYO0PJ5cJXeyp/KC+
jS7+KKmpZEIJuxKBjINr+HMe/Z0ufDFldRi+3Bhs38TiskvDRBYcKTxDBHLA5z958TKvrwYBQcTn
XDvsWmQMrQqw4mIZHtaCz01VDu4wdn+5/YmFUPtYjoK+x6yfq0bn79tX5X5PJoAc9KzfMlsTQFDq
f5I4iJPQT7NkZpdn8E+wsPEFUAPDBytD3/msW7eYaDqL8fhCE6N/mVPK7zJ/O/HnUXKSkLVAQH8Z
3dEctduU7UYcjhORS4R30PGCfneVqpELt+2sgSb2WjvUqrYimEneS3xsNmY11OcMwY0PKFyLgrkQ
EuP1yzWcsewnWwPdj/MDv/v9BTDgeq5aQicJBMqKD7JZc6//fAkHLVRt5S8Z36r8qRjlcce6Jcko
t57s3pXCEETGX2KMC0CFpEulzUcw0W2o8uHqS5hFQhQo6NvS0YwUKAuv2Q6UgPAjLlOabOzJcISW
eOz8WPm6sm5pnypKiursP4K5phNeZL+SYue9WgwUYrrETNcQM8rZtU0/qydsgV//tIlR/gMLNTU4
t2Md/GKRJk6NpcSgDtJQ6cVlf0WmO++4c24MXQFgYihIio9CetzblnpNEBUK67eDXfPeiNDdnua3
67s7vZgKDxXYtUpVnlKYua4+4Q8nFi4/y11oDwcJfl2J0Kge3mW+Wnj6+UPqLYgKNFJzTa8/eiYT
2yMP+IvbG4ksFfdvgiVPX6cYEux4d9T6iY3QA7Wohc1mL8Nups6qTZpjOfO9vfJs4GOp1EdQn+uM
2B9Hn3GchROqyDCv+XNjmalpu4t141a/3B4Rvk1NacnXEf1JquGKcfeJoKJBAslyiVGlo4u3QESz
a/+SK+j1A/hzjUT4iiVZvuOhFWicfrR34uhOGgm9gpt2GahnHFa3fdkjdhSxugVEeSaFmy7nBF1G
X0vc3Vy97kjDQCZNad/pQTKqP2eKlgJ3CmfVoRCi5byl1sxhBFstZsc3FPYiWMUZ1hCxaPXgzJkM
5oQrTtJ8SbFACinzazcx+NXNwFGOS5fC3yUlnxy3mWzLZnAkljT2EU+KNx7+3P3g9D1FyM+ylfgp
DOZy0fdSTAlmuxY/hTgLfvVT8rcpRoDIjJNBbPFQvlTb7PhC5vuVFCkClhPdw+CJ5tkruTuGihe8
iVkLe6qj2+mbMqotMPnQ7XVhY7QdQU6XrciGLPMfVHEeXR7Z8m6D4M5E5ydpBKFejhNNmapABY3m
s1mwC/pNQAS9LZ/RsS8LCoUWcqX4bMd2q4wJo5Rmf0Aa0PvR4HKBL6yhZtD/oiu55cObdSeaVBf4
Ipxn9u2CjTtAPBvApnabtpgW1/n6gR96QQ0LGG7JEjfG1oKBGR/g7Kv07cyn3u+580m3kV/wdJoU
qH90nuKqKidRTTsQJvls3cBm+BDPK/VIPr0wrbIJbMSyptAUqsFmesl1RwQ9HZ5w/wGud8SE+DKX
9QC1FH8ZgyiXPxfwqV9fXO2n9m+AyjIzzJrZuhq6BM5bCwVz/sTgacJUO2ZYwpoQVoNjxe0CrO17
E3eN6KynHFiMe/a9lSu7JqzWPV2zOkYwwl+48RRG9l/JgpqU/rDzJj8ODfMqOouvLXJwALD3mdOw
7CEblt07vga+cZ5O9oDVB34y8EIwzi+kyAKwBA5WUjYEJ0VkphqUY016+/N0nfHcolNlv1jDMVX8
UqYEj06eS5dd4gnATWmM14++drrEDZR22DGeLp/daAfIZydE9huw587mFahU3tz4ZpA6CsOPHTj9
wuqfVUobf+XoBpmg4+PnWtnsvaySB6mbSYInmJfD6U8nQfImHSDKGImuMKs4oGrPMtnTIK0TdeiO
juF8cc49Ta69LSury94gBer0RAzezOm/awsuEeu8hjsbF0sB/xn03reJNYUt4053vFNd+ObVbNi4
PLwZZIUEJ2a5iaRglOdnAXVPwktUa59IbomWeuRnRqkBxzzG9eRnUz6XcQklDbD/+u9I2Pc8mdO2
Y6rmVnL5+LQLJ2EUJAOc3xfG/jOfuVKU7YaJ/DGShJs9+JbRnxxRmXvfAb/kXs+mVI2ZvYkDsIy3
3Za91h/Y05W1vsH1VUd3blBw28Kwa3dqd/eIsxPyF7BgWrKUcfCtc/kYA9t7EksOXtufedj9UAgI
alWQZNN44Mi3S1H7G76/EwYc4ou02uad4YQSiHNDjWl9E/+RMeR1cXEPkRh+PHswKw+6qt9Ba/PE
gU1d376xGYe0oe7FClkO0gJRUt2IdsrtelYPlmNr17CP1MW++77b8tPcBD9YOsG2JZ4D+uW+3JjV
KXnFT6t4FmA1TjAV38Bi85acbyYJKCtkuJ1/Miem3vfy/b05WQlkLsvFFuv9I4JMFmE6LXtfNWau
4OWiD3palnb1S2cyOZeKRxJ+kmV9eQXzRSwZWmwAJvkvoliykJQWSTxIADCQEp2JZk34XVJ8bq8D
HRzWcoYxBPqeEySpAtE6eZnnUFWp83IivNiT5J7v7THjJiPYgpyFo+RHp5/8VZiAaH/VN4I9zqfM
09UTsjjfC1nHdM6zj0HxqbmeaSPDuo6ywIRG7hxl3FED/6KHvVfuXMyxI4/+SEZEC1zYraAuHayO
nexMRXRs5LTALjlEnCSOWUgnEv/79qYV9woPZmLxuZ0fCg/59U+qP58BuoOgj8wFXPDY88Qic594
MtmdaJLcoJZMeBxYh+q17P4Cfu/5BudZvmGgmLir9HXDeGcIdg8c2AhgPy4MH9mJyBWvtLBaHnsO
EDex1b+MdOQXe7ODGSVAVuTxImq3G7iZHxqIB7aspoCWZYi4gbJrtHv+R5gvJZtmxkzG8/PQ04Vg
tsHIpbdCvPXmXRM77bnWI9zMce2qsA8lU1rkhiNDF6J2eqFKtYX0Kd9i5+cjXSz5aoA5qHwjNyiL
YVYHcyhlowcb6Fgecb+UMWJbPAWeAjPpkmBYezMee31+rOYCiBHbPe//Z89Y3bqEyt1QhDVo2R0k
oX33nfRl6OKNl9tCD/jyfjW44Ou+01ALQCqIXP+Aznnnv5R62I3AxGNUJA5N/VzXsjc4ixuWiUM6
gf2gscHIedwDR4wXljB9uIQUoDFdZ5wW4k++gLjJRgPYYXlcwDvSCRtfT50J7lm8O9f67VAa+92H
mZu5UhWj9R07JcFDwNhCeNOQ2o3puw7x1b98+QNch4V2kiTqx+CuO+j1ERsGee7xXDcpgKWf0PtN
zUfRKbKX1S70K2aW/Zy65/QqpxtXY+jrXdD6u3JuqTXVzGaK2lao/ZahfyRprZn24aBLJs1qI0qe
EddwkLGdnPH/GY0JLZZLsKnp0sXhK+LMYtwA80GC0Gg+uNaJ6aOKB8EIHq5WextQV/zoVqPQcfxf
2V216BEM2fxkcK5Sq7hkl0svlXTlE5F25GKVPJt5hhDL6MCs6SWzOyrbH4nO1HylxZvQktaBiEM+
8p/jHhmYj8XbIOMN3FE+GRQFOXSlK6BkgREPatllhmpZbW6qB1y3yl85KbEoEp8cAL4kOxwUh0Mn
fhM2IP4OhBz40kSL4URJOpIf+uEuxuygvI882KfI2OUL0NZfr3QKiBOK88/VMEdQYS7aAWCa44aW
l4XVMzsY5aMxzMA4eiaGRYjmYhivdA9j1+wzdjqnF/tEpq9TYAiILKwPbQ6/DzWhx9COzNDn9rnn
fRkgH8L9A1uTQvilfSJGXPhbEgxZtNcyUrL9FxRoXjsYNE5TkUYAeLeszSpUyLmkgPtMIem9oeoO
lZXe24RK8QvcEE8how7onScB1YCJRFFEAqpwmXJeqOB5Ku+L3QBWX8nG0k97hWNsuxHHEIwt6uL+
9pLoX6RLXXMM2CV4laA7V15hVuvUaiV289Diu7CkvpygX3uUBvylrxYtPN0+VXEgV65LPU+3qKKg
/51Pxk+S7Od8uYO23+f33P+ACK1FJPPw8IHT4w7B55w42tHo0BHJpSpVOqRvfp2D9S1/nI5f9h+S
Y/TDY2Sc6Dd33gO9coa61MfeAcWTdnl+M3GS5faBDZDaV+J5V2eNG/A/EvKBJe/rJoNdqrDHpv4T
ehsQq4cDtjH5H/wUSJi/WHoQXl1TjJ3oncT1alRLn6qwANwNejPEa6JUZHNr1iyutaExd0oDv9ot
z6vDM1ncVaW0WzfSe6pfUo4/wFkd7oa/8+uiFwAH+3fLdJQef6ZuSGFPe9QXkMyb4VTIB9az8CZY
F0uZIdJBn7Q/ZObb6woI6McOIR4ZltUb3nCIUAdMghvUQBK18v7odGGeQ3r7mb0yLBUFQr8+R8EH
iHzSVagvq9WyWRY6JpywJmk06bcm+DddX2faRs/iiTN9UDsul1S8uoM8uHv553wgjX1cTCiuXH64
QyBSkF5p4q7ByulI7ZscUWqtYAlswpBR36/b0onI8XqvU/BMdj2XYFjJacbF2qmBuD6FeyuDe0+S
Iq3SzFcHcl3y12OwK8nDT4VOhJ6JdACqx0n26aXz/vtYYxH57lLDd+5O7y2bDWHe7YA8znXstkFX
aavcNFIMfTFYP6XpHydERYh0n3aEgz15i4DMW54jHOquewwr/sxBLugHhryIeHTOlUc1lequ5F7j
DVyeUSVqLeoy5ZYTyTDIwF4KQbKuFitzzyxpBIiSeC2+vvHJuBRNzA4473fNtVNySDbVikYPpRC+
KD2fblwCJX46g/O1J9jGUcqM6gbrcftiCl6OMig3OvZcSwzvKoK8vwIOwkqC91rkewEMo6EayL7v
/FFPHFbX4K6N4YCFZkM6AihB65QbqdLVORBxWSjJzqCIlIbBE4IlwRU6taqiwE86QUISBD/tyttr
pK9jXv5K77uwPRZUonljZH3CIXMnhsWRqO2PbSI/jgBxvsvr240VpLtZpWFAlZXOSSUrdPApLVWW
t9+3hQwqc8qT/ib5O2Y8TZ+N4REHLPuJRQ6O6nmnEd7dHWp4aEObU0HfttN+Q4lN/Yr2yrjeEkJg
iJ6oD3RaRfBx3NqOEtpFqXNcE8T9VlEyQENFP7q8mFQYxGErl6pv53sG2fPN7i4pJgtWzhEoM9qm
ohFmU853fk5UcjrXOYLvclPQuCO47vgTUQOFITaRD3H6+ruTDBx4ZuOHGQLa9ee2sRxg0vhf8A75
Ca04FhzcHfLBwNcGzsDRtMEIl8kmPJN+CT5mdopSL1rW3z9kLSYi9FLM+UI3JuMIbwupjrbD5el1
18v/mFKiUAXY8vdtplK2uzHpiKhSCFbxWspdL2BEa/2E7VttycjWyZaq4p5Zwkhf1B4W9XmJ1KA3
6pex1wBlEmxY6kG7lkq9Hwuyc9hB3o7YTDFlZWRkwHp1YZkdge/T3voCF6zDveIpCr39X9tGB5xH
DIB2zmSdqLQngCo37OFs0QdnsmOE0vJDlGAN+fBLmloykP2JwKnUsW7Le2+yK3hJBA1p4A1pOymI
a5b2flurUv63qNjFAjkrnBv2LMVic/i4zQ5MwFt33fecN94QWTBPLXtQj490LlmYGkaiDS/vyban
W9xzVwm4TTWkMUwQjEUQMaD1VPsdZCVWCyUQZqRKWpv9lCAwV9wMXqid0OIRf94FV94TobduIEIV
AKXtN0FBvwzyoyEaoehMH8bXybLAFX1G/e5CYlHjrQJqqWGI0fX7OwiYEY/hIBSdHkL2bJnsBOcW
ub+vSawui4LK7TAfMUbW4vDfIOjduoqKjoPtZ4QmSvx72Sv5SsfOVf+5MdbcVbPzKF/kbw6x6jVs
neeZfTP3yTYHeANpA5wpvvNMU6L9tfm7AAP6ucZCBp4GEUOvUGs0TCJjMlxwhI44dJRjHUadW+4O
r7HShgz5rNIHQNK088ZBuijP8Dw7PztbqVh7MczmI8wdgfB5QqFBCJc+m0UGg0yfo23/2s5PT1g5
wzWzW0A/BBXXPKX9ZaqtTeg1azr9WXm0Mxsj/mh0HIzRMAodTRU2/tQ/eyn/4qN18LvkfVtntUfu
pvnMcDjH3UFk1H2jCfRKTDVRHqSBLdhjgpsKstHcgHW1bNXA3r3CNNwVP4Cab0Cd7hljia1GsaMH
brXxCe3QQ4rQtUP2NA1kN0QcpoyK1t9OEn5adpvvypQabT9d5WJYJ+nXUdrx8mQ3DGktlD1GKFk4
Cf5W4dc4zqgRgbQxhalRzFR951D6+qXQOKpVIODQxBkao37X19VQntms6uKZ65kW54SJatrOySOs
VVR382fjc2E8KpgQHvfeklwZkdmlbKS5uRQqDAZliUlzqRvvyJJNSwVI2EXGOIyPlrVF+/8uvkce
K17krjimbLjQwZOeteVxfFk/MkTsOUxFORMlxLf0RPsGCvMCjLfWXdhmvY2ApXao5pOjnXJH90O2
rgcAKoQGlYRm5mgw8zQHw/vfgA5lxXFfB+acTWvVK6dxoIgNs9uDhdEyb7V2yjLUwYKJoYCuHtfq
KjwP4Q7N0rFX3Roj6jzwSabyz5HkNdBMH/VQzPF7AbeB9WQppG9lRsJmhG4vFngjZTGhQcD3A+S4
G23tA64llbeG0h99VGwTFIPIKdnh8SF+WG4iEfCWKQRvyRCYPmdXFWDuky5ORog0WZWyt8Bs0FhS
S5a2OmR8fXMI7aWrex885fC2ggjfZ7cTt8O+lW8SQOLZguu0h9cmFAK0SI74ffU0N3p1DZvyMYFw
Xa0bj1Mb9gAos5bMVlKSQvRmKAcTKAXtbDQXowKdjVVJqPs4V6vZKvL2371shDLT2LqwLXMwjH5x
50HuSehaJF8DqYKP/yd2rzRBYnKPp3yzaJkOY8SfDztVA5/wh0ZbMkTh9da/DnRr24nMgeqIMwMt
l+LlZyX8d50ZR2xMY7/zHdCQwqpEaYWUtrZ7d4ZwHwleql3vPo+AhIfph5b0LPJYFnjwSoYYrTlI
7ujQBpgDqrQm18bXMTutco/MEFAOhBhg0rPZdyGKqXL00gfivw33Q2bBiKIOq2+Du5C6+dW6Rlmk
241fb9JKw/klRhCE4lu0z9QtZ8ervFTkNSTN8pR+8samU1K8N/85GPK4/7mdD0NNDx5Q68XaL87x
AHKGbvfmgm/UeC3DghEDfGx8xycuS4uSeFrl37c04VhSNb9JW+PtGjlMj8gE6YHKpFXHQapSozoD
DZFTPrWv9yQvmeRKh3WPlLESN+2q2GXDAJNg18om2vUaphcShs2ODMphZSTbveUV4R8YgnD1bNFl
Tj+SBqe107QXb4gQa3r/M+kCC54NFPq11POg4Tkc1G1xGSgjjPIca396UNIzlEpnargmWsapz9qx
P7aLDsn+zJ83UweuT+1AbcrbN0NFQidC1QZJBk+LL6TmVAse3EH3JIg4Xn/i5i/CrL3/W93xS4rd
PwzO+1x0lUGocZbKg/9qwXZqp5UV81ILzY69NKS0zsx2deDLiW5AWYx+sdtVdpYq++a3/PyJv5z8
i4YIArGMAdRBp2zopHYie+XbelumBS2og0czBawiXGL6AbyfyOBr2IwtFmMdIyBB6U2x/yqraq78
KN0pwxnBa6yM7ScjxM/3CMAoTBSIgdXzodbdQO/JV35heveiX5QXJY3gTdaedwGp1yoeJdN0hJ9c
fqDByWFCbe1ZNiO2SFH0RUgCqj6fvE8C3qKiKcVJSzY4pFXkgN8JpmUoPH7tipN7CocYrVtmP81p
GcMkVNTiTF+zWEV0Y75ctDDhHfcbZDMKu5tAvj3cfUfZTunJbNqpUz4npSPJ4mDJL3wCRDKKABYS
HiU6iXx9P2IKeACWwIVw3suhlmKdtbZDVOI1v16LTHY0tetSgma/qeqEU435TnJcZ4vgpV2dXgsS
izWWRdjWKj2HhP61Zig+1PJmJOf31DbucxBvNEilzpMI9ZmM+tEkP3Ogu+P4M47NIgTCgo82QYfx
5BGvNDJYVLgSJNJUYFpEOHfk6HbzRSMgUg5HdC+I4c3yJrArIEPTr9OKT/ATArxBuQmnMHukh13v
aj3cGAOcjvC23rdRjh5HgcsRoYKyPHkVsybqjTHXumIbhzX8VxtK7ujCVVEn0brAMIG58j2iGOyk
uaxAsmAHDjhxASPbvdBDetssh3Gny7or44IkDQkIFmt0Opf1BIuU0D5kA041frUXqLfwh5ah8Wwj
RaEiUG8J5wD041eSlhVGUQLxAFccExI2tbFGnwBnJiztrszUoYBhEE79E4MY7RYa29DFvh4jzuKX
Kof4E5uD9sNdVuOaWItaXEvR3Ma7jzIcfiIv53M+8BhJQGDNotUuj3rnpRUzr69m94aQqayssbkI
2Uts4HzurJDNebeWD79282iDjkKqMMW/++GzSWUIivq4zqYqSNYV8176XJzoW1ow2adgRpvWCrW2
ccQLj+NGoWbcFVOohdlaUC9wAMT15I8M/fy4nDo0LHV9rWrlCZJeW2WrQsltjm2/YejbMOiIFTby
Qi9gcgAbkz1TpPwClz0q9Yi5sKz9fsBS0+v/ZLnnxn3k5HRPnr4Ru/cNc1+qawlBqxqvThKb2HcP
1MVQ/PTK6MeqyiZTuFlHwEsGhD6Lay6tMXHFXaz0q6YhZ0jUulpt9JLa4SLyjmW+0ItutydOoOxA
EdBeOlyJEWmK/btLrKpoYP52sxy+nNdnHqwa7UTaM96IXGGrDpU+i3LyDMA9xnCZEC4WKAAxiZA0
Rvhx2EYYX98L3m7ciWqQ2FGwQu3Zx9FMR6hsULuTFwHTLDzVfLll1WZ26Plltn9puUtwmTctIkZg
iGIUvzXtAhdXVwSHB0PN6WK+Wj4SvXzB1SNeyRiz1stoBl+WmvPUFjLMIq7bkmEyv3OrP2NLNCZ6
UvBFV3FYRQGoi23hAqhMgU9oT5MrmqM5vfxrOm/08do5YlJrfsopKWcXPtsxIyCoecqbdEnfCk6Y
xOH5c/Ly7dQdmhhLg+GtX699NvHkuka0Tv7w1YAAkvALDarlOWTAgibPnj70T4gfSJEd2qC9wGjw
/CnEsjF6b/hJcelBe238XwVAQRzK1q+xtDkU85PK16VwEjNQDXTMOCiQ7PepTaFDA+Sk20z73jA9
Acqqa6SxbIaUXPUsN/qJokgftqlktq4a/Tx04gj1uuUhacOJTHiFCda4h9a6chfS6tJrRE1zYbQu
jzLMTvuytuqjejgxnrPYnYAvSHqnbA/6IQZ9O0OOfuVDjkH2ixOc8+vA5u/me52wtH6f4g63x5Yq
b5Ty31vUc9uF6s8LmxtYTCDCUxu5oVDBwmdq5n3q/7Ost0QYwYIfweLdcIe286RBYyUuyKI+7/qv
dchGzgf23pEp0IG0rl4xboXowQytpHYAJXICW17bwDuWYRZ5C189rWsg4SX6qapdlWFLhjPOTn4j
mOOaciDMcnOeahJUF1xWBK2rqy87Wz9ztpQRlQdWWs6EdJKmxWjD52/m5rdE3XbA0eutyOZc+Hf3
1Rkmmpgx7GwzMgQfTzHsjtbtaPvOoYF9hwDgi4QpxZceemv+S/2bsWCJexQcj+sZ4evBLR5AsRbB
engGKYqUyx690bsgbBA0K+F5P3uEdbgjy8/zMr2NZuXxOIqpH3iSZ91b6yz3XNsmT+yUzty2yWfw
3V0t9mmUCR0lGVz6gmeBMDx8ysL+eGAwU1rg+9D0w9EbHXB0NaGjk0W5y9wO3BD8CDDV0MCtiFIl
VcktJCBEuiTdyj4HzGijPE6vrNXK+2+U5OmjBFMlvdXRlWHj8fO7kbsR1mwuA3p7S0EN2s6Qpzvc
GCck98EZRRsrU0oCj1CYEihPCvXS4r7gSWhotqnJ3QlOvb85RbAejy0ep9R3N7XCh0G8kiVCE6w1
rg6V16aHeiUncQQy1u1OFuGb4bXoNLQQyLCJh29SREmG/f/ufGu34NGXd6EI5L4QNxOgX2ygoC9i
PMZad2peiRXLHUwgnFaH4G19DWZKmIlMWTGW346lx/uT5zs/ITbXaDgvd2d5P33xwes/urrL//iF
AtfgnIf/ycqH9j2zdnmeaWCnFMmEqcLtQzjnZTRjLMB/UjmiOTIWRjCZuZiUTsRGu4o79Wusy6XL
qwi0EeHS5g07cYb5vMztlT6fwIPG4JpHlrX85bAkez3/+K/yuO0XPHLZk/UACdr+qGdws6oGd0Yf
/mR0fpk12U3YvzjnMphDeLT/KXDNvaTsK398jJrRNvsv+6SfX0e3vSZc5ZoYdvHZ2nKyBD4BO/GH
fAvP1AZumdoZz7+RwfHX6pwOOjeb2RQQMVhdggeCrS+EsTdq2KQqJTAFkNWWjguYK6d7jhQolP4B
d6RjMkjmvqvILtU6g/2XjpwB+dZSJuLTOsUKjbZAzQJPGv1sg26eDOLNqwI95UKp/+ciLN998FFi
/g3sYqoTlTyfEGwO5GQrzze3RZ7FZXPOxlqHX0E66t26ezxWR3GbfQRUa25DLhGGf16c7d7zi97Q
LHJPbYgcq0ioj3lXcdXsHX0RVMITqE161TWYuK9l9/C/HUBb4JU+L7kUnIKSzJUPBKKngW5TNzGC
O+AkWkTJTIY/z1hOiUZyKb1oD+BQyBavGc1fv3ds0TVRSW6XOF4ojES5Gboen3/aHmiiOZY6VFI/
HChB9lSABwbtFuMLRwa3/qzm3ZfvPHY6FyuBCDr2b+i5L5egWFEzDGIPG9P1un+vRzbvmZciZXTk
xhbwbsThQmFXhemlk4FQvwM1m+2+eRZKmZ05Jeqhe4aG4OmuhTtLgXna4FhwWojc4J7IEIzMotsA
rm3qlXT27JwZ2+BM0VNA6PFCCJAsA6lQQPK/PpwbKWdiPozoadeLAK/5aPbG5KXnG+l40dZMxdcR
fsXCTBSMficCgNI3RkExmOx4TRF6TeFXMuXaBJFWnoiRaPVLeYtKq1T8jsCx5bAbJJaK1N92zLg7
W9FlKLr5UKHC4kOPoh1fDX6mgdPgHnzv3kH8MjGJOgtGJIRwNHTVR6pY5fIwx5jXG1wkVKt9ssZu
mJiVpITBFjjCUvjGfFrk8nxjBAC2O8WESKl6IwAqqyviDYkaQK4w6i4rX6bYBb7K9Nf1oSSXQUy6
0dFQ1nzg1vLJDVn9VL9MA7xr35bkTO78AS6jS3yf4OusrXCOb/Mlv6Ruw1NOAk3WJdw3leEgDsUJ
BopTp0f+24HLiPZWeCYpjfi1nHu7ulcsw4NSO9KBsgArxUp3/CS/3T4aMB+O1wtDSaFqjzYkCBTH
eYVTSK1wLxnYmWhPZstUP2rXl8psicxsEfWINQSC6q/BfvCBz6BbP4/VOoUlREedlFOZklfHpFq5
cR8XVebGC1V1UoIsj5kK0Hv403wnPYTlTzzW2Xcby6KiW71ebOoBTmx6DhdtIvUUmnfgE4oWmHe0
H6FWOhtj9aTTFKlIfI5cgb6nlbE1y/dPzORrYXHDpQfkF1eSChozciIWizQvka1CxG4lAps0uSb1
s4YtJN9GLgCfSxU+JCLvbr0UgRDiGSSmmoreXT01eG335+kfHgUuW0silOtfYYJa+XTvID1DtMmp
e7n+/+pNoVOfHPwf7zmfuYx4/ddd0Vm/nbdZiBrJLwBwVh9k1eMczsz3G5yb66x8M81s+BHW4z9a
HHHDbEjT7dcmSmMjPcNpbDgqX1N3cR5IaOqe8tQolenZ4wdj3s5SPNVNXd8zEvy1x5wKHjxMumxa
tua58PpDLbiAkomnq99nOKu39/Amg7xf1eskw/t/VeYP93mKLaYf8cwl/nnja9pH9rpsAtJz7QcR
bUhYIjSKMZDNXYG6ivR2MXGimRSnCamA/fwYqkMNHFl2/Kqgt0caCWGwbIkFVzC/PkF9KNj02Id4
JnmZKxRDAzW1YLms7hOeiFyMipJZ8KrwUaEzT3mPEhxvFQNhHPquwgaWQDh0z4IKbGUK+iOtXEdn
bJrb6t1ftZpCJvZRPmHULaERNWqaI8frxHodnan3uc1hTpi5j2UJmUpblllKjTk0lJw9+uAFmAy5
g3wATJOrjp/ctF2cjHvSR5jsnBMVo+gaxy3sZFPykKvteV/NKICs0EMFgzMP0Ki1kmB5kroEwZ6u
8AOWmNAfPaoeRtzHKpGavMnX63n8A1q8UwO3OrCMN86gMEfdQIm2ngi/TJNdJbxDFolphvPHEjIL
Z8kshvjaZJIEhmQU5E5Eg+tZtd1TmcEeLzhgQAdnys65nE5lJu4Jucvo5WM5wbYJ99mDb2+Kfjtv
qSg250A65Hp77YRCSTCWfAg2oYcgE19SNpx5PJshO8hVA45S8EpiXHuxyAaj9o3GMlVwl0hOcbsl
VtrCArs5x+AIOJ09DaKRZjlV9kdfeuh8Y3DT4sz80JKjkyG1OhNbAYrv67LgiLWYOLw4RWSYBNOY
OxBlfPbwnePWkobmIrJrGhBhBurRjT3W1/RgQ0qZGrEkV8vcthEs+Dk4Y9mAqFkY838jlFIgd/Ct
J3a/98WhW4sIJOSjYSb0dWesVyMjxDYB1K+QWJPAdWJpgTlpK8N/PyReOe0lPpKNCocvIWJ7ONKT
mdhtwtenFiQl6yoJKZ6fgUl7VL0tCiZxoNJ/+IF2vTPGwHCOs0J0JawpbzMZMlJMrIPBcycFZdh9
H3HM5ky6QyP4uusfEU9rnSUUqJHXHFJSLL4RKTsvd94urDSuFNbO4jaFqMybAVpKgG4bx0LsBGgX
+kHCb7Z8TZDxDZaWhjvlPO9HYJsTFvgk8xB3MZSQcn5XJtkNiSrdtHsITSX/O9tUOttAO0fE5RAA
lb6tHHD2a/WMD0D9zgeE9w2fkDDAwLBym/IWb7om5OLFdD4XOzPgVviKA1wVM/7jY+91GhTKLze5
f34pAZaqghrF9Cm+CDWEadZTLkMS44stl3/iBAxg3UYmh45E0690eFByMC6n/w7fU4WeFNW9PI1L
hNND3g3CGgBPURbCVOF1RPvd8i67zRXqHxWOhnLzN2vu7pBICljmnqcn2x1EKQipVlM6iu5YonAe
7dx9ng8ykzgavHZfiqVkRZfceOn9ldjqPK8fFsAXuL5tglCFrg7pLV4uewWL0kYHJXiOaLQJcc3W
FicAdQZwqaVWZDhBiHdmH1U4+RBhHI540zJMN3Ie53KwbEYSGmSTmqcm1FIFU9IOt4WCXrnjJxnQ
tUaSS7T4nICI5IOvD7fP/u/VPsEZv8TsT9Kzuo12l1fJ3FD8fGjmTdAVRQozWzctGw4mwhDBJOkb
fS32rjqgpq38B9UlK2+3WNaJ+dUYH7il5MGCZXSBfi7rNaVgT+DKuZ2k69tLyrDUGdo90DDSJNQ7
72BT8bsLkZaFpnPaJ84KFmT5bp4ptxNCI+ffX5lbes8Mv1aYFZUPIPOWpORhktnU4a5xDMUpCoiu
kEst8RsdK87Bio0QOaA1jd8UsqzNpDjx1QJArSHfkYv8s7GH7gwaodnEV3E2kuxNNP2D1PoKVWyS
1VZY+76k3RgFG/GTiaJBBLo+LnN737ndcStzq+ASDfk8Ix9Y4O6mObZ2kq0TD+sGt3k2H90x1rX6
2uEAwzdBmaDrEv7JBw9Us2xNrgSKq+hfhTdMz1Y5OMNI8fcVEXvMHOx7kah44jA1U1QI7Mjnczs7
3bMcHWVmKi4v4dREabuA6jONFlYlPzN3R/Ab3b2xM1W7cxG3Lvcc6adgVYxkaWNSl1IHF/UuFPER
ixf066JHWmsefsC4/w6z3JwN4QpEcb0u/R/lIm5iCYxml8IeXDnHd3e7nraTnmfMfw6R3WREblZG
x1Zeew4csI1igOkLOjYx923MKPVlc1BPy4Nh1ReOkLc85wkXi+zchaG30XcXKkRBScheTKDozXwU
WUJovnU+hAej6KJ5P7rB0Yf6KVnSYQHdsu+aoG+tq9AoX7E1HkeBGYKhoOyfCrMeuPRHvpcuo0ns
+I4KIsMK/0YOqLxD3SU9VGWbdFKjXN1ABZVmLrNC0QJ3U3HOmvyiCq31+rShuRqjMu1eOwTQKPEy
c6EhNIlzDy620Jnb8lVcdph7DQOG5qdErJrIP2jIbQYa6OypL8ggZogkdNBJVfXTVGpwMg8Ia+jT
TbgghyhXJUTyQ6MXO1WUZtNCEZWb1RcpDSTBDh0G3r3kxevCPBw3B+3AnrT8uXOMSONgWDEmYP6U
5r7yToLMz25FEJzqhamCEqQhmBIwZDGK2a8272uBCuhKqYNfj1gik0kQJDAyd+rKd4jrw6xxgDZZ
opAsxFe/yCCTksJtO3NRtiGFEXT39NsN+V1Pyu3SarlJEoN/PnOmTuzlxeabz0elsMwYuTf0Gi6P
QzHGiCeXNXgYfrN7/5hDTNSK45+jSrZ1r4sxduNILSoJm9GKcIgH0X2JFMdbAcWgVcytcBfDQHp7
otd8e1xMvj01Mh+Up0/bXm61OXUd+H28MciwBDOUEfFtHGxxMthLds/z4Uc8wCpvrbW9XlunF99P
E3I3M4mDrMs5ttwWERYZMqwzoYPqCvWohrCjwnIHTO9w9xrFyByfdD8xc/EakwyNdz2YU3/Mo3t3
0ypC2OfMuZIFUPMC6o0H6jdBxzih634GPU/InSBpBZH6u/vBlDFOlWFiZv6i1DGgz/SEBOKRQoZg
iR+4qvC7I7Zk5w+h3XfZPW6PF7btLxWz8NkTFAzpmIbQp5Md6fbq/xrD00aVvc8m8DtRVe7D0Bpl
6UUon8jkrx8wt5FJCGdRHTtyb3p/fnRKrJmhAyLGQgux3vojWB645TW3WRfEag2i3EmFvvcjoUiq
lIp4818Zip1HJYictvMtjPFL5V+6Mzr2IhCZC9LOZm5eA1eRi9m2WL83K/b/xxK99VsZ4jORC1pr
knxxgwyCm6J0EmFfK2q2e5rw20FIcCiD1EWovKePXCAz9XnP8YUAWqeUWOCqabkzTWT/Gnii2ERE
FXPuDcfjFGqZpD0CRY7CSskF21giUFLdZYifyLNBgNNmsNY5dcC1YX/Xriv3HVbnnt1gtHPYuDok
L/fX6oJM5TjcsxqAS8XThCJGMHm4JwIKZp6UcWxDTUuNnVENTt/s82IrCxtFefXJ6qeZnGvWf7bT
Q0GOfsj6x7huNqGoTEztnojPcP91p90YTYuhTDySJGs3jX3sMakl4iMworS35mQQYDlmKhLBKS5E
9gXH6wO8fmobqLeJjRbtvxdrfeiioDHOS+4YyVz4XmtlKU6GrC4Jv+brlqupNbzltAXvb84DX6m5
kdpTV47p+FVqdEWsQOH+LmK2gWNqsY5IMvL0UWPQUP9W0KUnm24fgtPqpQaKNGYQNxpWXihpvP1Y
KzmH7dl1uea3SHIilynXatLj2Lm6U4n+g2w7w8tSH/A6qIQG15ZWURXCqMQhPF0yzdTXs5nSPDXC
BP2DyDhlr0Xh0XGNQ+OyMGyTTbcWWb/HTTwma4DIxFAcpPq/nyB1uzEqaFnNEdU68nuPJhX6rLXi
oNTtmLMSVS/X7cjyBIxLX8+gL7yRlAGRAgaVfHpvc5wa1GIocIE3+g1Bc2nhBuHU4R+xO8J1u7QM
haB60PRHk5dTkw3UHvbReBTQpXFgNvT8XfEGrapuTebpFvBgpbDM8i40GwWgtjIQheUZfX61kZDw
ZL148q/EfXrQ1hLKrKfu8jiwWoU8ZqqrTEJZOKd79xGfFonx1gnGIvgizvj1lpItRNLX0CrwsYoS
OodFHsftjA6fT2GWdkRZjdyG+ywY6fBcVNdallQhvjOCEiKZoFV7W2VaNcdPPMgdJuEcbxCbYSqE
+gFyEid0+4jF2ndX5oZu51cF48IdC5UVUrhPHudymtxD0FEqGczb7n/GMGNjTLsnGhKKyi3gAh1+
kCbttUddg1zMbxqf3WXOkHkIUENpSVUsSiMwDb4AhiNziZbv1TF96VL11kvvXlLsO7xSVXK3HNiE
7W3xb9oa+FBNSFxA/9xNWvKv9nfEU8ijPu777+sN/i7BmYiEICU+u88zVBH1FulWY7aoUS6DFWuX
KDWdhdzSIDBUmZf6Ak2XAKVpdCH8QgUE+SRR2qyVVs68eEeqPBNpXM+HGT1P9dYSDrdFrh0KYaR3
/YKDUtqw4erPd9r7mPtDI27WXPo3wH3R27N53oWC1ADBg6GefJysAhhyitrhrr2eYPwObGJC+ugI
thtyErO9Q5yRSK/NRqQOoBqmKxjzlCfKwOgFplU8Ff8Rwja9YQnrtbRl5LhObMD/8nHbEgEgFfBa
iBTVQVVjONIqNsr1daBeHXZZoNBrvxsmJhwPKoDY7OausPXgGZgTwBbd+P9tucFPNpw6DbrIeC2Q
NUKfARxTLAxX7FBRcKlYqzUZDqk5yJW4H/RCLznqRpp4t/CZtR8aVUWvgZOftqHqU4LJw3ilnMXV
dQRV20rOlDENHHBRSxMR/zD0e/kttpZLklFAVCORWFcYG5GRWK5magQEJJN5m623QbBSpcp/Uhxd
oIS9QjMUfTkJprJpNw81WgceyE7FCE5Oyw2AN3yBiQSDGzQGHYwAEqPEaRcGuj+XFK6B3DNF7SiQ
CqSvjpu8sQf/ZnDTC2WIUVbTBEYi4m4bZ4RrTfYNZCWGyfvkcOGaEye8TnzZIGQO8Xpeys9lqUfl
6p/qa3xK9ZSch7ryQwVGVUqQEIk1TLPiK9KFZmGg8+Q3so18yn66lIGieXO/6nDW8eiuQkVkL/J5
ebF2sjAdzfBjh5uvECgZn0IJUoxZHEum6Hi8u0Hpo18hZagOC/YYkmv0PpOeZnKFj17ox++5s6Wo
Xc1MQG/juQ+PV8eGBpt8TP9gCWsm+Q6+4sIaztGLbG3i+Ql8kyYTz04ux0kWaiIIN7lwQpXHgJIl
VLdSL1ScWYy5UJPxtZlzvNKnbxx6HKNqyx1gMA1XTebEdKZ2VpOJ0u6lSJzQG679VH1T4Kn0lGNG
8NMJLagxUw8XslGdbSshC6TOUU9dMiOASBPEjRiZ6KUJP16wVkg8bJm526baw1Rv7IPjFKP3LfSl
p0F1qbtxbx1Qvh9i3RsbRqgxTcqMGgH0rDKTh2rKVHA9t5NezUzp9j18aV4xxJ1dupIm/H8hN1nT
v7uADOG9OGeuxPyLDde9CH/KVYaMUc+xhRwzMJ+sk9jHPeuFGv8TjqiPGVbGPKb4ZFuVSVx4wC2r
7Ohseh2fEBb/kSeuB4ygqMBydT74OpKSk/RSCZesPSJF4jfbIdEFrU+7o8XQSdlJZSjFGViVPcGl
9iUhv6nNwLkKuuUWu/9uATeEkYYB/Oj7wrXxegnFOwqHuzg+6BfPEa4x2W6WXMeuojIvak6gENec
iI1SYixnJBZigGT3L2WBKN7OoqAsGYZY2AfkjxlukHbNwUy6lYQqKMzu3C5FNoGHsqQel+mEhTWr
j/+2XUYT4ubz8Rh6cEyrWAEYEq8Jh+RauLlwqLraXP/RWiTGDLmHGbCbzuF9PVFgD3OlQRZ1oc4A
q6XdSijSjriF7z29KkoSEznGgOLm5TceRXEb+Hw9fpnxHjOF/SSnlyXhx3yYN9SQ6Nb00X3AD/fH
xIDCLtHu/AR2+RmdQy0TzJGoMHxeK1WqEyOcJYRvNhIW+cKv9JSqjnYjW4Z0pRGSUsk0eJgcHNy4
NvOeqkzuut+32Mwv9+LubDVCPMEL6QFG4WywZ/I9iSyqnNsca+zqJNMMphtH31KF3KU4T+9WNFyM
bcH/xct7ISQQXfx6hZ28zayxojzujFx+XeIxK3Giak5OJsgq1tN2hF6FN7IfEOvdA579N6Fgbi8/
fBk2PbI60WMSkb6uur+qAUrrwDvlhjSp1HOpJkSU6+aQWTwkwH/ZdCr9mPFEmlPMGb1qzl23apKT
WEUAugHBbTXM5va+YNbquRV8cVnPxgwG03fcCVNGQDAPmdlrVshxX7dxH4ldUk9znOHv7RpMGs6Q
l3wjKj1WJ93qMeI6kcWAL08kq9MtKQ5s71dGTln/1RionzLjgtq7iRfO0ucg+yte1S1uDgqgqADS
9hUupFxzJfLi90XAJ2HIZrzUUpFuJjv65TgyTzezP8l1cYmlKIhv+tZz2wrAgYQ1jvM6091itPLv
OACJVqoezfJY4qiFVBZs/w7f/TEcqmmDyWzRA0xVTtFzPEmUQxvfcL68lljX9kV3/6YMdxY6Zy2Q
6QVRCWxoDfC9g7tGcZbj2QSQyD4QaDLzt1RzhDHXTUyrdMchhutbmqHAp3rMVux4Gzt+U5n9SwJC
0ij8W5qv6fgWhUe2v6VKqsSJGLfxAAdXpYadzQiY3GrSMnbfLlIcCkF3Q4p9wUBIHAtH3cz5E0y6
GEwZWIk2CdeIh0IEYknF+OkOPK+R95f4eU8EhNVar7hFCMlHGjkWntGKL0hghlKFIFVyYbmUY9Jd
Hzry7Hqs5uFNe/rw3bjQa3sVAEa/+wOfhs9Tx6z2UTwxEJjcO+ZetwqSiP4FCQFyDxJIINRi7qoZ
Yj7HXVboGZZZh5qd+knTM6CE46QndBa06JWoIJcTyMovggQIA934w66dd7Fetxy1tJKfxl5JzzxF
zO23RJ2hXJz/gIgBul9/VJvAAdq3XsrW544nFgrCGUJmL+BXHUqTdJK9B7WduETIhLezSmuaLAlA
aAVUxdRHUhBuR2ou1t43+waY01Z72+n20+2JVp6l7u3giMtb7FV5/jQmvTNHwUcYCdGy3jan1h3o
fgg5LBqodoHOQpX5xzlZOwt5T3lT6i7QFrfsk+2N3wWwQrglIxl9tnroiZhJGCTLOy/shFC/VBID
U/OqVd6CnCC+89JzULBISUgJpUQhajlbmAPu/J1az5Nau9YEeMIqH/jZNloBLg+077wfIiVKm+BI
Q5ck+2mZWUnCIlZjurMKoMnR02TmUUEj1fNN7bx7mRiuA2wUFLv9pdXYU0BC8WCPe5AYbOpFbQWj
HXCUNthxPwfx03Nt07iQrdmUtPonef9V8lXNXWbQ39e3zzdHw2emYOl6TSABG7KojyjikM+XA2Hl
v0rBHtHinUSsML1mPm1m5tgFSix35NESDueunHu8SW3bu3o+gcsULWpfDT9eLlcisdrt1tLqQPFY
XulkSMbyYPJgkPs1ODI3hgWLsTRNQRAgtDI16t60jVsV5TRUxlZ9JUWNuJ0xkrAfZODC9wHwmnGn
klHrA9JSgRF3LC9jGSq9brqU18ENsW/9SSA8S3LdyKUKLRqFKcyvrw6nFrOOh/i1vJ+ViyNzvtkL
ZX+bEqMwUQspC/aZGWlfp6/YZt+gCrXQEJIyDzutj15kuw3QqMXlz38M2Ues2u1AJyNOyaRWNssw
C0DBEJAD4ys/k9JkslGDw15OzDZaBCiXMOzy7RteiaDfiu8K7Nv4fAQpu9ut1pwJqxqDcTdN7cgj
YYY7IkmFfOta0eAAJOnTY6JFJ11l1+LK98TMWpr4aoTvZB1ccVax0UOKj+BN96Kaf8USMT+ZmpG6
eUqibKFz5xpVwxdmSfRdFNgCg3iD/Dq3+zrwTJYnJi6fIQgybBSykhh7A3ycKN9ucibGuWNdxFGy
56h7i5WcEcJRs0qE3MXqTC01qr3c7nybNsqlZvV/6yYPqrCkGnAGGEGVmRW4u2GDCyFAfWOOKS2T
Ws80pQTCwMYuUNUT+zQhs8hFhP+/INEblf4+7lXWzswT0SMwkfErpB+nj5WtX1vLIZXHNpiZTHuf
5ayjffBntji+ypIoQ6441xlfsASe7g8FOgbJPlwCOwhkIMsjlJ3FkzRKd3+wqXsxO+hflUFHaQQX
EY/t4g+hPw8vnOnbwi4RfVrhU5z2+IJoJdQ59vQYJbgcKGyfFDaOnJAspaI18emxMMeHr67u2iF5
YPZw1ngcilratciWrN8xW2b9wRsMCHI5amCnajABTXkF2Exl7MntAgUmuM72YFNVr4x5R1MwHvbN
FLN0QLQRz1O02KCYCfAqbUvvgn/rWJfcgmdqHyRUROW0V7oeT/c+JqSt8TYs+FWF39wjoAVsozDl
ItM8jmL30+cb+42/cVyBfiTxQh9Dpa7G16E5im/CwTYLPoPcRvGnuvXj0xlFSspso1V+oE38dDLb
XqSPz77iKiOpJlycG56VeEJmLvvZGdFk2EZ4e/IpxVPZiPvXnUCKUO6ronCIWXCjwnk1Xj61jt4O
g5fwIq4XvQfgwhO6qM0PDjf2auPYV/xcdT65pyNnzugxJIdtAxnrnJAOeOJ7Ko5pf68umBfKpohL
+NQB3ssDZbDHGbRWoWthBXs3Aou4x4hK+ARJcrfoMdt3KD3iTIzvqMd7tgyRXR4w5O1FJ3wKLnln
vTfrL3t82xkHhmpYuMhtIS+6CyUWAB9t3OFPcNLIGC2ieK7IMeQ3x/lFQMczrKayama+zdq7FhJl
mxiSMKgaK1HjcHkwSiORxa2pg17+S/a46WxOmn1DlYrob9jxhNvrifT9Gsw917pt0mmtELZtAP+Q
gtcACwAkxrlIQ4GIZuyYLCYUvNc4cgJU4iAAD2uaQ0QzFeVTWGH8jlN/ypCWxsH5/z+7ht78clf1
i95IGjB2gbSXiNNLGPdDKnzqhRYvbtVCSaW2H4JwINafzt9WiqmpQ88jeEUc6YBRxYnXPvoGXBXp
b3jmZRSfERz+zO6stqcWVg2AfJm6qLCrpd2DNnhF0bP9iAqKAN+mkwLmqIL9lEMXfJvZeeKPtp7S
SS2BHbRvWqMfIxkSJyVPeGPQh4CwlSKxnzJAAs7o2U/1U0lGUZB07jMX2O8HBwCSnk/sfNpCSgsN
uFfE6NKUNhcp+wH3kjMtdhILGWvFNVfb+99mU/mR+iM2EY4+XLdZ05QIZXW8C2VJEfcNZsPdDgsc
nWRkQlbP+XuCKYZzzBrIWCa6hRRC6f34D6lzjWO9QaJl+IPVo5tzkMwWKx/o7BfMWH/fbiDGFCYn
k8WU96HGSZlZp2VL9DqbiT2o/x3qRdnz9CHnOXMdVUPe/QM10oTUhM/+mN0/7biR5XDtKmrJNrDu
XBYHVVEWiGLSLZP/hqi4BLsyvnRO8koHsfyvvJGI/h6magmEc2GdodudMH6T1pXUkPjGbk7zpkwl
ULG9PzamajLbYw70Xg5C446Ol0/x83JuxmoEUfPb9TQL6XtzcocdFindW4WeaRSZiNapwwCZgSbB
tMOc7W/gs4BP51Q+t/M22aGn95gsTNDCnVndy9w0367wowUSoUHdDQyBlR6Cdw0n9XxT3mFu9z9M
phcIkyakRoQasSzGPXTnidD43QqYmYRvTPjdmJrIWgSQjGjn3jcN2OOcNA6Scg+hNLBRobwB10Hj
RZz0Akp5whpub0EfPsYAWbV3Sna6v+LNFLbR+VcvG37daV8Sxf/OSqOAFgbaeaW2pLrygV+mQDNU
zi2cHcFCK8g52xcNb4Nfx3kBIiZZEA6cL/vgO87COHJGJ0LI0oN+OiqyPiBTjvT2AWiMo3f76PrD
GBKDdhFS9CUKXk8ltSAu6T6WPgRperfMWM4+a37PuhgEHvD9wyfgIkWwkRAalAwAhtsmXvnTsceJ
cpd2ORWUzBIL6aYF7CQVT8Alt5jCyPHwe35TyilvSheFTfcEmGPLD2EFGnHiOfKZMs0tpkQXdaqb
ybQp7FCjOLBYGQJOIskdzuzlP85wDvvDVfFHrIwWDQ2nCn0U5PUdXSwEBTSQD5ghMhS8US7+N7T6
cyiKhZdHgu5RBTUBvMcwSPC2SKhyMnQUy9DPso+c8QvOWoyJnQ56OrRTuOl4N3MF3jAHZyEPT6qh
BkncLfnaUs7yqqdsfUiEkl/sjBuxAZdINfzIymGrHSLbf1v47a9nci9AQ0OzYvodhtnOGEKiyKWd
A/RZgrhd8PsctYciM90+yrLDfX5iIuTnQ7699xmHAK2l6jvi5uyyH0V+93xiq53sByxiXeDl47t7
RX9xua/mNHCeD0pkd22kLtzqq4d5GrmOQVO5REMX/WSPg8iQ13VCBnn64ztbZhM1z3FcPJGzOa72
zFl5ofEX96xR8eE1jLvwiq9PHfNUN5mvT5xMdpELwKXnLWsOtabaJ7cZoiELpQx1Tk9vl0dIXFeA
Jq5F+hozC2xnIhaVAkvqI90a5K6lYXbkWK4fF2OYZvqjQa+zDbzd3bKecWdBLNHnauG7UWL6v9FN
32gI4FwwvcTUJ83XBCrHYsY9JIYpDCakeQoBsSCPRDynnDQvhIGUUz5ErFFsVaRHneVe8JqNKqlF
iZo74pEv0L2NMf/U+odjRcqXK34iI3rYLg8LajJysroobqoTZCNgoL05hEW4baYRpGgEwRvgC3+5
W4JZ0Cv/WoDp1rWuoMVDkYfEpmd6Kn2NUXEdVleDb+ItydX77/Hfs5MJUwP8u9qrdLHDr8WCvenC
G0gCCRtmoyGIHWim4w3EteWGAC9nfCW0WGs/czIhqKS49nn4KldNQjpBJmYy6g5O7ZEQgo/OB1tz
oPZXxM89BrR5tRTbJHeOyZLHL41Q3WCo5JEKmfzF2vH7gkNVmpb4D2QZ8Tr2f3SHOAivX9KfgUTd
zcdg+ZMUJABT1gmJ+7AHM8QI0HtRbkLL3yYN9eMy8NPwh0IBVl82S6IzavaMw2FGz0QVuz/TE+hr
B/Ph1g1+rGWokjrL0GSiwiv3fYs9Lrjj6TNJquzHYvKdNePrjbA9UxPe1y6ojCxgtlRgLUYbyF3D
8iUj8aC5NwF6GLtSwDqj2h1oVCda1BrcHx8wo/3R9DpBjtldQy+cW8c4EKT7ctqnei4WzPG19r/a
y/gF04Hovl5kYfWgnvvY6/LKdYnAkFTO5pe3owZD4E8yAxv0+ZJgy/PoWEmmkQRXw9Z1AvdLdYce
iDgICoHSn5DC+MUZrp/qYVtoV9oNgNVR3rq9VIi4mn7rPxbKI55KiXnPpY1WtYSRDi6Yv3lDsJ4r
vPgcSUr/kRg4PfuX+EFh2EQnE8SUov8oJlRGenlHa+HoEwPS7wFChK1SGZ6RCi5IkLC0gcdRrdoj
MgEfdnIYqdsqOFC/O19s8+Hpf7d696BIVABGzj/6SlBnWXg0+DD20XittdpzdF0AD61/rXPrGZTG
Nv+egPpi6PJ7d9EDecCYKQNit0J+uymkzI1D9QfKcoi8J5KqqS2CYnQynCg57RHkDl6zwvaIS0Ik
ru6u7xlnH8BRKozamk6UjUnSsuI/e55b5Q77sSMwzo/mwxnqlL5k7H+tQbyLzbbUardMXrw/a1AM
01ehfqi250TOOGNUBuXuhbciHKBtAmPVzCAwd9/Dpe8epv2uTBClqG3EPEHXX46ZNeY6QXz6Ir7H
tr6iyU/0Sx5dZriof9ui9OiZF4DRMZHxDXsBux8OO4xtipe5GQY+xqsb/ZNG4xFpsUbO9+7xgKjp
3NQz8RhWFWXRjwsJYlCNoJHa9H7nF8aiEsUYVJB00mTcPgYKq9WxSYKZlUYxFcgszzV1ZlLLTnqE
x5VnY66Uckb0E7ldPNEov/WEv1eYWn1FW3fV4T7tFgrWwxCAsKZ6G/g6hgqEXq9DD4dr9PdXS9/q
SuzoeRa/PPijrs06O5uJt+I3NncbW0nf8cEOewYKEyRpdLdcON/scjJ2KaSAhhJ2Tu1J5ozcQ9L5
XiGGEDOgwpl+7tlE0ex/XcsDLhTammc4h7i0OlKJzOkZUbhh6rySjYsDrtW3iKpTpxeH+8pKwQuM
UvYdt/Sgn/DBODYDxLlMQCefU+aZr2msIGIj/vUvIV9yrgGYXrLVishaYNvtDXUegDrUzwJJwQHt
eWUzxpstc2NSrQitnqYzzLqO6KKHjNhLVRmOPC5noPXJe54ulHX6XlYJ3UyFsl1gqlXIS+jDxwwc
g81Rdwh9j17AOPUgXRU1t4Hjv4b380lG6c6TzeTYviAc/+BmY6WN+dkgdEWwqQPV37OEcVFT+8W5
lZkW4hDPcUzQo76ALyJueJKQR4WqlG3tPhKuy8oFazZjGqEgOMZkpJOeScDL8+hyKB4Ke2wlXG69
tE5qVsLj9IG1/DqUEvbRBVi+vOx2VKth5V9i3DV5gOyM3IQsGjB/Ymna7cHNSURvW6Uk/dHyUSIh
a2Cvov9EmVYGEHDkPtz/UamsYietqsp4Xv9i31sZZdyjz7sUIoV+BbxX3vyy5SMMZn44fI0fxNNb
me3cuhfOzdlck3+7KHKxobBjbmJgmpSMnWs9ZlMFtcTMkUZCIiCqmg4yKMRf7lAVDjOPIctR9O7m
RoR0XtCmgzUWTOj3o+8zmgPH6ZAtQiNsA6Lw4sZH/OMfC6UwmMWVAQ4LSo/jX+zkPCwtIGEw/Dkc
RxrKQXjEjtOcYWyHLtVYvCPQ4abFaqAA+/iIScR8U8NTIdeEHjmskoBcfgexYRykDj8viwCxc0qH
Fu0sXXGyW04wzRxTDNV56abOy6cjL0xW1pZqE6BBEg/73mJd+6TZOnrmL9YVeFb3MdT9BQWe+3Jf
WPTKVGGIL6aT2VAc0lJBiappiRV+3NyMw7nCbxlcleepZ+iPBCGZI5k7OgLRMFAFXJUkqHTmUcrc
olEGAzKHAU2Z8Zv3kCqwBx9uObdYfVspyc0WZbtohVG2Buqv8YjbqBrjZIE8MGusQSLqw+a/4262
dZ15fKNHDjdsfWBkQkg8rba6tTv2V+utj0K3msHlhQ+HZZuM3F+1Psqxx2iusn9Vl2cUweiHvrTC
a4aVAevBnhwTEDxW3n2zehW5BLcXK0Ut668mEZ02ABU2A0qYMsNWZjklL9nugs1QIvJwjrJMjT9H
ZI2Aj0JWIopn7SCvr8ZTrOU0LeDDh2ePj4rg7GGxF0RsPIrXoD2gtah/UsFnJNuT9O6A200iMvM3
b6uahOy+L06iNbt8b2cTtFiIcq2U1D8JiZNtTnh4abKvu0azX0VXyVdySorEwHcRGPXgjUfpp3a+
0ax5/MVEb5f5psA+O/n6jG4NnUl9u+ZPGFFdzThnwKQxHnloy3xdJP9SaO2tmVDXnUvKY6870R3q
vcIlpeOPmHSLqUvDERxYaI4aTcCHdk5Y3g2CkzXQH9ACLGyApsy+ReZ072SUI29EjwZuRxXPHke3
+rhVforgW+LXFRQh2P4ou9K7nHGQSv/+hvtAA9gQgR7WhUT9JASmNrAYtVeEn9+YjzYvdQ8AOjdw
LmkzX9R7CCL+C6CPWUFLxBSnBiNGegmcdxIev+hpfKs2agI4EhpjVpgRwry0TL+qcXvpLA5CLrog
qWGHVjMQu1RO4oigannSywk/RqaTUtLCJ5FN4KyngQi+G8NZpxkLuM3cHXzBWk8Z9OpHEgZjCILu
Uy09so1/Q8V2qDJmnriwW3ZioGPiL2xEJF8HaQ6ADSzXdCa1VeSCDkI+uZC6fI9hfILsNtKQlf7r
9AJ9v/gUsnF8mQQFh/lGEkB4ECZ/vgvtALnv1WqovwqAQ08p25WKghFuXtc6KPVbrDvvuuGMUCm/
X3vxPFL09wkb5AzK+/qW7cvZPm+p4al5MASRWAGdNzVpKoMiJTRGjfxuQw7t5rNi6KDLEVh8XkZ1
uw9shajdC4hETEEbVwzbDt9+dDPF1Rj+pDclkA+sAPf6hD+7eNAzJgTu1ufHzCvbYzMLDTad2uDf
OLcQ2BrX/CigUi6Ea9HB9kY2SnNgFmKXwbbNV9EL+iVHuwUY+CxyXhx6eUBxxTH5uD+3Q0ApxRL3
bO+aPI0V9VJLa8fHMDPUZQM5CVCUuroFv1xpeHQHb1074MOIZXQCPFbctF2gZdf2PjnpwBDfGCwT
eV2MHKBlfSWTJBaUAZ6lwoLx4gAOsL6y/xQaGgjbyUUe1CGusSNwqnUVfwxpOjB6wbbJLw5CgJ+W
IqUOZ62GjibKod2ihh/BvKx/J4nnzdIuTbQSOtU6AKuheRLsFEgSBeAGf+eFn58WbAyNmHk36L4U
aiSJk+G7rebZsDywxiToGZZuBT+xYpWhMKAb3niWMhYGKH2MSFJ904sqXuu3O4l+r6dorEzx4+mD
1A5dHPrylHgAHkyWcs6eynyidl040FNLQixcqn7ayP2RbphPgjrZmbrqFVZn1OcwATQn87dxbiDD
xA4UvM4IhNpZFLBCAviBYhL2dZ3NThZEOCF+Kh04mLCkC8gXnAG2zZSQcnIt6khD0kdgIHAqYFTx
Jg9TuAi7UKQLOa5mvvZUBy3Yl2ZxxnFTGLNZw8QiSYH22p77VqcjElHBeqm1FgfVt0GGXZDluyIA
bli8X1oCR3mqoXzzPcp67UpFHiiksy9CBRyn5AQZy7o7OnqJc69AvlDHc5gGcWY6tJiOHtUyd1Hm
/wcYTrD/32x/VQC3kSDiro6pCsn98m3c4jt2Jw8TeLErAcdc/IlBcU83Ta1IqEDXFfXxx2wGVC8o
hbSccCOtSYel+/Cad7TpHmvHDgusmJMf1uikKK05QYKgOZCxAnHu6t0dktAD9U0SIDy1HOj7DoR6
eWdTfEO+MrGbi7Z0fdhlkYiOX83Ck0eDoC3YZstK1N/bm+0iHLpMhxzwya6ufbI7qgVyQDcupxnv
/cwndn799rPh/2ciKm6KA+jVkTFZxBNfBkIijP2Il3QdznIxT7xY+nuY3Jeq6Z37EZCztv3/aOPH
8Z8Ntw+8D/2lj850u4WjTUPxpdHIEUXMoaXSVILgi+J4uxvPAJJQTr43TW0ocZRJhOoVovZMTZiK
PbQh4u7mLKatrViTRqUdiCrga/O2ZiliaUndLTwSjugLMgmSYxVwlahHaonQMLO3Pp9jYNcXK2ub
c2i4H7wwYPk7VZz+jrhIqYMsbKb1lNcqRlc0DRaM2RStOalr02Vfw+RzIgzVOlfMWWEOxIs3b/zv
AHxltU6mIkVmabB/nNbbelIO+7ND4uI4Ya4Cfx7XrwvPxp9sKSouoB/KlqxUjVu3G+phnRusdg9e
yfAWvDwMHo+VrH4iZNZmuM4UA+X+gbr90bMJwbqzICgLKjc+O3ytYw8NUeokYQkhiUdu2U5VFh9I
keVuSwWvlqP/gbPXQJUhLG4tFitYlWL2UKdF77v1zRj6HNVDmYVC9TiThF6B+CfBTytP97PIQD+T
k/az+8DV6DzPmqyLS/+PA38OJW4QYYazrCkasFFfNNvHCNrT76XcM8CKJfvmmS6aownVD98+Fa13
CCsbqr2cQ0hbpQVm2dIba8lt1C9CbgQ27MVug5sughz9EUcN/XCTKbsyAfHgQgFKDXAlVWOcKdDP
06MiRnPHmIX6yC7sR/F3NbOWcqNQ9Y8fTB1WYi/d3U2+nfxzBz1TDo+P6jIVswYU9sJh8W76jNM2
pMfyJkuXClviYfuevOwLwgk5BQZNLcEFKcgbRJGnpQi/8dvr3xd5yDNjzWOlXYGQkICB+YBEVwfh
KIYLwpQcVQuExtrCJQrn0DGps7/N5+I32rE9AE7VBv/6kKKD9TwZ6n+gtiDOIijHlESW42ZXDD5y
cY4FlqtwZGVl47tlhZdkkBtJamwXprgcZAKVE+WcSw9fczhRZMrBqcEZU03Zby0FsYMdFTMZt7+m
6prjAWMeOmpC1hvCwvcIdcRGiOEC9q4GstP1PLQ7y6b3ui/Rgb3amhsqL41fx3tNEoVr2QxlKv+7
2gKZCnfucB8XVwRnN7w2DQ2/NR6qE5uimDNkcIOegzH0RdExpwaXvRblJUp53Vpe0guMzg9gqs0i
Hkc7hn4YT6Wcwotyxk2tITvXnxnbmZQEpSucovPOXS5BQgNuhYd+ou0hE4ajfaqxAGf1zx3467fL
gBD5pzOk6hRbpOQDGBqcAS5pKIlYMsEbeQjtGzKEEnA2N55ZEG/6Vgw0jWYFM4Wy9bcXGteuk3vM
WAMjl0NpyUxsdqsvsWojHBO7702RrI/xKf2Fa2WYL9zhxzdgcyM0xej/TDj1rOS2kEjKaBboT1yZ
f1hEXnn879y9oj+lq41uY8AyIZgs6rlvB9hXDSZ0AeZVsA3HpBCysv1iWBm/S4m+uV0hooW4caqM
TUDjD9vnrC66T5zJvYk/3i0cII6EOn4vvsFlggrNLyAhDAopJIXEuzV/KHAhB/OGUP55fbsLKrRb
HoVZcxo5aWB4oHXKkqzmtWLRjOIctMgG6GY7cZM9TRR0yOAOl2JoqWMJqqkv+Xx6KljBMt8AF7TD
AiKHFnV3hjex9crFPuh9YVLT76sCJxcusqbk0t+bF7J8QV6oBp6PwUxxMOfAbDITHOC7jlr8aPzo
o9Zn/A1qHG3mJW8QyTK6Ogqf7QjmSyI2ihLrCiYaq4NWYkJE3CxuKkD6OqmA1YLFJpOMO84NbmyJ
R65YNQe2FEz2uTe1sSzPWDC6p2aW3iB5hPSxlzibVfWdcYl1qw5SK82idLXoGV3I2uPxViBXbCzV
gUPWgbp8fBQYVOPd7pbAPKWfhbGUJfsgE2Tc8LRllr9TYrdGnrgH3LRI7nCMrtS+ewE8tzdDj5Hx
dZqgbxPx1+1eTHVhxTO1TOk+GZnL+WWi5URPWV8UVZKT6a3OUbhwvkUaHyanYXOR+pHOPfqOnuv3
R2RiKWG+Mfotrm8DPSewk9n3IW8m5KEL7MtH+L4d/CrfgU8iCO7Y3vJjJCI21itvkEq5E/KkXY7O
O4dc+GlwvAydi3541zpvlkiTaQwBBHlIs21ZAs4NsxPQtD62xHQqQK+8o4ttev+eXApl1tG5oMnn
yvvde8NlRaPJBMl9wisjHv161oHlVed0904wKG7+d3P1iYcYWeRmf2BVBM1qDNI7mM8uP3JnM1T5
d2qlo8AyS/k4T1pistrBSBN5CEAZDVPz7B79JvnXPFPcZ4G+CqhguQxKvGw3NLzWOivqpI1jvLnk
nLVPXha8+ngT+qlHJa+JBLLyNeeovjsypZwo1B539hhogRlYVSh+kfg/EPWcOALNStN7ZqlnoB1v
q25acWI/LCoWzuH9UlJxucMZN7ffckjZBU/NVC3r24xG2pxolO3QNST+kQLYNFqijLQRks/DYMAw
QwNNeRAKkAsIEGfTpMaB35ix01ahng6ziyEsPOmgVwqIBsYuEzkDBUggmXM1raynEF2BoJWC/JYh
BDwx+GBYZpxF83b1gXqbGbMQcQVRG8IajpKoTFLEuEpvnEFjzGE34mJpgI+dzYIIaPFmCfwnSIFV
M2StfM3ajsG+lsjEEA4ssW2dsrre3YWrbJ/AvTc7TMqXEKQFxsXHKO0KPMP5b0KYZuAcakpce8Xa
3fT4SIlyF6o31d/XjF3Od6sIsdD8e/Jmx7YrGVja+DJI/k0cRfN9/wMlPKQOipwrxx58MkIdk5U5
1PJaOfL/RXmeOtYKMl/a/2rccf9Tdj2haC/nrATP5btiwG9fii5VuBU7AMgsXZCP3IIW4UvkURuv
q1UBRZHdk5pAmTInXAetVkK5TmfZC6LoSZWguW3UC5padHr5AJ8H6gHRrsbH4NruG/+tgzdU9Vb4
38WI8noTUUo9FIabo1MG13ilm94SFfnGrvc88ASDIaU6ME8Fcnx3p5JBR5fo0K0Hq6Bq7EzL7hgc
IIPHOmR8YvUE5+1TfjAiLCTygCWn/nrQKbxOhmkQccTMsYOSe3VtpAspDVyfq2ixhAEU4mZR9FKT
VXmSHB5O5wr82jUw/fQxONsyM6esF57E1rDZ4yvvb3WhqEdjKlN7qjmYU5tcHoxaj8pQr3r7vvBz
9IIrK/Q+pjuZIJSgHh5nDSZDRmxjkIfLLPo281SybzRRWXBahC7OBaS1R2XwPYDYfDjV87cPAXTd
RLdKCO8u1YwMAKKzQfj9dMFQQBymlkpIQ0kDogAGWoLBhF7hOalPla7TsORGqKRI3C/IF4g6Ai40
qb+rxrX+Nnks2RE9lj1l/tMNSBMyxpx+If4vWrrR3v/MWWBeGr9+HO/vYJoKnsKanS+cbKEhcnF1
4aqMT4zW/h69FvgNWZqwEWm8hF+cZzodrCNlgBBv3nzbzkK05rtrOfSL9jWgeGUhgC2Tw4oOCVDI
q1poaOPJTYKBBMC5DQg01hLHuUWwRLZqXWD/zuKvMX1ILzjUBiWVCcp7ImsEUcwXsSwlrRJqBW80
nfVQSycC98J4c+qLCkFzB+ScBpK4jl1/0lahX0h2PzqZFwuaSmE69K4AHElDAZzldln8h14SruGu
KB/RFacvHYWs0IRcB7xS4IpfKqxX78h53Ym9j9cUXXHxFrusj8m3BU8HWevCit1AFYz2dboRE+HG
iOqAkCeO6j3OlwfMXGgDMNSCVfiCHXgTrsj6iGNVWO8cVhMMOnScTT7krihsKJ/HTPK8NWuuOExb
lSyLnBGD3VxdR615qgnQBOg55XF7jmnaBEC3WCr9nH23jlPQwzbAIRBEwsOZWWux9nVcRMngRRG/
R0VLAfZ0pE34+QKWiflnmsZauThHkOLnY+U1CJkq8v8B69uDYN2TCPrIhrB5HeUVR0MxmWmfpQZk
PUakYwwS9IC5J9FdwRBUVH4xL/ymImchbf/BppaSuWJkop+P/oxNIQaeOc8Uk/J2IpAdUc6cKBkr
1BlURHFG7EMxt8YfNlZ+KKN847wvLw7dcoR2nWqDKHv+JGEe2CYVaDkzF5NW7U2VJoIqfzFd9mWY
cRDH9zJ5Ezmd9Mo7JxosU99VOwrWcnd0NKSzyZuAMreP2Eu/vKNk+SYCTn39grK5Zw5uMlcy+Od8
NT8kC0h4Rnm/UU1Hut2Ag60ldk9kK9ULxhD176UchYEjbdvRsjKSQJdOfOuzUu3pcJjFwEmDEpVH
PZQofnSEZeptEx/mq8wE1WOWqM6GiIUHBQ3f4shjDFkv0pj0q5LvYIydPRMo0lY5xf/oxzDHg6fk
+OVfbX7nn6SsDnVFLEO/YMkZkFFwxhdIUs+v1EhqWFghLZQZsTGLyWFdlQzSp/Q1S9+JqdOeqCp8
BVIjFf/SRpYMzT+0P3bAszZ5P9MAvz/xg5jG+hcWofFZTqYhjfbSjnhuKbUoD2/q6DMupDKeT8Ur
+5O3QPeRh+KPJ1ehLayKP+LwX1r+4kFvhbkvVGhK+8drkkza5aVV2uSAQu8sOafCehG1igmWN4QX
caqmEJYwSOKI2RluRWyIiNCUuTh9ji1qjhcIXYz5iUyVUqytwruWtfYzxAFtjSkXUOASNBlSQvZC
hccLf+XLbYCl9cfMLwTbGx6hYiU97wO4JZa6WyyRoex60P2ehwhC3JBniAzss98XazB8DB1z2W81
CKVZnZ2/QsjkfZN/zsco6OhptgC1rcJM98X/gIP/QgZjKXQYJ1d7PbmLxyR+8LWH8yo42v9so65Q
IBD+Qnv7QS/FG3rqcT9mPf5yEiSHHKmxoHOl4ihGVm0S7zrjr/hpOfWAaOiMAITCsHlOePgULFfc
P1hHvoVgoeoSEnNz/FIkiOKKqqX0MVGsCTy5T43kj0CoVL0KrzG2qWOQUE+5YWWmD6ztNGUekqbt
WNaJX/n94J8XOQQs/Gr+sy9zyCBFRM8w4KzQD1TL6w7gNe/yAfEHAwN6Ae81u/KfwglSvKCkaoNt
N7op3hzYO05cyrjipJv8WqQZuDc4Y2uIdbAzQLdkCxiliZnv09ONzUIXpQ8J++Bp4uZJ6Gr1XtPN
k+FO8Jb0hfCJ8pgVtAilxgt4yBi3GoI2Jt8/vamhTfdxMDXLp4NoL/12njUMrSH1yPAAeqb8u0cc
N1tzofihMBdW41zCTxcE/TV5wd1akwVcY0VhXNl/zI6uZ7EPABJ/MSh8L/P6wZEPp6cBy+X7jdzU
UQSPtPfssqhD2D/+GhrTFJmOZ2fZq2tNshk+a6LB4H3kI2dI7BplEm/twn5o9dnTAmxTmJzpNLz1
V0WdNmLcC9nOHvd0kpoMYT5ObY3mhArgL2a6nEbpXTUFYpF/bB3CIzMigLxxozB8rnwySh/+tO+z
cj8THy4+EMvDPQR4whsm/7X5sQh6QVYD0XXT+YF1PwSQmWvv+t0FwH+79VIWkwSLVLYTuzC3FbHX
1vIeLc3/uQxKvtbP8d84wnyP6Lu3cyT2S7u4v2s6nV0gQPaUA4SNP/3wrI4NyaKQRhxOZI/Iz4IX
JEo4QJ0gGgkj43/ACX6uR/+QWH+1i51BboULgwj6vJ+gal2SC8jP63+hQ1cjD7UeqcKOkPsrMiqd
lwSkdQdCqgBa3YxA3TQ61aZ5XqV5GY4WOs6m8qUrFySlvUw/VTu75qJO6bK18g+QlmgznOo3cEg4
6oWwFMo6w7puZ5ZxSHaQyURFj2m3JopcWn5F2IkzG2Uh9rN3WmaREGhJPQKYX/DJjuYUOJ3pr2fe
Uf4DXu+kYzOwbgMqilEM2fQyTZsvDVlOYwu7pByAbagnu6QJPKm6MXC35TeUO/CZizZSZbrANiKo
lyOAnt10dUIbXu5uFTw4Bk1evQNS+2CYhHidFnp6jpUDJuv5b3jeeu8GONxNqW6zqYuFQDwsBJYs
hsJuE4ytz5lg1ALQTNOWSQPHbWRZTM/gDpasX11a1EQpzJJYj7/FqaR8xNtbtIPZmLaddZOkJN2c
w/z2km6rVbKjHWo52Ht8yDeX6EuI74dP4TSqTn81m/MoxO6EOwGD3m/D6swD9MqeF7oell/I7iY/
pR8stPjf1kMrEUw8ibU5pt8zTjyQ+Wr5o5/N1sAhNvwUsUkZwASXLFPRKNCwlHhDP9nPnxeRecgW
+r7E3oE8X9KVDlnQlqIeugI5gAx4hUtD0+NCkEvfXFXY203DNWVkL606xYk7QgALzdUD/zDwYl5R
nWCKqaNIx1ZjpLgMp3UX2i8RkefbHFGViTZ6jaMZKxL0JpK/Tu93Imp1af6dTZlIeGF1mLUEytpX
0DM1rkKyZztU2auaGzxX6VA4yX8YdQjmMh9YcYSLDY9Xm6zVJdTBJhWtv1gYMAcYp2aX/09HkU69
3SNSHXyDkDrCwOB1dXKo8tFazUGMXil8ymeZwxLpUAkGlBnWljwpdxiBimmQwIa/yPgh1cfi3YcT
Bmz2PPrpgTT16qnvFH6qn0vtTRvgu1HW8PEhoFHSt3sd1CzGxT+AK4yvig0uH2hkBMBojT6Nqnvp
XS7IP1GqkQ9MWGWqzcABtJD9KVB1Ea2eXg0vjr5tYPXuU2FxJAGaufDQjQJR2vs7xb0LoqNbFGmK
5QnnDG7OTkMBA4tPfhNTN1LSSNnixB20njGjpGEqC6QGwGOGk5QiJUPYkmzxUc8RxX7XqemcovVs
DfJeg8OA8J6F8v2K/dQqD4GYiTBNwl+d7s0zr+N3H7bPcJYb5XCGq3OO4r5Ke/UGRoevdbvlc7BW
B/ZP3PR568y6CFzAFO0vRWAKbP3sK8CXnHMSg8EeNiJ5v+UUfinRauZWmQr4qOwHLbh5XhVxVjIE
szNiZ73skBk+k8yx3iv150jCPG6uZ9l088DLgjp6Xx5NHrGIR3DvP5XZgdThgFUp5qVs9vAtsyHr
lL3efnlPEAgwNSe3XSomvB1GQqjMuiDmmXdp2nLFarx2r1PU3Z7QebtzRxepqz+kEHlljtc+dlB4
A2i+rXKu4Xg85LRcaolp0Bg0QgAYDXZRj4ZoP8n6/CdjEtG6DCAHJrNG1xywfZci631epNe/XsGS
ezKGovnwIhj5jbmtgIPnfXNOVFNvaKZYK8wMM6U7RVYN98Cn5NTX65yJOSo4FWaxVhwLr7/RABg9
eKRDLJRgwgrEWy67HyvK362ERcsZoSUQTO3fl/COumj1tFI92gRRryA1vysFwFBqVegXpR1cVADf
Kor6cOnR0vmmLkbwN1KrWqwWEUqJHTic53/k6P9OczlDn0741jPUHSymKBXS7n5J4OCwk/62amXh
VTQxreLhHs2k+db3xaULKQ4aIogC4gwdTFbYwhNRfgHCGMQbJ+8/HTugzhy2XqTSrHq93X2F+wdW
wxJzMPlfvi1nvGUybrEdi3/y39ildih7saP/epKOAvjuvIfa/m6EgfXQo23DOmxUM+8ZhchgS6NM
xOe8tPA7gH6RaO1jMndt+4a0WnZyZSBNVmQppR9VRSPQQcnzF/04XCB8MDOMHKBvXf0bRIOuDO3J
0zr/cU2WTIG9g6SEHxaOBGOtvHY4j5c1Dwq3SG5kVMop4jBrvvoDM+bG2MJpXINwb/tOI9hL3KcY
GjrqCHXDz8T6EUyrxUZ9klMc6HL4tEoCB0fOLy095jq6fEVrdVAOmM9Dvl6BhL63wPts3RGi2nbi
fsEoaJIxDbdx+ufJwc9ONkGNKtLpRMqxvD/+SxeGCsCYwyROSBdT1fkym/yldQuhLbOuJfltJ2nN
xfjqrFjmSV4kcx2KMl3q+rf5aRcTLmm19Lg+ufLTj2I7y1VL3HnSTWrYNCpvts9rzKnWT9/0ZvvG
KC7XvanDnKW/N3yUrYtk/Fz0wWQle3s2zK/Meaim0xLbK8lTz83Mw+lplVYr2Gmo/BFPCQTSK/au
J9FCdT+UtvixX7PdQMj4bwRQZyfqX7P6Mpp5GOa4g/4HiEyRKoZiihc9FgQkeV4jNFU2oNT1IQVo
rcgxgGB1jPDXX20M79xj7kZm5RPOzWZUEkQByr/WkIZyuIfHEbN9eNXvIsCMn8WeM2FSgn9pbmno
Lg2T/j12X00eCMA04+2ehj05cySy+ZC0j4IiAE0EChr5nTHpQzT7HHv4D/kmu0x55nGITu8UX/Ox
eQz+9ffHUaYBZsQRrMC50PX9LhnN59FVJOwpdg93Yso8xDT5svCcVCSW27S6XSR544saDu20gmcF
SnUBhCJ5K2L8u6vfI6KxP+9CjeUogsSZVBwNoYNErsStkA4RCwiQ0MYGAA54/xxTReRZfxC+LDEN
yWPLdhA8AOL16gkDq9w6tfXV3pPSsJ2u1KOmwTadSz+dnmh1y618LlXWjG4efcjU7vVWda5hisI1
ci5/7ljqLF5C8TlWizdLS44SizoF4ylYv7MaV3ZacLN6SHW1rb6AyNK0XNncLEvj3XfTwJpZy+bK
sBLqysZTNX/VTID9JJ3QWv4zpuzaIdzdtc21ySrLKW/cPHLRSMrN2ep5wB8Vk13q8y7vJ/hPUhTC
CScAwEjRF0rXO8lgTp+zUWZYCJgLCdGq0qip948/HfSdFzfKd8cAYBgtt98NBNDkMx0pSByEIOFE
dJtsE4CjZ+VdNb87EeNrTmMf6TioPLdcErWScxTA/tAKKylMvqNfOeZ9zYejs56ETaPznin9PtwG
bcZNtHkO6CbJzbQrE+0Ra0irBcnIRob9jF9fjIw4bBhNlRYuuiX6D/NcZsuaCbqPRLCZW8r9/QeV
TqV8AyUd/N9oVaY2NTMDsbICEWksvf/hHrGkDL3Qre75mMHCwws+HOzdma6RY8GutyY3+i82e+Xf
h2zixQF81P1zbTK/+NNKuey9gHrP6o1zafII/Dtrlam4ECP3764LavCA6PyhKiCE+YoFp/MkvaPN
JK3TJmyipkVYpJpIzTzGxXsEA89IhUktnTxf4aj9PHAgKcJa3C9BxkKkt77oD5IhC/7Z5AOLZefA
+z5BigcRSxka+4CnwtEDm7wbPR/Wz9BGZaglV7sHy7IzBvYNRcw9mfYwLCePABSqUOyCXt6V5hDl
M81MvnW91ObBI45X+LO3wdKh+Aw8QOy03ZXmjoSBB52PcsMToFfH5om1LYJxBbuGKeXJRDjqFsiF
yRc/BkQ16YM5v5+0+sSAbkt9fBpYZSUsrrBAbd+Qk2jbnCx+sqhZc2BOp2CPg02zlzOjwLNlJP18
OwLExAFEyq8N4FLDdJ6aDAtMB+hiWgigBLez4aSGewPrgZDNC3ND7CSF60hCpzQnbjm5rsGk/Hrx
XNf65wqTkN64FVMLkObUBzKaoijayv1VfVcD6kDV1724EjbAM2B9G6TkQHcBakQaYx+E0Dltc/Ys
kUc8A2Evu2ejBk8DVQ/ngLc8SC9R+oFMf5rF+I04POehlEey09Jf41igYKPVhU0JPas13XHTfcik
bwR3H0TqUGU6t2KvTnJtKZRDr4uEJDrf5ET77Ej3/FiHRYHbfZ0T/09zYiQs/bsxTmzuR9PjFjni
6gI19Fg3DYai/SjBUMoAWvOd8Ykw91ML1ScVEZlLU+4wPPJWkTZWFZNeVPkbPEYb72Qjyh5dz8sM
8h+sZ6bfQjX1YYG6qcL3Gqr6ULAGFhYlv4r7iAybs7QfXUVQLZC5V8BSEuIM3pKtRJbP9zXJ5smK
RGLOow5VxaupJnNRSYZHhnPzTzN+ZhVBWHw7SHivIyQgbXQX+DgrAd+X02rSpJj5Vi1Vb+t3vOUK
W6qZAYECcoxNOaXBB0bYEUdBv7F8mJL0Hr9WTjpZYO+KU9hnIfcH/Svzre7v3b0opLzaToyGwmqx
2e8OQkrckMrvhfmXJNRZoJwqAwpQt+PW1PvEJnkMwgZ36uLHSjZL2AvlANoO9nruThYQcIQkzcGM
rWrrR2w5/Q5d0WeTZEjbGpjJkHrkg7kOMKc7Cd5TWk26+yBm4vMdQ16Yno0h9jC2VtXUal68ZOqc
Qk69pMedEoMzr+arC1wOUXo0yYhAdgCMZutmfqBVpnaBu2qy/wILSyBW7qKXDF6AhJPJzCID+A4h
Kx2b/FO+AIAgSFRAfGPAIZCkrgT/orkPqP9+BXRNQrCDcGyjnMjuAZa98i74o/wFKuVBuq+8uw0X
uWyQ0LcJX0uZNOdZdLzC4p0Jddvz3GX1qaWczIuOLdplZpyO9UTiFMpQ4hdmsZnTO3SQefzmI1dP
H9XdbMtbEdnyMlkRKDMty7AwEmlRM2/KeubVAbdLGljoE5uidShpeppAtsUXTthxv+SP/gc0tkxZ
OFe8cbfzmLOyRKhGXJOAHiWtGJblDtPIoiWrC62xc2p8C8e8EqjG+6W/n8Tli3Sh21T6byJS09il
cpB0HJuD1QjQSqvMzgxgQX87PAxwpxzZG7yAh87nOh5gDNY8r7Zvdrzvc8Pnlp9BN2kQpAvPOPKG
x3XRZztAKpGsFhYECK0GjAeyIEmJc8V56HQ5aedxtq6VCxC7F+SPdfA4o/Rn9bEtmZq0swiEOtTd
hxpZ8exepH8X6Wu+z8JIqk2P/J6gki9qv0E+oDqrc2HWwaiMSUltEPkFO0IN5vgEM+8s9bb9NCpj
Vj5s9A9kTZ9H+tm8wpni/d0Pj5WGBzxAMveAwb9LKxGdLGASAMbdeQ+wtDUv5JfPYlBeDmbxmhSI
e+zH1zasvcAQYKV2izvOKxLrlP/80e7T83kq2yxlLMehC4mUdgpPj4JOJNbIPjrNXnZNk/oqi4+k
XYkFB06CwYScJoZa6EfGqm6v7VAO4evd1sxw0/nfUP2DMziIhr+UkjpvP6Z+wVce5Cvv/Ad+/AEF
VVY66knvWN+bZ+qG2+NSmTGFtWHiYQaijONprcmA76oDgd2+e1uFrJbBah9Il0XV+pcJTq4vV2Z9
TCb4XmChR2rwR2MNr+g+mhe6nK7RRZcuTfaXqODTV2Ii6uTpZHK0XHR1yd1ZrOC+UAc8SWW9X/G9
0hMfwHY5xj1U5MKdCpi0xK4JQT1cBwBCL1GWnxoZhbqW4tDUcfUj5z1AO4FwXcHwRqdXcsKMEVVI
dzKOnb2JblPfrcPLWfnur05MjkpIt2k6c9dXwio1iG1fJG6O1jcpck+Hm+eo4T3AcO7db4EAkArS
pNkP7F85sK4ESm3vw/ybRaiPrZZD9MtjKCk4GnhcMckGnWQz46JJEQvsoxYRqwp/kbo6mcthO+JP
jVwqAaMGkBcgNGoN+5TMyZ2Mc4g+BFX0vo2OBGpM1pgJvbskO4EkZhMUXstCqhoTKejsnrAlw4RM
QPAK9KfmEXO407cv6xma6y99JG8Xs2XRwzVIQ1p7pG2vD9nhj5TElbyZ8dXa0PYh7C/k1w8/u35g
UBtaUOtZNk4yjUzbhSiNpAmIW/FYxMzpp3vf/QJQNgtQfLT08y2WerJYCePBBw4xPqS6WHrh8WFi
FmRl0FofW/1WnaMTpz6IChoruCDZ4v/rulqt46fKs6HcTwCJMYeCro3yEviV5r3iJ57Td0nsDuhg
hdodwkLI9xIKNpyVhImByrMTsmdjY8DLB0pnaXpn4ZJvVuq82+BxD3Z4u+TKj8BB1pQkBAjlYZhX
hrehWEcqC74kvB1y22uPjiLitqB1lR1FZot1tWEoj/+cUZRSherGR1YUu7nrrnfzg/y8ovzyA5Ke
oSu6OEWWUKSU690HSCix3T6dWOLOPZOFeiKD8xyBPy72FwIYG3rKsPRx8bZADGZPSiP6oZvd9IAf
MsxPvGX1KFjyJHqnmG/YZJvs5Gw6fZDZrmXE84cCkOt00YB/KKS/ckN51OLb4pIIq6p4KUaTQb4Y
DVt6FYw6QtBTWHuJFMcz7qhiyahqVftEQnCxAb8rudEsPlxDQQ4N1XCbntWmVxPCz/EByB1ulCy3
vw5akrOMDSfMHOI3ckzADBc7zs+Rq44OHN1cr36NwOqwQXXBC+NHBLRT5tqC5aNwJG5nZAzD/g9f
zuJLttLz4voeXaKi2xsUNLpCwEEf+sub/1eLFTiVMXgsaR4dc6dCNYs/mL1yZGcKe2PH21MQwNOm
uOo9IQeQACdKe8tiwzmjD9zigK/6hBuBECSnfNAMqIrp9W5zupczuKdLMHYtpaZVcrVmmMGiAWRm
3dNW/XAa28RhRgQt7PMmZ41q8ylknrAL7lbL8+KfWGMSpNWgUESQ44XPKqpsLJh3IPq47TDiRF66
KcXLSeyhhLpj3ejfBD8j7dJOiK4o89OYm6P742N+NSUD6Ae42N3d9NTIdYC1FxRXB9pa0XND9pF0
IT/CTrse06WXtI9hnU3MW6SG5xElXhnVBhU/ybC+2RMKe9wx7+gAwio15sRHkOErFRLRQ8U/alUm
ePZejM84etWSPWq35rzAxtCauUvnYmlwZcDJ0FsuyaisNzygBn7cutzfqDhdwdWCnJb+b/imkE1Z
FB0j9uALy/LFYuxlStU15171v5oGM7psgu7QZvDBymraUTKYTT4laQgRfUCWcYiywqizjbWK5gmZ
a+ffg7ZH/BNY6leoSudjCKligqIzVyhasQG4R9Gp0Q6DKrJRn8ikN2C0lO7Ua7N9L/HbHw/3L8aa
BgH3pE6i8ZdM0QawE66wxukH25PohctQNuCY4oDSLx8TtWyBgCqPHeV5B0AW9zLOykzGjqwjz5f4
G38ey8Trhv4HGifqDGmQ+sm91AWPlByJT2gDgUwJ77Uk+/Lr8hC/JGVfDwLmRkSuuJy2b0+rekH6
z0Cvn4yJBq3U80QT1JNcFY98SXOoisYtVU4GUiyOvQ2wq1ssWrethJicj5mOC48hHWlYtz+FJxk0
WH6SJVhDtDGIc5qVjQ3ROZ8BmzjTg/uaiUL4boORwum8xmf3x6UYYb8fFWuyHRpAOkS14Y6r6Q9E
KJnJ+sBfq28F+GwpFJ8UHQhEU6HiqHuPPIZoBgnVnfM0R3mX8ehCRQVHuNgPnyOzck/OKq47iBe5
Pgx1lVWLT4tokhp92oKELr1WvbtV0C5W+LqXMGctEd5NBQt0finVQc76v95dzuYuIm28LYDLh1th
3G/laBZZw7IrclfpaSyzVzky7fjeQdli2BxoVcJndf/cfPm84uyHmBzWNLGMqUDL+10mvSTf2b3j
jvKh+6KM4xPtOObUc3RyqRp9+5rWCkDFFDZxLUy3zgDiGHiudkfL80kaNXaAydZEr3/aLgc/HVTl
rSGVX29yIT30qkUGIA7ytj6GEHHGAVkGfJ574c5ogArJUyh5bW4BPilHzjrpK9gUfWaC+AJYqMO/
e7rHmWwz+eS6dx74JrzpeFzs+ryAoAofr/jhECUeKgzjXUC1iDIRvw/lCz7zXMPhSKriPFmPBxTP
jhteE0DVJiRa/d56h2QGIY/mTw/V4SByMGIjZ6FjsNrvyglhStVkXso684uswyZLGSgh8oSTXubb
/bayd7agkdFo8HBDzQOtesufbdVjcSufn9keEn52vv9uDWrs1betaP9P/WIc4HkEZmdUmqi/IPn4
dhlbMXw8dr3ofxjhYSrXHY28tXAwRI3W5zWBzof1wEfaL4C22YZUNsZMP/Q1LEw24kfePBPcPpeH
Xc0uv3cPxWmU09hEcjtMnRn1GKmvuM5d8M05zHsePbEUTeEmFlZDDWmZjRAWY2HOs3VW9rWGcWw4
PwO7pDZfKDIYOBqo3pw/LDEKB8Xvj1ckOENClKBP8Z2tRw8+yfMR0aASZYyFMXwPJ4qfG4xbVsIE
2FZWb45jz2faLd/UAIZ2PQuR7kUqw0RSibb/1hKAw5TSJ4zN0ZOB+4xumQs/KSNDJsfZYXmEST1A
iBnaNz1+pfheT0ef4xJyU1MUw1D7SZqwEPu7bpDgpuSJGt/MMPYbCJDhzuv/GqiOT8699O58KQlx
EZxWzWURqDE26QZc/F4NdX0Yj3TgPHvG318Y91LySbduIKYRxlIXBWJCCauJ4stpsPbTTvsOepwl
RZISPrMTYb/okJ06ZTDKzI9+7DCq0K9xoyZJom8gN3fpA6YcSjukHoJM343FAb8Qjq3yYNWnaVx/
yHSzSplHj88Udv1TN7Xi2PYotMkK2WORTeg/Ic6+LtTmLRIdpxMPJL5YgzHv7pCYr+4ItNuutd0z
117c/7aGxcZHcDoxRW2l2o5C1Uat6jJr85AoC6xQgZbRazy7Td5NqZxylaE301Pok3E8KF8pzXp/
Tb6ZAg+woPOVg1R5/sMlY2/TU00TY3ngY8GFPmcc+b45833RQF/+DiE3phNMi0uP92lp80OWenJF
g/cVZe9bofZTgCuoy2ALAqFi/tP6EFO+LMB+jZRRJ+zroJSUZeGcIzO4UuPhgahZIhMQ59pBREDH
YzC96QFcz63x4AkBYF/neEyfDwuN3S3yRMDbcqyR+5489psx3jfurCjeuIdforON5exjGnlV2272
ntU1/F11PB+TtLj3RhRWtkbbvNH5/kbDx8T/1gxF3gLimAAybiiAXZpNn7ijpt8zqNdKFn8RXPIb
rRuRPYVhn6E99jYEFOeMdWFQmRiFKpa7rsZ1F/8ZramOw70HOJb7cIQC3BjNa/MTaNXkdNQp51qo
csOBG096yv7s5gT+NlA+9TeS8eDzVfP1Qj8C5gmd8NKt6rjZbfYXnLUrq3T02OgZycSkISO6OBIc
vnKfgj6/rhj0zc5ns7PCvYMZa/mBkzhiKWi0uLj5Dr/Fd0evrZZydhVBzUIXInHkqI7HqVQ+LqOm
dcXFpb3ETtDH3y3c9DLGB2acFtFa43diHNzC+JnlXVEiUE6kxMgm8wWOZ4BmdPzdRvzaGU3jA/sc
0ROYcPN7+S6bzK8lN/UYpXzIs6+LYJWYWohi/wFXvvbPXFJZqn4OCj0VrYulaXGSXotqHMHWnHY7
RFGHnyBHd8BITPxfuTDmtnydS3DwFCftLl8MKVmFFCHv4PkOkgPFlN9b/YnNyrmIpnoQzjSNfatv
rydHF8lUhWW04mFJP0tmzPXKdks45KeQ8SCuyGbtavr1GGq1sYEmZviTMwsLNIbGrHDuKdBRj3IK
lRrDlS1wW+5GbAUYbdnknESIvDqUwW16zcSgQyVpvX2F9YH42tNcx6XRlb6ceW4Fkhn9kF9zkyId
57jamoy0gETokbhm//XFKkjrk24U+OGsWoJriy34mQgRFm8mKb3uiu2KhnSak69XgwryL4TJh7WZ
E/Qx5entPf4DI+jqquABNDTswK9Pcuihwp2fhYY/SCZykgIhK+fRLW3TxdZirWVvUyZSiZM7dLcp
RcFsl/+yfl+QNXfHnSNY1xXGfUECYV7SW6TrMxvmD8GT8DELNvH9axIsG27eKXoeQqmqu/XF4q77
F3SVRB7A82WV2oF8n7jiX+Td+ungA1N3XR7fpXU78CpNS31UG/DvrchZAJ06ye8uCNLZU74H1NpL
t2XSMIUQ9ucV4TN6J9FpE9thHtqghc5Mxdm3WJQeDq4WsX8d4c+qPjAro5FO12uxVv3LmJ1Zljpp
vQ6I115+a5kPc9cCiEs9ye7HdyQsqN4e84S3ZMuvEYmQZ6BMDM9ZQySx2rsAQoVVXsu2/4p8b6u3
eDDC+6icmc7C+afXHWE755Vdk3NWLu0zXlHzKoS33PbaZE4QrRZ7YrmpqzO+7aBPz0Cvi6AYPuoh
322t5qlCujQZRi0phHNkCgtdqVwUyrEpQsBpYEV+kQfKt4LZWIECUHTT4enUrGJ0kPmIr8zal8CR
EyvPHWohl494I+D2cgMzN+kCnMxB3Su2r939rfpwA4Bsg+9eboU7Xc/eGd5pVqgsZe3NMfXrU3Q1
jKjvi6xgP7XjdHdYFWXdFeExK11xCgYXFJDjQjkLwBTT5KkiQnllb8npxIZoglG4lZa19zgfEYc3
G1Qh+l+YoPX0CJoHV5eb22sGWUZmX+FHRQ6J9CagP9uzfDd0iP8/w4zKIxM6beTcHjy22acByUX4
06Fz4N9/RAJ9VHLUhoHSUotNmMfpfga65IAC9974Li0+vhNBo0lAPG7rhoRqUeViQfK7P27MFs8o
XyNoeEMp1v174Ftr46AGtzo307SUaqEW9XHiYkjMLUUxuPhOZ2nj3WoyEoohAJ/Gp7qIsHLl9tfS
sZh+mabmnbt1y3B6B529i45iC3/tZqFFvSzOzlzOu2CnPLFgNECOHFb6rFZXd9yg6nSVIKDb4l0S
ceKITW/R2A5UmxYHO9LUh7S7ZjgyoIUfU6oPP6mzcan+zj7e+WKQM11BX8/YsrnA74Bp8Boe8lwg
FudZ4tsIbll4qGPlY8PdEuakbi4qOPEogC/8WtnBFlXvMrZYKqZAWkPtvjiG38t8qJSZMFR+U8hi
6OcQvOwhpyX32ywkt6lLBKOwldX9TOMv197it+3O5Rap3cR4Zp3FYiKLou23rQA5rt8vF1tA5Scr
gl5DDIyAaxMvybBRpb0+NSVhKk1Mlf1oYAQJH9beR/diZH6rRPsyDV+XwlE/KTSs/uiNMTnOyfKm
wNWtWJ59Aye5n9z1o5OkJHVJg38PHIBtNvb5g4FdqIO75+kd79a7x9GUICDTthQ07iiyoqt/+Sbq
jhtGUG4CKuAETZ+cfyFJcAkGSo0M8sKBvCHGXd6XjNfCc0DzOt/8/tTM3q0f6JT3VLdTRa2R8nLS
vp2yzAyLImJhLQD1BFG8kej1efz1N8b1YUrphXNZSOHpCktzuezoOP33RA3Yj2AT5GmXi0Pne8GC
P/71c57zYOHFDmR4auqr1PrAm9yq8GNovi9szVKK7eInwhtVAVegv5NURYbL8drwjHfJf6Yuzy7o
NWqYjzDQ8BkqbcJEoM107DISHAp8uvIsGGqiEdWi7P53d6Ofs+hv7J/bVJbjfpgX8V8cURjPJ7P/
J4HVbkQPbp2mA4pQCEAIiE2VPtarZJuaThMgn+EjelhKJN1MpzJHfEaYOErNJrLcMHxnqo1WmF2V
eWJu+R6nNdEHAjt1Fg3zvD2+yyv29fHebvcpuHEe3FutR31sBzSMZqd6ZeL1RcL3qjQsZKWiEC0V
TbwRs4pgeVlAdkHadwj2X5zxLaJteNKPbq5r1pX3cI0UdDgWHj+Qba7c1oPIUokwpZN3WkwtlG4Q
o8oMMVMX01E0R9ZrszeNnjEe4ZdtvepaRkdIK1e9sP0JowX/m9hGMz+Q1zIaRFgLWAlez5P63B63
mcpYn39mR4uCOsHGgb+2aWR+cGpcxDzhrkv7BcC9cFOOxC7otNCSOsr4ygSuAZdAuXjEDDBdTWct
SpCcs4/3LiBIyY9lmSKkZi66v2emat1InUn0rDXsepA7KWqdFOFNXhvlMir9Wqt0vNxByensHI51
Nepr+oqXMHcEQbm4e30JSo8h2/udig/z96/fwn+e9061mkxaGIaL+Hl2ag20Ey+7rJ7DDT39l59i
7qHJ9D3ydjJPW0Atz6FGyvGtOdfCFtV5Ju6QsAV2APQgitxBQWZ44kAGleUe44AVqPuyrRcxRqMB
MNd7YGmnGEui4ZrLKPZ5gc01rIwArcIddlMzy4Hw17zgQQDizWA7JXzXcQsW0OQ2gpdxLlmHt02Y
wzwJwnV0D2iO9MV73j1S6/htll3Oj/RBkDcMIAaY1xwjTPQxWmJaSc96qQ2Ibf1WkLKh9rbzjbVH
CuTgBkb+/0bEa9jr9XITVXeij3r1Bb/1uz0j1KD8bjxUvJyWxUTg7+k5BtMVXL7fFXmAWksOHzHv
pgpEscjDZWyAxc3CfeNikaYGPFVBXWsfsVWNfSUiLPo7cegOtHHwqZ//dsST4/ZTbiNyIZsvi3LJ
30+sB0EeW1m7PzutdqTb+tvfnkg9eHvzmUur4jxUBU9ukPBKuEWEQFDGSXAm74PgguVXEaYF+bmo
0rCxm5KMXt9q1SxyyAN/oarykQ3zLm7LrdTKsXFLc+348ZQrYkRH431Ezt+uLVSeVkHscKup30q8
Ik7OQWLZEeghMIodrt/kubTsB0neLdqnLbWOsM43tQrrqslj3g+9bCsLLltuOX8TDKP2Ln80kZJH
VDK6QeFI3V7yTrW++n7xR7FNoyEMOp+R3ulMTHYdDsnNjTiS77/F492CjjmFiSVTYC33rK+5ZFqD
7a8A74xwApYX9VDq5nEBpPD41o/7UacjH0tEmJUB8LT//csJssjX2Em9YTLGtpFY3tJEcxkDwQLV
dxNWGeLmAWXn4w5ozdxjLvyT80ROHH0V9SMSGq39G+RJeFmC1wQhqnI+wSftvpXHM99qfT7L1hoO
6kxSywkwBPz5vrGrvJ/GiB6uDIbQ/hmPWFzDxs6kqCbwKn+qp/87CHb2jk22sxlhpEMnSPRj64+M
piTZg5tGkgWENjgOjOo6EOEjTdZSy0lQ0YtAQnZEIKG1TGxdpqTjj0A5Mqyl3rJs9Jv3Q9HdWlHt
axq/OyRRplkQpCsIc+LdnsNkZaQGePGNIEvLBpnHGd7HXueZMsUE7e5jBKMoElyovO0nGhyjTdFU
WmVGu4MV7nd5vMhtq9usDLRgEll42HBAojVdBOcu/AaLqL24VvMwU5CY8UdVlD7yCAr8o6irbtkz
jfYCxs+XcVOkS9OjgGSql1v3wmN8im+hBYymqC2no3+zqQgnpAJXoAAHuou5L84L51e2/lzAjjTN
2wzLW0aesx42dpaaLSeq9INSosn5nQKcqGK+3E8Y84rz19UrbuXZqYS7k3hCLzHjIa5gvIfizSGP
vv/uWFNzNWfsQOtIN5GlCjkIVzZjSwQD7YgwnEwLtAfcBq6EZJLenVJpspugR+KIZRCgs35PZbgR
YinumXbH0kTnTVhFrsYuKXbQqojYXP480nt4t/58Ht7N/yIaDOt+gV9/sQ3nDVEJVBDndqyBSGR2
i+xYppgVJA/Xwl9Q51z19q7GMer89esiIn/A2rAhfzPVauVLr/tQ2dXLncoimHygUPMnnJC3Y3Bn
1iH5L2+02wgs9RlXnXG7Prdthj7KOEEAlSF2cAkN1NA4wglcs6YqwPT8uHeEaTYxdZVPXCSbajre
37xpoVIUyF1jmTS5iQLTMeXSovF2dhX1ldY7pXu33vvUYo3mpk8ORGvAez8cto+LXBin63Jcmpq+
FpkuboJ7ALqnO7pBpWgGIh4AR/IchVbflCMl0BcFBYOaXVrdE75DX1lv8ajpyhjZAwUR4dZ4P1eL
usPZ8fENdkdTiXaBvFAaYFknvrn5a2/IFh564KdkUv/LE1u8+NQHpL0A4OQenH0VWqQXw2zswRz1
DU6zboGWJg7ZXrMq0OhFBdCiMUL/e+I1N1uibtYj024aU/kZzQgVTSK4S7jTLS34bOvoHf7s7ECM
0B32WPm2uNOa3o3NXe9RAWXJBjJVL0NB1cCgTrs9L/M+cRYMHKOVQLF1xwDoNaDYGzdj9+OTXdqk
iB1I1S8eYSAAizuTqyuRHxUm2Dc4KbyLpFZAjwta8pM/6WZjAwnXWapi45C4c/WZdgpBiSAOKAau
XTjUpGaj2eu2IcH94C2FrWbg8EeneM5MP6WOWKgJYlSHMmbXvFm5j9ZoBwnk8kC+52rL5OxF69gn
+B5OkGHA7uwKG47khHDhrQ+UFHqrgX+xFVivIIOn793nYW1+HVho4DBNZ0lcABAFmsB0t+yyW02P
lDEHOlAxnYeoIYJV+P1F8vpwSE7F7lCgdJASY2JJi+RDSfyLhZv2UZ6itHj1WkCoqgu3Vb5b6OD2
scqITmxC0vjaKJ8vxAr+nshbVq29aE3UXimNn/Ig3oUtg70AQumkwYPvWhdqNMuzF7LdiABuz6C3
aikaZYVvlL14S1eAEe9f5gmE6Fpsms3iDAph4BWwvy9s8O2OEiIpULNGJpBzivPk4Tj8l/miPbID
jOJrRGyJYh5pgRcnv34cMIGr3JCpZR2cDtcLZm9d9WiDowFb0dRfpAQ9qKN/3o1MnPSlICOD094h
Tz8nnAr7AwcmgbzlYIcBEfrHP17+LthZrax+UWaiNmU8fAXscFy4JNJ20mYM7KLnbm96GpXHTp85
0RfYr0JrNLHBGhvOb8K4DleKdztBLgCog7tTE+YqQjLTy7h9osHM+Hs9avu470xoB7NPgcGz11cQ
Zp62iQbCH00pQyBHYogwic3JSWdIwSJfZoAO6ZLPvTllcMvuZDHyVePDTCbziOfHrrWAxH8rYE07
Oo7kgIQn09gOr+j5lCZ2K485QPTS1aRx6k1hUiBzUF3PfgqxFrNBGWTNj9y3AwNoKTLPZ7bv1g5k
SCgencbgGvvASOq33rWx2lt/e3UgNhHe7ZYfV2bmV6xRpXhUifO1qxX8pmU104dAVcAjdbXYoEjy
Ja9Hkz5JhwhYvd/XcLjDx7GkOUWOFKfeT6s7XdtiUOQd+yUQ9iNzuyp4bgHKCYn5T3AJlG3AGEbO
+soMjLbwz7+GSG31b7PgJScnpApmtdSflTkvWfSvWjFl9Pt1vy3lxOpPpCs1Ga1hx5mwH4xahzLs
j1tnwOsTkRtTfz9NhI+7bfPg2dhbvpdRhiGxcN+GR1N5KxP4TDPSHbKxeE0UuUnfBU5s1BkoN0Zx
i93jihe87/nRR3He412LGpiZYCB02nXYJq2qr/wi/XJoHl52+uscznCDD9ETjtFw5b5dXIjAhfGo
mA0vkrpD51lI+A0wtnbQKoeeR8s0rwT/oqK8r2rlFOPZpBf+Ytsun/sAkGbrZ5YursoPqXj8DKI4
CGAd+co2DXc1y3rQVjKPGNShQuPIzGsKN1F0NUTVB+x9zVQy0XHZyIYh0WBkWkrcLy8CGd7R7STe
A47xtz6qy9LzHZ9DPA/HEx4UmTca0D1LCx5Uj5cRsjS02Bh/ENkHIhekW6wCYwop2mpHd+pEtIZs
AUKo9YjV3cLYFOGPBQaRsEqDsxRbP7N04pBimCN/nEv3nVkGb1XdY5UA0XoVbeMylRLzf0iZJJmp
iq4qfscK/u+i8a94aOc5Bp9TW5QeSq+HZF5llmcEoGYaz0qFFuTKArSJ4F4Hxu5tc6l1OpQWhZW+
ZIMzqN8RHUxRpcHwDnd7jcESLcxKq1d9pgDqvQEjXghvap1BOeV412+N6cG0gA7Q6T5pt8CL5Pw+
fEo98n7BlrhiVpxyvUFjy1C2HJcDWig7vodKBRbF30XWJzuCxjkrX2M/gLxe7FSNRM2CXZmvzA2d
TQR/kkQh/YheyzQP7P326ftErFVRzXpD4uvSfh/Q6vFs5CPX55SdgrGeo2/0W1BURDcFRpB8QXzH
kYBRZN11X9xr9YWpqWqt1IkDJIH4a4fD+/yHn91cd9lCr+5H7IJzAwNoKnWo1gI46a72y3Zk+Xkj
3Flmc+WDzSmJfsWbHwcmho5r3zY2NmwrqSLsj6bk3e5+WRe0P+mgtRuOnqtr7MB+Bb82x5dAVl1r
w/zedlDmVD6MO8ZWq3/w9NTjpadaj4UQEDixtkeDRvxpvukUUpMK0KpN0ffJopTGEwUdHb6CR+88
+MbHATtTJOpLsah4/1o9/ia7RA2da6o4qdcx/PmBcitABplHt6DF77gmk1ycONYfhODjKx0ppFLi
t0bQuBAb0iZaF1B5SrsACB2+W5MIeZIxeWtbeNfopAbU+lLB5lInFpg3aSSDW0ZDw9CtcDhHyMy1
ANpTBBoZjH0L8+QaVO9XWCjIwDnDFCUUhVB8BUdKXNYaApBby6HZGF78N1hHp49FQxHqXRfN2tMX
/lXxHWi/YBDAUP1VdvoDATz73d51BazU7Xp5JMXGd+nS0upYf8luPMjcKKW+YcWqfsMaOznW4QlO
7ITN+0JoVVCixcZ72DiKg161YgajXt+dTNQ2HGxHrd3JZjqCCiYCR0VCSlLLhub6JHmLPVNnW3hp
JrdEHSapgRpprZmK3tXwNOgo50t+KSI3C11SkCqgSCFCDWGcoyizxHZeQzjCpYyLXpjq0hOTNeIB
L2RD/6MQdhwHQDPiZh5SIszWOokJJ23aVzuvbVkX/aZXljMTEdel49+sKU2uMpIGHjEbxEGTTMz+
kP2thKJZ8+pm9zzMcZzx+EWM0z6MPDYP7mi+BWVuOmMmODur5Pi9DR7e/CYo+t1FPHsp6TxxWcqa
km+0wQzdd0taA9nLZWZYAqL+vMNcQmaCftJBGO5Bk0QrZHR5w9nKLmBuXUpWOlKArd1APiYduDNa
6zPtTSGDO/1/j5gob5D/6RkU0dXk36sp+CuiGs0igIkTdcQVZBxhWjdVHQiYt+G83ypU+OoTb9xP
sJ6l8ySN+0FhZPHBYw6aEnEDswCZAUMIAt1V9oVmW9r7EmWC2pk+HxixGU4IQVujieGo7rZj5IpL
NTqWpzB/DO1IH4HSP0Xwawpxmp6Bf0HHGb7oe5PZ/y2PHPCqtgO60jOZXpEHUHBMKgmINNl7uZZO
l/0Z3yJ+GykmCSS4jGylDJv9KidRur994OCOTOwFDdDPq0fccwBSyhnfNY9oDFryanFBlaQ3Yatz
fyCOOBn3uxdRKA1TPn72HXgrXwnWlmDvI2yjS6WSIXUJWP2+0Tqpkh5sC+SYbiEcwNMTocKIBJ3s
V0QtokDkb+uFB7YMz4OM/+6S6CQiVugvKPaFPtojhxdSP3D95YPMXWhuc4O5l9Zq/tbwLs8Fso5L
Kol9nbPZuZ7V4LH58PoBhT2Da6DYniAL0ewTTBWBkj6OMUBXq0STT+v+AqtRTO0zrN0t8xrHPQWc
kVAJF0ZBXwrMC2xBwAaUgFrk5LLlBvk/WaCIv/OBR7jydNWJdG5E2efFrtARqut4CuU/SU1bBNpN
yWqUaLNWnrAQSDGzjqh3Y8ONKbZYzL2nLTxf4muEVwutW/1Rif7CMfeoacurcjUbHsvVCb1xhGrA
EjbvRT9NDfx3IlbhpC2ppjTfbUV7glC5BZ2WDvu6UjmdzFK+JZ8ecVxIB9O5zDOdsRFnd52HvHVq
a6LPqzcKtNiGl+9eCBUIaiK3YojpXqew9fHAgubdtEJEtfpHdsyQQ0nnYrxEHPPSUfS6XT4JD5el
kPXEY60Q/VuPjkowHiRCJQ29UUSS8N15lAdRp2l9+FPG9q85Nvk4pwmWzqkqIp3odMG7ph11NMwT
lfE+ngUI0Yp0Kxblx+BIy+Qpm1z43SLhlZPkzF3M4R0N8psocb9wDuCWpU9cgYZq37baXpcOi5Lg
cyVHUF/L1tEWu8c0d93LgtxO55iidO+XWT9cTWO9seu8TIOgTX+1+JDljHdF1Hg4mJSeYgAeYUpf
FK3JY8cYVeTFEMPTXXywpaO7uul2FPws7F8fwmaOZV0vc1gk05N6e9tPZynqXFS0W6GMvv2QJfCk
ojRG7peaki695XT99HxbCZug9b5+jVZ7pcxIOeqLeNAQy/tH/nwX/QBV6lIh0lc02GivtF1yOHWk
ZMndQ7dEDMIOJPX9ywHnSrMPmEWf4r2SkIGKpw5g7kwK+VIDFpShnXYx6dcfBntW3ufq74qKLbf8
JB7t9Deo1eU23DOHAXhTpUauruqhU2np7KvxKfa4fRK/w6xhhisJv0ZgfEMmfbCn+ifym9cEepQO
BL4bsVgmJaY7sdtovgLbYqv6UL10Rut8AWmcfHQw3KOnKyd4RZ7d6oOUvlkMfE4ExHAdumhMFuFt
SNO1DtXnIugWQCjhhubaAsOTDjEiN6Tp+5TyArk0ULyWSuwicSjPqfpSW497oh6K9y4+Fw7VE3BX
zTUrHNi8fCNQHuUeoZYTINCThdv+soePYZa2jYvNpLrkhxCR+4zjdt5reEa7bLJ4sZoV+9ydZmE5
FX4hIERHod7CqvsNtXn4c6qOO2hye0eJFa4xN8ozuxQDo1T3TYo8sAmuU0r7KbymKgW7mDEpFkJo
tGj+plJEBhPWEKoc/g0Eo/TL14pN796GsnG0G4e2J5hrZflRSNLmECTZkgZqNjz/FxlcVOQNCQYt
uzR3KHQuqFs6AEdSg8E2abLTr0ukjE7oYki9YdeZfV+DLrNhsPJgGVmCMr9d3VyGUefgKGBTN/YY
NlqGgY47PUYwkhRi4pXVRYsMMa7uBHlCmIZO2h5rZh+YNEr1ZOCNf3r9BY9xk/70P+zX8m8cYL+v
gRCTFDF1y75FDgHArA+SUS3p1E7pd0f1yLKQVA/jZ93EUHj/Zo1hQPdd9oVEbP3B63lIfXNCEZde
b37S08QVvDiulkfn8mIT38RytPL7UdHUem2Jei4tASf9iQrkxs1LLYlNrsE+wzRReY6OXx6bwMZ5
yuphvVoyLHqvjkZl9IaAr2kt3/XVc5rphRF/yPyAYOx4+gYxMt3P6pcnLKihHqkJ/SkSwnjJvC8J
F62nTB+wO+nPl/9b1Q1/qhB3SrFFaW1uMWi4OboYSYlkNDQDYns5MmSxf4M652vUSeMw+vlqa/fK
lai+UWfYko+WvamQ4W4E8OpsuNkrNxwyHkEWNwfn/HtYtDmmwTZN5AqD4vYcbxCdP0veIvdBntB2
Kc0Eb3rwZSNROFoUKtGuzd4vmVC9MiKZsTHGOO2S7dJi8DadLbJ1E9uOHVh/3O0q8IsH9rBaZS0W
4S1VcWnYEsNhrAyYU5ybK0f+kEx1q9JY4Rg32Lcwaby+d89oCYUzHiqEtVCMdklHdmIvvFh6EMLU
l6YooPN6dUcJLgT5HaTEaAOw7BtNTDM772fToHhLBmu6jhUF0SnHx02uWN1WwhjMx2drgAMXt9Ix
+6GF41IYHAI0fZJGP6zMUP3U632pS4+dppPVDu7vei09QQuB+CRlUn/82kjbBnBrR6M4DqxroBhi
7Ddf/+ktVGI9IGa2Y6KJt0oOaoV/5YDr8amq1aCivb+Q2y37/y3/EC8LLcPxBWE1vYLHLoQGPve/
50tuteHRvInn6U7wCDWR7BuwEfPYeMVrX+KyCnqKVgl4Ruo5kfmL0EE4KGrWUfeec5rJGkV/cGdU
IsZXWqEtLZ7+AMIvCKPYDakuFu+xQPLhhkzyQ46VAniAnzzRiTukZ8Fs+q+SzM5BwPMjI6QhhPHC
CbbWAQ4syQVrLF6xlwWldh6096/vg/LEUlluD0hJflXcbu3+AQGJezLLC+0nua2OlnagnUv0O3Ox
foz4RsBGeUVhUSNQ3AzWNcN8U0I+tkAUKdFCjnG7nd2qMbvpThHkCgZTCOCW0YLfl20/4ra/Nk3j
xsEQnpMucFaPiX/Bmja/NZGq1cE6VkRRr3phACkZrFBtDtAZbtAd/T/plmhSKeQviYAN9F794lDx
5/1+JrJMVozd12+nsCFSOq4TRwIev7oE9SCocq/i4dxvZyLOV7Q44f176sM0y60mmRwJIKYa4WP9
k0IYPSUGrd1yJVaheWX0Zj2/wUsLjv7dcToYuBYXPKdPouw1vWMoZ3S8pQqIQvu2vdvodN6PXh9A
azDJbz968w6s2NcxahiVOMaEWJ4XvB5LWjuQhYZ3omwDBSGciZV4L+LRetrTvOYr0xyjgqVv1Jll
vb1gm/UxkpTUDGNDE+RBX2yLY6U+KxKNT4A1e/Ar51dxp4et8MRWpuFdnC/jh1Fv36BqNfGUIjZN
1l9A/coKYCG0Y2TSZlW3XRMRJCA46c0FqcERq1ge1gGa2OQCI74PYg2QvriF84av/JVkzsaSXkud
E5o2xvw1lwfuUiJWw/AXDkX/e0o6Tb3J/nds8czzXsr22qP5SELvnS9VmUJye7qHAI8m6qk12zDp
ijxIvNR/sNm5bkxtXl7PKER+TmT+w2jygj1wTfmLmvgJg+i+e4Zqy3LROV3pnPsq4lb1GVK7fGzV
zCq437CFvQtd/dMNHIe4r+AwJD9hgClGM+hHv5l+mO+uT0SrzkDZFYVfWsCwgW9gp6J+9z6S5wVM
/yET5yShOjaJAl3/Z9WW2PuVFCOw4Q5RISHU8yu6KWS91UfDl0uhLBmEXkKymXQLqzYY4LlPIm0S
96+9+zTIR7hSYEitPpP+SRW/oNK/MezAjfMv4uWqrjmH1zkdIifLkIBa21Lvfzj+9HjPL1flyLjW
pX2arabj/ybY6UJmBkAFW3XCT9SM/djp6vG73sUGNNk5AIcpaw2Hhz9HlnslpaoUpbllpr9Nvvnd
dUvGRHuWbfOkTekvMSr+Q/Ql7BsAo7lV5RHchh5cid3FsiEVGepopUn89GAeXxtefvOERnwo2QgL
PLLiyHFh297hDsiZB5uXdh/Ms6SktxS87AeniFFoNJ17vovqihVwwKCdUDKMCrgB0fYSpM5XurnY
36azqLo7sI8r8D0qHWGxeXxs76uYcij5UFQyvBK+1LbtEfUQEeQ3+RHrLkKoEKagthC4Sr15Ga2T
KVcwUGA6b6jSFb7vFqjLErbGzRV1w+PzhTOJ4PimfX3sF0gsY+GhFrnX66KIp5ICPW9aUx8PMlmo
VBaBfdSORp2hd8geeu1c/GivRZlW5zXJ+0Mjg7f8h1xKXYYxUaIH37X0ovoCKDxcQA/M03lw3e+8
RGPDn3QuZiFhckAMFxB445h9AKoLsxduLdRhUVPGF1LKmXh+7Ijx5O9vroQZXjB+8oTOlQ5ttD//
WeDmiC8Wj310aq42RzOZWe46+im29eEoKUMVJY+M0Q5O961FEP5dxrwWgujrTuPBne+2vjb9zf3Y
SL45DoV5KMUPOZFJENr7AJGNVG8yu/TjPkLuw7H453X1ODwa2mQYuHPz3m14qzsyIVKRXZsOeeFT
gMvN8y3QI9Lbn2TO84oZZbAwMQp50G1A8u1Px79jeg/rppUP8ABQwWfG92Bj7Ca1HCkUsryfwO2z
uC3+2k4jZJQllYGHtfMmnb8ysrNJH9FRJcOyUFpFC61Glu9aS+aDeV3zFXKYgGxWHsv8069kjxjY
54Voo/DN4VQHPeQJ+qlBDL+GZHg3j0EHiAGvEu/tq4A/PEEwbDrBMZ+ucaeX+kQVbQZqTIfotGBe
e6M1n3sSuYYcybGfvRVlY3fitNUXcvUABVTNCTFxkh+Vaf2QXeDkid8xFftjtkziJgmrGB+iNfQc
4vHKRSkEBqRyRKomlGup47BYoVA/dJFDAgx992SDGuk74+JYnGClssYFoyVWujRuuM8+0LFRQFa0
U6ppD69otA13v2NbVP2ueR6XL9hvobs0v1Fyx8joiNPa8IBDBJGuFKTRlx/lW2FMsWU90Zy+6aCK
nJxZaNUexvRTXju0L0pN8Tua39eXsRNoSSQ1b3cBGbKc/j0ryEzI1b5THdnEh35hoDZNkw+ojMl7
UyfMeZbXpXqSZA/ROX7Owi/9ST9IsShjPJFbYdIzXfzIRkZxUFt+u2Sr8TsxyCDRd9VyZpDiF+6s
Q0R15jqtVUzlKScb3XHfFI14Y65AsJG11yjS685PHGWYW/WMDMU7p0zYaLa34d6If8+ImQnYGd62
Q3JS92/90dlQEU9hEStgCDekWjHM500asV25wEam8A2Sd8FAqgjapyX8Gj8eLDT78UuUEoxHF2ed
tVRVb+2Wm8dzy5+uOinURLrYIYUjkLsYnok7iaXfnioCh+eTPHiVEe/V2Cv1iqVPnqGXd63yE/lE
Gu5UT2m+B0v1BpN/RypoM+dWuU63sEOcDCK5z3/sNlOP/eqwqiv05GBCs4bPWBQRLjVMGHZPZ/pS
RV9eHHS3F5LuebJTHzFHIk0OSR9BsPT0p1QlYq+bRSzBMuwLbxGDq+c81EBNFg08Vfi+9eMqLh8M
J2tmtWy9gLavMdwK7V+YENdmKCMhJ7jdIusfv5Db+7K/p6C/wNp/7wl2Dwfd9x/JDwJW5InEkrPM
WX6bt19JX7YA5ZTNI3xaaMrq1Cy2l7nSIeUK4TjIsCM8/eGeiacCLrvlmOfVx/qLltc6DWTUFMU1
7c5bd0T0AGwCt0cSh/nQTBRaCkP+VNjDfJDKRVk+Bx9tsi+tlbF2VkWXAW6YCIwh+d6FhERaWjif
wUT+U4S4t+7w6FdGPspE7ROrjDxj/D8+RJNhkg8CEPH9dqStxvpt4djk7xv9HFh87Urlae0t+AlA
fDgSYBbpYSLMSOjboQM9KgCz9osHBdLMgyPbKVxzA3nrrx6KOVqX+R21FXIneaAsVoReKRWCWFVr
LF6cose6vxR1NWTpozKUEKW88pE3ALiRtv/4UxOWdkERaaHiSr3f+dKbT3fY7M4VNTN5MyjZ5Bsu
SKHsG46nu/7J9pvWCJNT1SwX16fR0w25Z9eVy67+7uWNmT3s1gSDTK6d66HU76FdyQx37jrwOdC+
Uxr3tgo2tKZ/GfvXK9Ww7L0I9FQZ7ZktxKX+YlQ2Xaf7Tgt8nK/E9f5hGt0e6kDnIEGaWP59hKx+
g6wikfyuP6auFfBeZt2lnZGo1xj7apI+dAw/mbi2NvZLL44Y0gAdrX22V5KcZgUlqr9pEz5EvcfV
SkQY850ZC50/NCR57lava+5tyATo4Tjefv8IOgc7EnSD+76w8vd/vDw0Zw5a8ka85VNjBi3Cm1Ip
MfZd7ttb2CiIUW0b1FmbNjHImuFx/ZtZJuZRZsgVYbrYgUg9CMFfVAkoLGA5Ag/k1GSy8Sk9YseW
E8W5k7NZQYq3+OF/oVEZXIirQlL6HQLAkFOpc8An7wrwI95cm9pjrKjJp6pOQTFe7B7WVkUmUooa
r+Lt+q8rSGZQw8dHV2HuJR/emQXiKm0TDUtioAMVemLq81Q4DPp1bggEBpDssClA4hem6vSJ2pMi
GoIJL2muOO8FT5OTjEr0gPbv4W2ZdxzT++5v8EKOrG1z4f5MPujwc+qKj+1OqkF7PZdcqGGSUo9M
oN6l7QKOiYRb3guwLZ0p11gHn6DSioY7wLntSBvKwV/Cw9gUzqyLwz4nKq/07FuoF9h5EPhmq6zW
vTtOQV942YogPktBpUKiSGVFxUZjU9IvS3hy/AxSh0uleOpdTr1xY0PkByjCqjnOIq4T74k52tKe
NRmMo/1WThyIamWrheemI83CaUG3AruPOy+iabzDnYGCI76U7yj7+7jXDw1GRg19aRLbtfLd+Lmu
2ldUbSA3mC95od3ZJuNSzRYUX+2G43ij6+zy+4S6wX5x4NSU9FSHOOj9xzC4e8/cL3F89SmkJdNB
pND9T5OSyMaLbey5eONouxU08IolPfJ1P0noGZ7P6n5z2g+5EppHB3f+UMmqlJTP7Cb+gASp7BdN
A2IwBm+rvfZtCll2Wcko9jrQeYH1X3SJL/9aeedcARQDyFgT5CDzYmE5EGzSuNweL7N3P7U/UgJl
gTJxaNZdWEGeXgUUZQJQokY1WkMCmUFnepMat1sSF3KeWzCtwdXno75m2k4CqHHHwe+ergy2D9Zc
p3oW9fPrpyEd4CU8yzhIA0RNiMDHnhTnO0K59r0Bf+mz29Pq4YlzzhSecx4nUQE9N+A6JNpU5Ah+
5Q9OVJ3Uzg51z11ALG3GLAWX4mVqj/4ercVpJOoFdOnd+AlIw1c2z38c7ttAtKWUAuwzOGFmo9h7
PUowusMwizGiNEx76dah1rDrCguRnc0HB1PjKyZ3998DukBCH/JxtZQeBd2SsVaVVJcO8jxpIjW0
PXjok6mgMA7ypZdKKSWqNKZHutOqHsCZ9qY2dNoXQdC2JiE8/9JJrTywC+TpJGGCzGbXlRb8Kg5/
p1hsFhPIUbIjqEOY5jPY72ygj7yB2Ef9tKShCSa/888B+HZiPjxQFmwwOhsG3sxMlnBvRfkUGWgC
m4qs0OC1U9idBL/2mt1/fJyWEXDc8isv/Xb5AIocZLoDohDsH9EPNxGk2YUDolloiaswoLGNSbUQ
zs/E39u12a61JAmsqbOcN1gt4TD8TO8/kxNeVt7PjWmWpqpsWIjE1plYctbwnjFVcFUzNFG/8w5t
4BTqaF2gDLHDL/xsUoFhFNj/am+mcEowCd//u1kcxDA8HDRYYHFdQpcU5FmWJ5Nw5T/HUeVIXGkG
S8mZ0Y++pMD8Ub0PNfHMblgIs0q1hr5kUDs9yI6pEwQ8PYDTHPirLooefKqmBxnNZ6qcEAJ59ZXB
rJcYDTMHOS9thIkcMqeDB+m9TzooXGC/yNi6d8gl7kJJtnISeqfxzMJO9Txu6BT+otpwZN8/P/7L
wf5V19hzv6Jtk8UJjOVTic3OXkjbobJe2D/kS/ywjq7+iRkeOQIzn8plAe5SUHf6uRumOOXufEL6
XPZdVAALbpFcEtE1uyV+L4Vav8xAbNzPM5uk6oDzsAE/i+J5h946HApzz9opXDsvNYNByOFOkeOO
Se/deVUqCzzjFL8ugiphA2GQsq/OdHqflqBit4LBJnvg/d6nZrsv8sxcNRGtFYKtma4nIkaHaw9q
7l2IqvQOZM5q3EBwLT/WddV26PkKTDsDZz6YuwHa6NuPIJJOBIBcTPtEOLsPzEkssToWg7gtP+ti
LF6nJ+976VocDq5hyLmXB1MBlQHHy+3r8cQn6VLr4s/e03+l/yBvrF7WCp+YzASTL8YTxHI6KBB/
Mo99xS2sKFKUkcVEqLRI23MUe1S/vf4bMNnJpQIxMY2SLIModMlmk/eguSdYewnL/hRyCTE+ag6i
vFFxsfOWuwnrDLgt5PyWTu9rCIfj70azOSBSFC+YmUR65riYXKFg2HrEAUq0RJt6sSno9ZwQsNBI
bkgGyP8XXk1/t0UiRpP9T5UT44TeupORT8wRv0ijSkFcHeGinUj/VPBvffs5tynk/sGs8rh3wucO
FdXyckIa4Hho78ztlPJgbmYkYSWWJlpfuJdMOF9XcOlDAN7w2qcZ/Ng+Fgn5CWzH/LmKrEjNOyEE
dkyyVtQ3Ga72Q15Q2sZ8SmjCSGieyzEvq4voH1HDqxOMQTpaEBKyAnQLq7RyqDhqqJbFTtMq/5d9
AiSEWRcETx5fwmnKDS/l4JnYBs9pKvjF5gE8QN/UggPh5XSI18hhk+XP/H43QebSbhXhsCUBLk0w
mboqGPdn4FBHdIlA7HY0Nu87dsemC9gefRWIZaKiiCDnyy4n0UQKwXuiWdbsy+tTNgRXPeHy28J2
KGD3jqX+y8Kx6gGqrvxtQhkjgEZeiQIEh4LoIku66kuYLYSaEqlAW/yygrXzYOtrda91i526lcg8
NarrTi8zJl+0ZFjE8JnzFphcNxZyb/2kA/Xbyzbda6+rlY33kMK2qaRwkfNddgPRIEyH2JlqUgDM
NBWDBVcrXAUG5lHrxRjmf+Z1V06m3WBgOnCi6lJ5tw4LcDRHYyOiLxTDwXy71rnwhosa8z8JQbkz
rH3mSFKeoaiyGW3ImAdSHG2UI3KTHvMWVp/SpmWKYYx/2V1TEeyNOQBwH9E4zXkJ6teMkTPcEpXS
945LY3AgEe41vDg6cVPCWJBxVNQFVylbzgEAY89Ag3o4oyxHOVQre+uWQL0oNAvcdMaE5iLANG+E
qq34irDXYli95dfrcfDVCTlESUOT76N0GpZ+TK6850B1xRn9XH1seYLTLLyxAmC477dm7qAG+fF3
72tvNx+PJc0wPSUnFnMarfFI3AcqXBgK73psBOXnWrIhOJbrlzVgjmIp6hxTYqyKJ7jT3PlBIBUR
ycF7MWTultQwFDNu+Nc/3FyNaCZ7OQcRmiD1VOtINv78OTGCov1cikcw3nxj+gRhRNsV4o0M/urf
nENMlbIdxOMQsasKDSFlAJMlErDix3UmRXGYd0UcGY447g0Svom7FoIgVtEKOdhQw8fGKxQIB/Y0
HFL/9DA+ox3LeoEK1/dlElPPa485ZH+SHaJmxU/1q9KeiWlAjUzUp9gZ5u3qWjIdrB5wSj575XHs
G4SMJ9SscKGo3pl6pYCw5nwrh9aawgjuEUU9n53/zv8xIJTzwYrnxOObb9UeiQ831YTCOMkZfjbV
0jjDWw9etG84YIYcKEfVmBq8hhfp+Fc4Bb6dIvZrvLNTeGqSDHVEr6qpJP+cZ3dGrkGZ1nMpQCVa
HJP8GWbgYEZDSeGnZe5eLEWzZ50yV0zDgws5+HyfJqIbLhIANx3tARIrIW5uzsrswdCLNQ7K7QKC
dtRfXUaoN8lyaG8eyoMkUJuJtwpLANDXFd1gl66xTqV37SBcfOF6HvCbeDFkRYu/xQ7+o0cPVW5c
gMOdvUTVk1Gc5nVYjLD1R4Dkkps3hOWw2qUk+e5Y3H0ZY1ZiTxYR4w36Zi2ngdfuw5mrox+CQygD
6CPfsm1iJtvSA/CvGcrdhaBZWEIsAdJow/KvOdBCSovJf6cERt6B1JwLNkDSCKdsmPNxhdy+VoPt
FmB8l7r5DROfiu/yS14iZnuiPgMr6Q/9ca0Ta39f8HwPfyb+ihPGu4Dmwh6Wbjc2F9gI5IC6YI/b
VZGqtfZELqzmboPHNl2j1zNQqYnUKnSFVAfVTF0VSHCcUDnJqE58xvYe5b48tMDHoVE2Yfuomp40
kstXjx5j3+JbF11bJ09kbMFSZWAKe4XHJKtHTfD+H4HdpuMYkBW3oe1eIDq4ouVx37y7HGTR/PPy
S2Z/2BPhW1IWAuZfH8gtlcXvbZFeNTcrzscPKSSU1cdvcxj9UnKYU8UFZP57fVr0Kma+8uW8LTLY
Vyqc08VX5O9AxniYVecPQYEcFmFvsV3vIiblKZ+Cd6yKpl+Cw+EyX7MSWs1AAmIJhBGKU8WpOOTb
R1AJiY58xktZ3V88jb3Tz0wX9jBh5gFA8xiEmRgJR7S/F6NTEnH1cYSYQ75vFvX/hIO8fuo7ozvL
8M5sY4AuPceRnodZ1e8I5/nSK2mdM5c+MnzPvPaf5UMOQkiwhbOD2OR/S3L7xMSBTTRNXReOyJDI
fdva9jisDhxqAbc5j6x9WZTRZo6pDunknTU9jt+Yq50tC73pc0SQ/7IuTJjgwJl0IsLFQ/wipluF
JJ4S54efWapyCIS4VQRAKmz+frEFESP91LZCwNKQXQUywfDUoWGDjd7dJaYMXrf+MSwPSb2Miflx
Z4C5KZzgRe3v4K6PqbDN9CHpU0K+ICqtm83AKNtn1yP8gQ0c7hXWxJBRfeOY21q0IADadvvAphCG
zsgQWaIJaZrVYCm91nv78/OEmtHiRHPtRkuyBKWD4LLirkXaK0ggKVnWaTRf7mspLs1Hj4uwYgNw
vuqKPmMocHPvKx9iU9T07uk+YW6toyHLIDOL9O1nxqSqkYYEkHBXPS6OJDbFv4so9X3Xpkib5Tqr
Kw2opXFda0mccZRj9oO5yMYDnbA7XfH9VvRx01ffcwS67olRBUbHz/NdWKP4ObKD5TPOAGWHNKG/
vd/w/g6AVSo1MVnW4Jk5jI5iCDoMBZBdVFnx/9gNmRmFnheiOaMzbnMk5MY0QPh/onbjSYc3ZgWv
IW3LBEQpFfMEJNcfHxJOaMWJuydqkE5stJkggcS8HRvxYpnHANHhdP+ZWuNf9QDG5v46p0iI8rK1
dKAT65KH5wjdutCKS0JfNPuJK7E1duaROO0CvRKLdz/pay04/Umos4O/TAEkYpVfKW+cuLsVML/q
SkPQ0L1G793T3jOZT8RUMt6rxSs356GpBk+oFIVm41ewGNcf1iG0U8UqGgF9usxSZLI1A+1RE3S+
lNGZCVzRsGqiPoJFv2J2yCjjRZOgd6Y9SfiI+M/QKm01VStg3Ym2AljOQHK+/47zY9CrLV92etz1
Y1TopeciBVkthjCSBqU3Om5dxgi6OnN9439Q+7OsdfRbvkbRxyX/GLVZj8UXXXIQQSIk840tLu5Y
+Cb9m6k5B+7MxsSU3zkCSJBCJHnsQ05HtR9muD417l3JGP9Vc/ea95x2xudoYUqyhOMA762Rr/b6
6j3GN7cfJX9JP8LqzVrAmoLRfsloa5n/cqQL/1Zl8n3jNEfgQ+sXxaptbr5Tcwt2hv8ngLfSZGHb
fpmYvOYTS2LmsKopbX76hBqv7o1sCgIJUBQbKk2sF0wc7qr3lx+Kaqtec7urC61oroKa9FNzdHHV
dpp17Q4FpqtbLCDkaL8YtzZacZXUuuzt7EnVk2Jntk0+p7G9drJ4dbMQfLMzVYovWrGVjHfOFTKs
+ecxsoEYInQwH749BbhluIUZPvrQefxvLrocxL9s2+zR8A7rXCiDeDJ78pYN78I0XCgzeX22g10P
P5xFAz+neRkeL4cUqswl6y9Dh2Kbb9TDRw6A5IXOGkVgfdNZQEFwpON+2O+UYLhRN6VVJ/+iRt3f
nMqfqy/hSKfx7DZ6XZAHPEwkLbbj2FAXxW9l6PcDGoqwJr9D4nWpb6Yww4ptXQJri8BDGT8mu3Vy
U2Wg5mMYhl9LD/j7jPIrDSNzOfbsuZvQNZAARz3E5uZ9sn/ddPzS13A5biveme5NHP03s4bVYl1T
3GqVoaEn98D3YWa7EAFlafHPmki9pr2dNaxfTob8iSK4RQs/7GD97RrMMN+4WeZ8JKR7q5I5/za9
i5t5krCj/NX5dB8/iXdvBiwkCQ9KKW5vRVE9e8erYxTpfcOCa+9LBHJl5H/n2RCTbIekmkaYiCcF
SKeG+hy7srwQLBxqEkZEz50u36L6b53mx+f5hVoLC2K9k5mUw+f9cHrsfoG19N7ypKNa6jRmDCxb
RQosbn7uydSdGGLw1guxkVoRT5m8MUiqB/51a5/sd/jHMtXAEN1foD82NcYO55G9UmBEITc2fFQY
bqxun16eljNq/1rsmgPuDRaodciUgECJ+dtxlir0q+NJTO45mQXpT5kW6XBr+e68dKijl/jZg3MA
FJnnZXYwx/JRDSYq38QJCcZxJKr/rFYHIckyd060/kAAJK1lB/eWija1i9N82j/GkFec72d5tywm
TaLfk5rTxRUrRw57UFB5OfSqjaP0YXCF1GjeRQgmL9vlrXRvF/Fhpj6omSfoVFoIssWlZd5umfum
8AeBX1BQ9h7M6ihxqSvgjbA3hgUJIZmHePvCPgpSwkXtgDNMB8qDBrdyY9sEsEHgwEgevEfgX52+
D43FO4DFZDAvpgQRaBYBjd4wGlcRb9y9TC0on9mL3MeW7MHpn29bNUhNAvCBJzsT5w5vRVWw03Dx
NnQVzmQhl06N+0DS9ko7L91RT66CcZ2Q1956G/fCXWa0dd0lG79nqJ23010shF7IxDlATYWyN/Li
bzQjH4MCyzLSkMBT5XpMfMci+fk2w5z5mJ/+RmOwx0oR1vs/6aZuzGLz3qtydgalTEIPn5HnBVRB
xStlJjkpzAkpJBG2PL4kq1K4zyS9vNwFqzp5tUeue+SIwKwwpxjTutI8zp+HB07YEHeVviaurS8j
AAIrwh12BvaGSRGfQGGKSWcaTsWsEdP9GCWtE3vJ71tkjQhgBgINzfimi5P5JUSpVfUUojCVEOJZ
tZNxxFNM7EwYyO/VB/QRPtslDEaBL8RsrzSEBcGmWE9Fzb7jRhEcepWSeN8MkV/iRKt9leaVOyHa
GnrPnpi8BsOUBwY1MFZdn620bqLMMLzguJmfZeu5qaUR4LWXtuAXa9Ik8nRBWHqaiCG65VIfs4uM
daalBlv5y/nCKMN8RefPSWZZaRcVmV+vrRRIMDOqD2uPufMR63PIx139WxJisYEULJ3JuA1sSYVi
Bd9VJIWHVQvnKmM3tKoRdBIIA9n8iO3xmL0u+F5Rj7BkLSGbrj2Wqcz5plXIStelCtJi+PzIqwDj
Vw1/LuvRoUBrGx2JyxeijFy0ijvUGCQ5iHgJs+8TgIJxA4bAcWtcTL5LRzm9fxac6ljQzVGvLocR
B6SrQ6GVXL7ZCjlyq3eEdmHOTc7wTiYI40JpzQFHk+ut63VEl2kqaRew/OZTDrUrz6uoigK8fHXY
vLJxQoCJCcLdMppfRS4H1ymR3sCBE+ow8H4ycyRMNSXd3+E1AM9Y0Kf0bbV+wPN9QIbGgRJe9W+/
f9kOWjQasIExByJFoaEZsPo4ZoBprRO3+TJMOvDQTO62KG6p62kJ2mmwJK7uh+pgGFY2dDPClFYe
M+kcIxHKrVS/t4MARnSkYnSEiP+PDB2awl39VDYZgdFbfUWh4fUFgituJHByoqtCCzMXMD3cYyET
0U8VNNBqMMJjxDOFkQ4ZfsctBR86OaawbLUTS3EATqMu4aBexbTabbgSsj091P/KCNNqfHNwDWb9
2opLGn0LzDnokTEUK2VTcQRRwCCYVPIsdCWVWuJUQkrb36VtT/tQ9Nm6S+yhcOJ1RlJOc6fJNNy0
hqr/m8CXZgp+wynx3MBf+cLhby+Vy3wnK+8ofGlNfVjmWV8fBZ/S1rQSNsW4geUnSRFFKDCrxUaM
WIDo0Ts8O0Eo7IX3yzA6ED/3Ce/s9FGlcKAxTwj1rHCseWevcxIAoaeXp+Hj2k3dJI7JE9wYgzPq
V7hq9L/HTm3JUTRjS8EBt779kJo8AHHGGRJC3fh/ZfLLCTTaqbjygevrd2evGIhLmvvbFCInglib
yyUzhxOLIfQkl0UGtLkJtySLOvAJXa/iVtCuIOVRVX0SS/IaUALjhQKq5AMIH3ZWND0bHyvMvKpP
y7Cue4jgDVcyFJT7bfMAI+h3UuvLQfzfsXmWcX15FH1T+Z8EhyyG0Ya22eX2UgpO70wurOzxFksI
ih54VAY2nEAatQy7M4N46mrq7mfZpw41l389/xRXjKnjFeB56QwlMDThCd0Y9y5zSBZRjTACE5qO
Vu9vnz0NDKjOwtf0OajCSQyiKrXv1h2Uaai3zLrsD9R9+BwQHYFE+phsPC7waT8x1GFnwKrFg/Q/
ji3+1vfepv7PPCt9HcoqKz1j69VPFVQA76uYISAS1ou39de2hDURdFLkGS5DUiWxI8Tw8Vj3VSo/
l1CsDb9rs9k6cKhvajg3av3mTpcAgiH1UF3ISqd4fAdXr9TGN3kApzOnmNu6lquZ2wFWT4ql7xqA
+cuVGqcG8QuRq/o39UOgLSn0UH5nfeDg4NccPaygymNmWi5cyXBcExXSx6OXz/H1PysAf/AFPM+w
jdiChV/PgJTUzxsW7YxW3i+kK8ZtUUB+EeLI0g8qPibl5gXdyXwQ/Dzltb6mLucXCLDU73oqG01p
I+4mRJCRO97WDHym+CJASUwu9QT84wLk+yTcG3OrtfG+zfdr+xhioOwB06DtdA010jHtMvY2nKbA
Xq0nIJgD9mp4occPlmvATUMBCncaF8gbPqIogPIqptPXuIrofAYE/TS2ufCPVJrb5SU15PAEZMa5
TRk6+YwclKelraqhKkqeTDq3Hs04xacvcR/f965xRkHDkIte4Acc6aRpeueZKR1QzD8wSAQBbMcZ
zRxTUBDCIVKL4fZp/z2SCT9+OdhV4v6P4pNooC3lCMAHqYNKOwliA/+0M6/6QI7pNzG3uQZzipDV
neaYbHpxiwdcTWvBOFxG9BpHVM7Eecp87jRYah6fxFwDNY8zrSpBu/u/MAk46VwskVpU54+0xuaL
l/twZN6gT7JuAIv6XqJGHblWzpMyprH2S9omue6PsEbfBQMBdJcGYyl9PuPoAOdkR1y1WKaWf8uk
QzBVK3grJ5C6eJe/+7xQ+HiCIpS3EkkOdJDqUpcr9pDUehchfKdQM9PODxns6yNxmA62cQECVQjx
SoQTH5laWMqPCXSWlfLswxCWZMckZyvb+PEcQHiIzQkTSpTJNs9fhgHfl/9ANgsD1U7hES1VLjwc
YwH3GVypA8/NPR4Bzm5I9rdOTQU077XfGL286+faFrNLtxOIokGDRCVlCiOD/q5cnDzpERdXi4SM
n5SKOsfivyICmejFW+9IwdlqSm84lo0FfuXeUv0+bnnvS9IDkmr9BMrDRAZiwUIDuztHNbo1cqb7
Bab0FH1V1Gi6Fe29M6Wgo1ciahQpeCtrwnWbJGFE/nvJFqLEqhMMshZKhFA6f8vrQeASlDqFHfW4
r50wDahq+x1QUZcSw4ncxidSkjJuNlHOKR16xVTShTDz+SkRpqLzTaaROeXiy/NjsFdLm6BjIfKv
TlRUGRcPAgxUB2lr2BG5ucuAmGEbL5DQstI4Th5eNPTCG3UMQeVmxMLPBqMKndlmpwgTt+5fMUhh
eJVHyswvDW+u/1lzzesO4yVkhwnDykr+1Yn5hKhEmJUV5AFNEAGYkyYqyoMaIUQpCwuCSXkz2mDL
DsXbSZJiXYgHkeKYEc3NIQvlJXfr6F/riPlZffybsrmsBKBR3mLfxAgxVZbT0U8ccmOkuIuy59a1
pG/P/KFjffIGhEpPo5E3UZ2PVk5W7Va1Li5MeyJYEDE8PjSHJ4HJObIP2lYHtxswOUFDXc2RKt6l
uAKzdkAhO/qnv4euwoNBdnnvpLrgzgfjbuemfuqhXDzuE9K3KzWiYm+a9bZkjC/eTgi7zDQ8pt7k
mpOFgW1FeGGDoOuP140unZH61SLKf0gPJqwgREstvrpcCvFkxmCWcKv0KS0HoSRctSfOuCVC3gvI
/DKRajub/yUogQhiN34MzLSEOTQfXHCyY+v7KkQSOxLjiBO2rhhRn9vtkYln21V2hJr+gv2eTSQP
T/qpX8HTFb7mct9/+i4DSSU7fXJEfU6OcsZJi+ttwETCX4aoa8ulCdxvEF6eZNKCB0qDz0yduFBD
5BW8FvrGUQ4BiqY7AWIPBTvkWzhWnseRjbY1nEP0Q7dL4lgyLDuVK9zN5L9PkFLXRzR4d3ofP8dE
3vZlKd+y4hDWkCF0pLZNwB1XjT2SsUPGJUWgXUXeQKM3M1/IO/hU/f9uWcDAhhDLF6YW4DSMpdac
+BvI2+Bb2ED1hvSnEKyejnZbSqb2w3E2LTzf0jhipV7M5SZw6rGX9XwV+yG/06dIfqD2zbrMWSzV
PPkwLnuBvwxOJjokRTEHdyIiiFWu7Uw8rX/su4nExRfYgMMpOzZqTmA8BHEmB6T3U76DuQbF39rv
LYo3dw2XDt0SNXxMRAUi0RVflqzZi58CN/IlPWMOsHO4cmydLBcyINwR0hZTp3lT8vOo/SOFmLyS
QoZ01rmV4jxSOYzfnsMLJGyYR0dL9IUqFPLVWxPyxK42KPuZwEZPhHgU9g+wWf+rBUcPTdO6Ox1N
kkN2vrvkzWkbMdnOPocOIYJVu8D7j1F+tZIfkpSaAbC4m3GOaGFhpy1cL+KCNe7OFtvHSztzIO8d
KbafyEHlk9JXROsSVid780WMDe/UND/LS0wRqWO1TLXiL5pQK98iqb8Ab3laIOiQruITbLALMqrw
+kct+aMZCJCkQSqO/HcsZ3xewgwj/D9oiTHkzzwGQh6GdUIbpIU6RakigJWLnFx9I3t6xgJV0tN4
3sQpisEs8nT0Mn0ShCXlmXGY7MEK8zJJyilpCfE0njXjDFX0e20AnnXNI/Q4lkf8wLkAPoGNhIwl
V8lbWtAFH3kcXMZWP8oKoUdPxe9La48ayEtpMjTT6LIxH58jJ0L7r7eN2/DLvtINt2uGesTjNgBu
250pvwHXBApeQMx35ksf+K8J16LtCKOxIMcFvv4YJAffSHWOVBjm/zlNcnDjFPdlLbEMCiYaiET5
UyoUJZTAgPrZpWQOYBfx5YKf0R3j/KlEgj1iCsijifHNn2+FPl1i/KvkPS9ZGEaK3a1nQinEyMca
bcShXBxQVcP+TBheNUzsLHzLgQOPDkp0ZLTlQ1eO3SPakKOASZASMfhv4ORCZi1guu5HF3AWsKHb
iUdk187P6TQ9z+VBkM6y+5KXz5lm7hWYbJcTt/o6Vwrm5+5jWv9KJk4KJerh0kMJrb4R08REXJR2
fTg8dOF9sMO7T/kVOgIZGZrW3cYOomKL8GyPR3nB6e+FOiS+NuzRFAX3bzmMfZ6zJqlrV011udTu
UO6SKx0oV+XmHq3PtkwpuBqWr0BN6QQU1LDH3bmi85ICeHfab1YUwMKQwcLTcPgGHcFKAjINMpiV
7TsclIqAGX6oVW6r2fUaSdpG0JHvq5Gs7cHwFA/x7Lg85ZQv/DEGYJt6ufKODiKzD9MAb3bZldMx
6tJbV/V/eawNb16ANHQ3HaMJWNRUrKVjSnXLVDBLWkjygjJnK4D15OnCmTUirvfu7TaBiR8FAE6Z
b7c4NmKunjgEx11xnoqP+f78Zzpu/qZZvEN4wMwbFfiiQvRqA14GPTlFANNSD2Zk5fGrsZWwHCDP
8duWltuV0dZa2TXr9a0DmKsM4ZSneY14Hr9X7+dkryfypcZccHwayOwryJhBkHZbImq2pvAiLPSJ
mFpc8iO7P3b90gvMVXV7m5G8iCxUXysmGnXXSi30lZbET39pGbk72xnmCPu3NJTeRtSkGSchRqrw
fUi5R9rc2D0vp0BkYamK9hGpolG4ih/ZTJaOyXThSSS7HGTb5le/ApTp8rqI44MtZIJr8LZ8oke2
p6pRy4wz/Nr188mtU98KDT2BEopYED9Dsj/R/361D6TZ6vTmpG21qq7IYReTJJkSOOyFXdlarM6M
ktkfolQoVYrkqFy/zVBcCrIgS5kOL+i3CRqsvqrZfofSALxs6zmT6T8F0HI2pZ3xcoVnfYZFHYBC
m+udZmYn0T/qUWo/thggDMx7JUhmLT394fzywPOQuM9rCPK0tvWt8+4F5d1VbA99rv3z/iEsUenp
24ZzsXF8QnkIftiGtZGUC7/x1aXmuaYZBCURO8g4UDa2PRUDPD/kDVimoLexv38Ojmd7jhWkHUix
auvGhMfiK4AXaLArge824RYnOQj6Z888KaRmV0Ldh4pZMShbodQ1fo5okVLjGHCkSgwRqWmmhh3l
DM2lyKGZ1ywaO1MIk6tBwILQ+lRQ18kKG7+UDPBu0HfRHxJoiWEAID/bw0TeVelcNCN5Ho9XVMGc
jQP/224PLj0oL7f1dkRk3oo9KZIAcoAh262KbcaYxmZHTdiJA3IV8DJqDIuL7PA5gEo9kjRMXdj9
FLdpmDd9C8Wo6N0OsR6sVfGu2kGgfsd6arOPUzdnzMPYAs0IsMuLh/gzN7OjzBP7STK//95VlxEz
f01pu8KmhULFMOzrAZDHqyBxh7WJmwdeFZMQpFdi4eJVnn3zEOim5DhOODAVsYe/C7M3oJvWX0XD
LtH1XQpXp9p7OPkdnZ0mjCNikGkwAL23zM6nnPGGYJvMAZJ5P/EDMRnO1YXCg1X85/sUaU6YSHK5
O84E0ILU9mCgpOJt9H4bThfp/Idvc3psQZ0OHP51n04HjbauhUaDIvZ3fwDQiwT6hRIFxsaA5Y1D
jAZ7Z1Gp5QV+xN+sEavLLf1iSwN8jf3MVV2+3jcNx97I3INoHzdUKN3s/8SM8G9rQgONvn6doKlB
T02xIer9fbWHo6WnBJ1ftU9g8iqCwZIps3H0CLTc/Iq+SqjpjOJJ+PN/WTytUb4d0axRo9mySHJd
VVV3F7/jmKgLoa5OCmD4B54BbO1wkJUwhjz42G/fzvteE6tWy3zgZviG8j9EfYywCT5eevRg5JbJ
yNQ5iYzmG0tDlw56fKGYkr3x1sKh+Lq7j8qEGuICbO+3exoc535ayMgijdU6voZj7Mu4hiN9w4fD
oZQfCY1sOmJ28FTwzSfGGaiVhfmE30n26bvziD/G85+s+7UOY07BX9rTtoqAxUMJhfPo2HXaBpKo
VNiCHPxLYcirEaL3uXu91+7c/MVYTiDdfyfrAfaLaxhPxAzkKWl1VtqO5Mmuy5BNaySKYMFyuLiI
Hb8GBiH32rXtvthTv9E+xqwSkb8EBiKoQnTQFz0FMMg1kLFOYQUZEN9rRB8fFV0h29OGxBI4UW+Z
EG8sJSGhi0cohdBmpjU+0FMip/Do5pe/OOA4ZsgZYXu+oJ34nBlwAJN06fWG8Br+Se/i76VOTGIf
8Xq4wR88uUkD+xOww5YqNfgVhp/BiW2BDLxJ7fd8BhPi3kneUoo1xPysODGhYo/8qv6fr6xxMPgS
WW2XPdf79A9W++Hjjh3fxMobTGNU5hfeO5Vf94uvmqCEZk1wuu9r2VEI7tG7gnF6iNvTO/i+hwVs
PZY9h1opZgjsZYmQ6boFqUWgBOoIYUeVXtlnnwdupkJbh7r4BejLNhl8eDPM2dnQgUK6C6TWx1DC
X5C9pG1CXChe0Snic46TcX1Q6a01rQ8UyivsmxpDP2PeMTU5FRb+tdhw9aOXU/SA7K7Dk+5IUw/q
5AqCRJq2wOvJjOhb0EZXoaOa35pM8CVY47Cphkz3KaNURg3Sm+aUfjxU/FDY+QIrVB2SZCabMVzo
vBfnZ9AVyMJtCUbf+xA9O9oGwlNjUNVOP8eZ9q5ad9Ou1UozBYCFchqd7uavvQF5YriWAni1A2tz
4FVNw0o+yeaT6ZXLeMbALOPOMN+dLOe9OGKbg7B1qevARyeUxkYRgUKy7ax+gWkwRfsTLjzc2tCb
pXHR6lSezzv4UQ1Xqoik5RZxOihpY687kp7kDlzlU2Ue6I6nfKECiGQcWsycnBGo9Qp7hRczwXTG
FMRbKGsvUz0hkkzSU7N8V7uEK+r7HNZFnpXU/lxSn+5BNAoOrQV+d52zOkDSbMNrUh5FgpigqiIu
dBsCtgii/LTfb2qeBOj8dzCG3IdD2+Ecio4H9ynTx7e078hhmh5eGQDXkT/14hAUHU9yAmdAz/io
3lwISmSvQBte27mEDHilJ70EIA6WINtsJYkA5g4nTte7Ij2KuumDBE2k6wGQyogx1SZbTSkYEggU
D78WhNmisExBMzvC8vkADWIg8hWg7BvslUABq13VnI8JFLN5UgX8zX/3TwSyV87r5CqHD571tn9a
knBaFHSni0iyjOEQr99OH3QrLS8BuGiWCJemRcdohZ0YtvqZYCBGYpIDeBiRTxru4x/BR8bht3j6
Q5FgDQejYQtrQYCquXPvwp94HHIvfxZZ4Mlk8Omu83pp5j3ea/ONwr1Sz6tYYVzoQyQuAvz5w+eE
gkD18tQVXia+UzlG3ylDmpnYJpOkcaVHBT14Z4hm9a44NvklRb+V8coJYnppvaT7DF7MXhT45Uc7
JPKJqE95dm6By3t2nFchSPkv+JXhl3I0/gZTp5y9rnNru+KK133baoxpOx5JmauNmFNVuFEvudFo
MaMkSYPXSAJdL7Q+dL7b0+SIbEfrKjDdDCSRU7zjQxXb7NhEUGmmt8I+lMCnq8XOFstvfojAcLLQ
bGkNzBPps1DvMlbajpbqO8aiHxodhFZyzROQgey54HveZr1NisJ2xxwlNiGy/o4Uj+uyCburn84J
vty9GvUZSZ8a7CtTl4ErIcE9EWuNACstS98TzW2dZf/KkC3lHHA+ag6f5849uL6Q5ZfsKFMQIYmM
dW5DK0YHm9FCr3T62mGftHMNPQSEoDtmEEAy+qAKzHlFwyAx9OrKLCE2Nmhz8a/+33QnV3vRx6jn
qYH2rIJleN+Nlxz5AO/r+4TonRyq22BqAOICO/YGgzTY1VGyun91/R9teKq8EqiWznr3QrZHTTY8
XWEzsZ3cl5mR2O6CNJwijusBUfavdGKaF/28pkaklI8lPJvkQNFIbC2T2kSGIiskv5J6JMoWTSi6
VGfv0vfynitsQw8eq3Upy3avAYnQwXNp5/7pKdCQeEzk+pMPDR8v0nIE+N9ZYq6ldAvFZld5vhCj
zEJm89eIGKDt695O5Y/2o4XflXozHzrKiNda+aeGulrItZvHvqMaS5UNLlm0QLTWgyYwuY0AKlTc
Sz11NvuhJnaCDj0oJ36RiKXsD2/u7G93kYkubzVoPSeGOVOf2OW9Gw0RScndCEfJbElJSyIt0BOE
sXpev91mSxWuG2KFwz2GLCF/+lM0lFuvzNMmLErhAWJxBh0bsu1MLBzj+D9C5lVGjOVVBxcfOPO/
J811Zcs0PjshQFCoyWP2+701vDHVfxUOLRUy9YWrgtTrRxmgx/aYxdJ2B+F4UftO6Sy1bNZwsOKI
UZKVjPs4I5OxkbJ3rcoxdkKfvxDP9DAAVeI3Ia73AOiC1t0NNsg/KOabhGFofz1vNA3Iuhe9ojSM
P/4Exngtfm7VY9Fv0lWTsYlIEkS4nVeNNKG5nvdiIDYEMLLUJg+AHC4cpxMPMM7kvMw0hwkljaIe
o7QCi575n2rUCs3cm8rvVqItQg6jRliC8bs0ZuMp6shx4oQA7qR4kJTYVr+F+PbCR01Y+WbWScjn
eUNnn6NI37z52vC1Tmc94d0fnjGgIfL17QZO8dCPQuHCKOoGRh6xIBBdzQahr0Y0yoxNKtxqt76W
/MTsBWm3dJDrjm37LCoyttEGULhm5BvqpfSS1gcSaq1dY02CWw1FAvGP2/vlio+XiezZZHlsXT7h
GcHMSRz3MuXYVVKhP0zbhOuRXt+Znr0AAAvphRi/UM0g9wHhM5p7R4DI6vAQc1mv194BXlCc4+0O
ZOmBGTGiTSmcXR3A+ydRwNhiZ3uQ0O4vcDA/piFikdk7DF+mJ/IZUCgFgBucfveHbkBfxVxqwBrI
+GI/o4x3rhycHFNre8PZFX+1P3UYVhpt+gIODmIRE5qQw2asg6/uyOLhu2FhJY6jGLVXnrowqhXd
fRICzNJAYVqS/9+aEATBMJdbfFL0DKn86PqDCzDzT1Shc/lmwR+jFA7eXo069ZsM77aB+Z3PP5LZ
xj/SLX1sFOtXeqKaagVHw5xOkqEBwD0tuTgWqGvc6kYSwrk/+0ov74tz+xuyPqc+EmvrH0GYqXBm
1aGYjTeyvUziHgrBITIATcvv2+5yqTJbE+QMnAwJWGxRo9Ld8LxMELnvrgH6j49tSZuzXk558M+R
v2WWHdd9wOeox6aCR7lMQT1NeBqKNoPMS4/IPTa/gWEigXTIPycFXHLvQC5KLQAb0qVpvgqjwd7h
mfr04+sqyTmFi04jUnidCqM/F6miKuvdy5fe9ggt3oRzT/hbSXHQ2gWlh/Cq3A0hdIpB0kzOEJtq
8KM3tkAwpTPsfM0J/o521PLuCIwpgTX4LhpqwNtwnk8kFm8b8Q8IJRklU6MM6F1YLb3dQlZ+B4Ml
JSb0Qv77VMGmgUEKSHCRhJJfmMT/3m0ka+/eN7uqOeqjXzAuRWNPsKx6Jp7OP45wBUVzVwVClLjP
31Vj3SYuZmXSr0UWhJFxrHFU9vLZW8QVmydgpxIrRmI+kgL+R1FHQNlCZWJd9g5TZcqxpy461lSa
tNN5LA0Z4W0aGMVcTYU7Uc1bzlUbIksI8NQmyRs5eLFO5RYKNINWZQNbwomFCVIJU8T4pnl05e8O
zM2teSYs8An1bzaKXTX4SDSb/xDNLVe3zCy30+yhKeCnfxTVltHkRL3bCb9q6dYDxaXQqJ/UPJxx
X7oSJheQfzG4xG6WHitPRzLMFwib8Y06YeEygAFdxbbBDdA1SidNs+onz2EfoxWHLfZWwm8FxG8T
ov/oCA6CmSLOAi9QvrtNPtcfmJFYpgrimG9J8XsEEurtwF9ucDmrAB/jW3CoqnxhHZ8r2wqi3FkE
ORhElAPDxP5CRWKjegT0rjpoqyg9E+4NPVSA7FM35lnbrYIeF94iX91FDsvsMBHo0x7qWJjG3JPD
EIG+lTS9qIchXVHy9VQMwSBDVAc5WxU/SoCanI9j6CXYQiCEisYivRbIgAmDJxGAtraB5bhRL68T
Cca6RVi373Eh0cj6RNXZSIJfxtm9mUWPiU3LqWxjU5JXTRlycRYl7AHVHm03naiIGxNnyR3gh/6P
xlqC/Fk/Q2NsyY3OZ9JjZm0A8pMhoK8gmno+crY3xSr92x31uQH3nFiTwNYkndg2UPMNN5S/fMV4
bxD6zlFXKAS3Fv2+T2i9yHQJAQv/szxWC1nZ6t5+KsRX5WzZW0Sd2fYk6G1CLZBnIThXTlphJPOe
iTSN/fgYySopLMBdDgz/jmq7ayu0LXi8xa52Rewjxnw2Yn0tRpQlTT/ZWPRaxFWmT2BSctpYH4Py
OnOvRzWscaEMqN8VWCpw3SP3rBh+dRjKiG5naotA63kbGppNgZrwAXE2u9V4GxF/EVC/Nj5Qw9Pt
bzscW3OmvtPCQKUKoLH+eS5VU57L+iT33fx7c5JFKDr6z2tIVHnKgVJIfEZ5PyAUMrnLwg0UTH8G
FsdbQGHV5VLumfiBE9t+05pPo68ujE/FPVm03qcyHOJ3pyAXAqZDX60aty0Osza58W1BZ+IeBCd5
8uHizndOwtDB0Od8hryDCwqKJzRfO2ZQuIK050RV/VyMQPo6D++9T4C1Yr8ByeUas2RpLN/6e3qH
bEA8HGi3x/YvAx/W0Pqvayf7EqgmMT4IRanNgwqHWQzaNJBfRNBLvz4oHiVZAoOl2yRpR7BYUPd6
cyHIlAxhD9clIZV5tWbMZX2qUaj9iMGurF2xyiQdqe9TFtnFzr7ynH8gzjtYHkq4+Fd/YHBbkO2H
mBC/RkTYUuRXaZfhj5uY8V+6R1MtrIH0vd29Fx/65GD4ho/lFmkfcc1oRP9v6H0k7THv2iuoIWq5
BgeFAWUjMO6O56Kesw649xhiHvkUqpvdOjm5jNIEH1TjB1oxjYunX5ktDfcu42JmPRFRIijMby9G
KfC+GgzPOhWCD/CJN5TOpr7L6p5OCrGMu1TgrsUOeRS5ectnZjUis8lCHqvAiGkvjhmMUsJ24BiA
E5aFe36/uirdPnZZAwuwoJ8sLo2H+2aQ5QNWF/z3Jk1TMJx8lbRztb+wCOjrGOvFPi6nwBU2ifny
G/S/D/j9uoAXo0NZhfIj7FsrNqZK8A1rxkNg95O9Bmt+YKiCYZ3rdVZEwX7vox0vlA5S2ixal6+Y
yE36wV+3obu+JdIXna7nU1uTelgN7dIJu4vV1mQOlxVaJvFf7aXqi4sB1pDxqBPMdHZJjO6qRw4d
X4Ondu+OE9RyzstOYLvL3APeW2ZIyCLnYRCmQQGU/i8xkTPj9mvQsuNxzbHsjliYMQRG8fDR6Hjd
fdABZVZO+m6t/FjE75iAgoauaWi2e+updAONeVm1NrTxbIqu5z5kRXqWIEG6N/VT4TuVmIlj5RD0
5JHzGwvPv0n4SMUmfXUyg2PWLnTZYegqovQlLvHUbc3L0zM250nBj3p5pwodOMyLBsdZUB3ZHRi4
iIIffLNtsizzJYrcciN8J6UI92fVsGxprxybipn4YhaFpJzrUwanyIj/Vb+MpjIFUdpcxmz7vQWr
Q4CMHnKEF48BIcNjtDTgwuFe/qjB5eebWqEy9+y2lI1Uol2TsiW4bAJ6aZZfWTn51lBAnC5yYkqJ
mKmxNgjuZttqsmJrISNf5uEIwRBKg/XFID1vVWmAUDYkXMm1p5gEdgcMHFaY7rr2uiK5zX1PYmH8
JH4LkwzXjtaXSvMhX0j00p8YldMDC0EFFgiFZsouwgUxTW2dS5ktMb+tj5gAwegXjWJBE9uxexwR
p5m7DqR+hDz11CwsAyPakLoRTA1pk7+jzKvV3ZWmIIt1jyFqBudf/WuA8YQCZWwh1ivUrgQ2U7cy
cX+VF5iJjVQ5m2PamblhQvRNUxr4dBn7FL4+bh97bjM+wh9973cr+q2r+le6GaYOlAZZjRaem+N/
byBV347StaDFRc3f25rOkFC8umHLy5l0ks9k5KnEikmj1HKcrsjvd/2xoCXjkkEaU6FkFY275UYV
EwhyUOc+KV6saTYNybBxBh3ldKUqd5kwllR4LMYLvDTzGXYLj3kjBk9RhxQkYLAr59jzEKy3juBM
hoGThuxP8uFAvRQaDdtehYcLMJi2ablzrry4NWZRHdZdPutS9VQ43D/C207m63Je1QgIC41+fkro
BkyhidO+pS6d943eBtn5D9Yq7nt/fsDHDdH7cqP88hzGacRtRR9rJxoanz46nt/jcWKBQPsKyFkq
6XL4EpXjNqfR24dqJxjrOCDA0GTnKp2yphbmBWof8jwsiuMfLShZdN3NOz6KBQBjztFQjNgsyu71
sjEJ1LUDpYcfhsu/S5K4jy/LJvQoycdLsOwwNOWHn5EQi+yQNz4GIHFWdgNX+MhQFsoaIkldkTYK
2gQuQKx3WmgwIjLgOWyuCzRcwSTELhUfeEuyqged/ueJ810eZvH1/zzlNzI0WOvcxbj+8yxFU9+U
PkWnG3hc6dwQJjSQUcMBZsbCmOkOVg13sEaN2ovVgxk3gKgZb4pPAoetCOBDeEj6koRztyjumRG4
NIG3mAbz/1I+G4B1omf1EeG/089w/mstXymrNOlaVoo1VTNH/yhg731urRA9E3ySGbrkU5WPM+gn
xAfmpYTqqRjFq3hfkz5631yeXsvQ+2KuShkEjAbiJE46cHYDePbQrvAQyMXq6DFQT28oO+w8FbQk
trx5j4xQEF2E0TOpy4q3MG0VhXIVGMo9BKlY38dspGu5TL+JCIqssUigVvRHmgFSitsv3ujDzdE3
aRWQRuk1MiXsPZkLGNFwciD9EbcFybKbLTfPZDTnyHQh0EtHLgbB3CzoKbJ9l7eJwxDAhIcqgdoE
FAviUQnhnDPz1pc2EAMlD6+vUpMa8h9yNbZNogVRwoRHxxwHEiu574sbChP2apufI08A8rvv1PPO
VdWLCYdRPDY2XnUsTYdHLuR/8gTpKHHSSUdFEyrQvyIi1M50fspYQd/0+CV/aFXTVG+PR5i2CHKi
0Lmrz+jgvYJnGsj3G12SFaBQpY8gsGO1ptDKkLUSRYFhn7WwSDW/G8mmZC93qSwIdXVPz6ah/uMn
YLVNLtbsmFvXgEvVJ+IbJ1QMk3fwVgcZ09IO/iJ2/NGIkF8QK0z0y7DLR0RVHCN9n0AcxYg2jW9c
PtWnmpeCCCtnMx2TdUquQ89ueXexjTX1/2SdaGNs8H5K9sRoSm/f9IeQvB1Ilh0GmVNrZc1cbFes
z33JQtOybE2GZu2Fr5/9KrdhL17GL+V097On19CrG1OEUFa6uJgNBUkkhiRshK9ZZDX6pi3JylaW
9JbsGtlPJ/hilR3uUdCSGOn5OAKUCewQ2oxnNcvhQNJgDmo7aNrO+yyGO5r4bJMdL0qxlRIDB0jX
8ftOp7+Oa/DCZnREyCdUE7kw8WBqqHHHHOV+/bBuO3AULEY5e9klMXTBPp+/STADiuh/dTgBronD
T/TgKYcWk00qP/g999GAspz5wL8V8Ga8ZQwF9RSSfdEj1BhvGgDX8jpRcGDfqquHDP2jN+4+yjY1
i1MJ6BHjB71J1g4dhHSYfxg9NJbKDxLH4Mvniiitc8Euj3++0oSfIDl4LrjWzG00OsrAhaVYZWi5
XPdvNhgdT37obrFJ72D/gmK/rLQgSNzb+7yw6M9lMS2eCnlFa7TphExRKQ9W2dxS+xikJlKGDcD4
OB/OmUdm0ziLhP6j0MTPqQjnlMMZVITerbiY9ealS5FD5jHk3XD09IDCO2OymsYfefzUhn7agzTH
UulfcjtCoJzKJi3mQ2aUikcmiBmjIzYiR0L/8PVfPhqd2h/kt6tU37c6HJbQRI+OUb861LLulLeS
R543uBfazM+ePl4XV6Cq0me90dbdOsZV7Zt9O+WxLELMYhCYH3RBO07crThwb4k84J571H4jS903
+C9kjNJ5u2+EcxQzZlNcCXt+VFdRSu21mNEC74GT95/YXXPbGq1oSb2WRFsjAxJANgoEyOzXhbZp
PMYUQNUFnp56Phac814bnFUjEhOnGvP/4SrsukKXIDUSvt5WZr2htXu86H8UEatCWcmQUiU6w0QC
BwbZFeCVXhmG1PHx+x7U88iE1Prsi9svFr0zaCA5KNXH2aIg6kBFbbPkotspVNiD8aKkhHqZKFq4
/ueeRnA6CyOedTYkalpa59u1KF9qGcbjy/dYJbMqO02fnzQBY7TwqqTxgKNhDwzxBA3utgCAqvyV
DUX8TVmsUxOc3Jo4Ru+F+XkYWSBsmRL9arXu+0ux009tLBhehMiJ0ysuNj1PKTafc5FF9tUSg0PR
SznY3JSuuyl8atMtA0MJyxBbIG4w45mMqzQEnCW4Zf472bNEc9ZJJapDzJoJBRkdQb/Y8kOeH4Eu
NokabqAUTHgaSSS4Bpo4rInhAiBaeS/DKmvRr62gZoiDDMmwyfJdrPe8XOTvZar7M2dx4KLjKgaQ
uo/bXxzm4qnLPsEjG19G965BZ2RCBkyxYZ5yEVeGNUNHP77oJBeYSAM4mnYo5sI0hrqqh3bbu1QJ
kJx91e/wvDPIo6K9eTvjeffTRbleLgEHnaUdKenn+0Oi/06y507OC+rFk0+9qc7k6sOhhUI1Ux2R
3rnymKCYG/J5m/bArCVGDL/xGtnvwzAHqltugXnlF+av+uzH7lwGXR/yMxyMG5LlCopVmPIYCJ+O
CKQRPLiuEz2CHkbog6tTQya6v+lmEAOl4tqYpke5ytVDaiZ62zCj+JzjTnfo/TLF0pGYBzQBwK0d
Sq9AYl5Vxuh5C5pD1TypH+3sae+x8LvuCp2FlCjcU7Z9VDIJIk0c/VKdRLAs3pVF+PyLmLhJBp0y
pq5hbzKMdkOkDVWUFry9jMuvT97pnNi3FiPCqYtvJomhzYnGUQ+zELMvLBupw/eNkkHvD1VXpSEq
6fDKcKSEdIWoDwXuqfh3yTyz1meKKcLcJKxqfvBHZZUbWIuXqOzFn0E71v5MMhZB5Y3M/WGF9k4p
ZYES+BVMJjubmnUWh+wLHf2Us3S7yMl2u6rTIZyqizvAW9odcRZlDTaOg9yFRMwXrCRxZe6Oh11B
R5I/a9OWK+jVuq7Xn6Pvehgj0w9I5Ymvyc61lzvjoGJ8+D5YYD1vvOa+a+3eHDFRL1GazXwe7wmI
j1Q/EkEKOGI2e12UoW/pptSz6WXoOr43j2qEYFbTOL9i176DbL4H6wC3QMmEtV52h1dQAPdkoT7q
23OBAGKKfh0YlFh6el4oqb90GuXKB9abhFb2/BQC5OvqO5ExtjvoH2iaorvxLcJ+tS1ZXRjVg3w5
LuxH4t7bYGCUDVhcbjF4l78crgWS3NrvILOzC48+3JpMGhjf6uQrrPrlIoNR1rRQCsVZbJvXWFDA
XuXIvq+E1B4ATW4Mr9GmJcPCVixy/ZcwgdMv1qHQDNaANDcV8ilZ6oltFHmH0BIcCwSmXL86wWas
8fdqeixgDpEH/D2Yo+P4X5hmEZzPwmIKQKzHYKd7LNmCsq4lX9Jq57XfLxau97NGdg0F9MW7WaYb
P1pDA42uthmxlUwuxDKbhcvF5tAPqLANT5F8fcNfwkbFFY4NCBpxiTaD377f4810anoaiMlKgRtH
Duo5uLbfgHT2dKkTlcLjHknLh8EKg2uFO55/066g6IKMGQgxKZ1Wc4OcOUzRR5fyfJtiA6+QbqP5
B6YF30cKZN0scvzOAt5sc83Z2O0BiAYDu/zwVk7rHx89M5wQpwX8pDFgonzOjNQIJX6L1gRQ++UY
CAtAIBB+SELRknuNfF6X/DXtZXqGEXrhOg3xW9oa11LGND8QKqIYyj8ytb+a+1neY2fEN0k5AILi
C4kUG+uw4m8tSPf70x08nGhrchL3lj01t3oSzKr50SSkHWRHTBnLXi4pR6XjwD9ozdKKB5zEMpJa
kurkPFlOJcXKH8K9HXKhqkgYZrtN1iqR0aVW9DQMC4CsqZ5xFbMhzt/0A0QwY9YaZ78d4JI6JvNJ
pOkA0EMoT/0pRPh3CcnGa3Lgx8RxQ7zLw4A3o1zOLJQ+0gLeYgM76Ue2H7buvbDZwwKBu9JmHmTz
JhyPTYhHQmoWQBz4EVG+ExOmY31/BOV93vq53KaJYfpQCiAkILn/8XCPEFKTfZDU/cg7ixgO23ZW
wdaXu1Re7Y4ioaioq6aheqqEaZsNRsRH4iPT3R5dQ1XND66yJmqs5th0gP6xbmOLO7UPabfftFwq
HHswvexWvwWwW1SZf6N79pcCPospxe1sCAqEsbFzdFMaI/olK8PTg8M4dSXUy/UUKSdlbz/dMRYf
g1Vc7Y0twkLM2cya0+6/ej37PxvTLQ5ASLWXX3PYzW0eCyR8v9ExtobftwF+yZG6UH222DzOBgDX
1bq546kme4cPjA9lwPV8/10A7/aIvAisoiMCx0vd8GOzlfxQWIx6zPL7uvw5I091TytJEb6K2ePe
YsZS/zObGQfcxn2HcvMaVujZsKAK0xD4rzXKQUdQt4zxPw6dU636p95F6ZlH7v+kdC8M68ODPG9P
+bDNAmqw8OFI1ihzU7qjFra9If2/QpV0KyjG+55xDjGtY5AGmHYzfhfXKxkCLhbNhe+4oxwl2/ix
EI1qmj7+vo6ED4aGFwFa/khXKYaUP7VjJiPdmhexpYD/EP0L5ago9M/vN880lh5gv09n72OHHNI6
8rrN8hBs2jZDEvQ/PD93C4ELP5FuNV/f8qFbB6e7nYdb37bRFs65kSgE0ueLmRUcPtA6qyIrmy4p
J5CilQOHr9edFUhKwPGpfRVFFPzFDZV3bzEFcwSrdeoobpqMHt7FCXK46dtg/de8pM2iu8KDMOhE
FYW2p+Eu75Y2N587yH0Ps8/wGFfXRxN4yXzTd2TgmkyU9s8/KrH655JVo65hPYVg68SRBDciPOcW
a9XwHr37N8BCEtN/gIs42BMpJPRSMReXY56j26tEDj8xkmng9r5BgHknXBfx/l9KfivXOhFNtNEb
y8ou0iApM954HEqtG2uqEigQEJspMo37IN9YawevbzIGFA3feZ4+hIttI4HyOJGjyd2lHBGvte1Y
a/VvXH8bCKST4DVBWqSKMnf6wnLHO7pq0GgOuT5HbIODKeAN1tEY9olp6tQlJUlIrZ5N2Zy+cMPa
AGSa/As3a4u4jZS5Djp8sIwGIfSdX3BiQ5Pe5hx2GIsRzDOCVWfdKS3GAganS2ZeKw93BMAX388X
YNABYDd44vXAEAGmbLRMh3oEie+lWZFzCx2l+B88JaKZzXrVMUIeigBBYmuUOWBeiuUYKVIhSyYT
xBRfKT+K/6Vl+XDogV44jLAmrupdqMuiaUc2XazSWrOhENhsBk/XRejGkmvCn79q+stgHcQqaWdZ
Myq3SdaPjb4aALk1Ow/K/57gAfx60Bm16u3pafhXYQJXfUD8Nq70ChkhUf0aDbHVT8bUueLeoqqW
A3yvoUASMVuReBU5U4maGJpuGCDXnRyBBC6V6LzxbVp/dvDyjZSAkNzL+nUzLz3pU1k6KR2o8T9o
e9X2hTYT2eiU4q+VV1/QlPsUYE4SBMKUMcPYmOkjAL3e1llyfT+pNjBvh4NzuIrCHesQ0v98xG8n
OlGy0BpuFCcfGfYiXutw0c5KiPhOW95AM/FpbzN0FI04jJ2CkBwIR/XyZqJ06LgV9m73DXQ4KvzB
vyLZQr6ojsBDnvfNhlreceK+W+QDOb2FElAV6QuSOEhzHZdLszxZ4gFP/cADtx/VR8NBK+TqL+/z
CW0ESWv5ZvGjpe2m03iOuqupy0SX5OJqt0chWiwzXq9a5lEw5iq9+lsNGufwRGELa4/xT4TFxlux
QG9Ano9bHxQoNHSVu9Zj/G1qvi8sU2rbF4KeD3WCkcNP6opP6Y3nbn1ZWBO2LRtNFdOhhnCQZKUW
idhauqw8xo/LUyMX6n4iYg/sTAZUFIhKiBV1MG5M6J8ZmMWeuQoFNW60uNeQAfGAAWdG0oGyIdv/
BbB/aVAwhROGxdQBSEt1hOGSIH7iqT+kYRFcuVVzIpHdAy85qJa7RiAEH911BDWm+khdvGsccS3t
lqGTYKSfb3iBk6bX7r907r1TRldXuL/p4nWRdYy/BeVIFMA6KJD30cd5OTN8vw11g+yFJZ8Rzr5w
fxoxN+sZxRTn64LMvSeEV3hmQB8HXbHt8xd673XTB4w2qa2K7FY2ymzLZatPDIqu4ROboREX9+lO
S6qYk/UhM+ZJ48sh5JXeDz1ipYwzqGQBbGpRCEuhoVKZ8xmIot0uLE/NwpLwV37PVX5Mi7nxAgMz
20+oD0HTuunCsHcQjGU8q62xgw706PrBP4HcQ7hP4niu6+3xIuYfdcbRMDYNhLqcwQoNic71Xg4i
abwg8E60Qcw/nFKkqwtojHMMVWCiV9zaqB+Z2F978GaTXdQEB/xfCj1wPRkau/XqugfFwLkXX6Ft
2Ee3jUM1wLOVYCO1+ofIbAuwgyXrOsqCG9qzZlFY81ZJpUYxy8HEQ6B+KLyhPTW1CpnaGlOEkw47
f+w7BlZl8iXwYZOkxwrQxzT/b1L5HjmygZv/HeB+YhTxCSpky3h7xI+R6RF3Gk4ROb4hiwrtLMug
nLEZwsQ6LUGBKHiskgEur+yLsoU7/Xf3AiMU0Zr6PbIAYx9HBw/fcNOiog3TQjU5DchJxpkdNtb4
vbhhVeFvsrxlxwD+aCtt90xtFkrJG0KA2yDUm4tTcuoKnNEhLsrK8/vaL8vzSKQbtcjIGO1shu/3
P7zNbaB25er6u55Xp9IeHJZ8BrWrsRpU0jB4DdNQWwzkbYDsDW92+GlW8jrflB+0BPRq6H7uouRg
5T8Ba1OjPVFRde1TwXhLu5g/nc/vG37smEY60pItxXMoemkhH+WxE8Dzf3S03a2V3fWjkyQ+xDQ+
QnKzQS+T6jkGSJzOSgo7A3jHyp7N8gb2JfrlP9pa7Fw+P7Lm3ZYFoKFicx0g1jaW4qqRot/xniUu
m7gkNwQ7gzAtne/tfYitcGsMjDO4ToklqpvF6HyVZXe9cFbUlLXU6XAIJ4sw1bXDqDaUFV0T+4zw
mt6BDVa8iXB5XqChAcFeU7oFgwaiNGyE0q1ayYefLt6rDW7EWuUJDWzKM0snBDYNnDS1suPC2q3+
xtLxuxqcdxnIIEHKn2FPqD7ghP7nGHw5EmCoknm0z2uplMZI/nC+D7uMJwZi9N5N9u83nlaZPxC9
U2SzKMAqluaTw5Vae6tz+jg791lctAkjV370keMQsgaUNm/0hD0y9ZUpADAb1qBI5edIh9wSdQbo
amqqFtX+24T65ECJ0/ChvmypmgiQ8QdWcgBA6uwHk5GKPojVztxkod0Tc0MVJ37TFlC0qliUtCU0
3ac4gSMvhJysuAtn7e9Z1k3gDxFLogUZeT0mnsJ8zp7yW1xPl9LClE1tNtYKRZDhhoEZYWlG0IKb
C7xIokYqxHjJx52CBhd0/W8E/vBOrxzhcY7AY6WEH0piOsAOrSpHEd7KgkKOgNzzVXbP6yhHv2qx
Cr5mlicRuvG3zU98mlpLCyuXuf1aKnHy/o/+H2sk7IUHYN7fdrcljzJokQU5YqWjDX2p/pOzXNjS
lCjx552eqZm468tBCc3caFCX+9b36O636tmQrRSbL1SDofV/svJRBtYJBoIhnmgOzgJM7wxuM5Im
EpIXzBcCFec4oHh1tVL1N7g1pk3H1g4QUrMwQYfPnPAXriO70lbTr5XkuYcEevcoT3wC9c2tZVRE
85RxGFaniHmhKCiKYr6vuEk1oZCzA86Uj3Q4s5tqS371m9xWtsj/3jB378wpvQm2UrJCj9uz0Rxb
Gbk8EFIXh6LaUp7LjHaHaqcDqtvEhZdrjA5v866Diaj95aePWOzYKYF1lPwaTMiLDr+iZugPRN8x
/r1ufrIoPpoppHPOvM2ATeUSxl1pVW9H2CaciVCIzG33ONjFxUjiDveX9eC1VCaBGzKdUtWzjsqx
RowGBa3MDEW1Ti1gtCIP8NC3cEPNc096z6guR4XUqphrRLVXwydNDE0KsrZWLcVXZX6wpBCRc1TN
5xkPcUdnMHkK72NMLGmWKvdMZjXTqU0jGscFkl5BLEWkERpJMoePW2PryRUl8yAuY15DMgUbS11V
oBRJTwc9EjPRem2JKhKAgrvtafvuGEDFTjJ+gjvwtHzqciRWS9n3ClKr4Mq20KIvX0uAFlaxIISY
YJkv47VQnnIVZnOlFUD8Pru6Fq8/A6SXb6YxOPwE4upKiG4MLjIDjoHJ1xxnBPbn5QdvqtVxvQwT
NN9XMUKBO4J1KcEmnL6u3H5w7UrYpiPk01iqFFmCRHMhKDJEhuOWRdymCM1v3glMSSY/VM9LzTeQ
KlPAG/j0wufeZLhRBSVK+ZCkxEwQNn+InXsnX+BpYhjCWfxwk2mLemLJLIeZF8A9RhfV0j2Pwigg
l8QhOTbdsIuiGu6cEm5CJkXIQqVfy3svoB3k35vVt31UDedIc9Ft1PwA01+kYsHTI1M2Jay94YHZ
qSq3rSdGtSlEMBQu/tm+7/JhvP9VvLx4es662J1HzMdPfOhd6C2VXH6sjwf1QBNmlp82WUkScagN
segcU+th7nmmRjv7MXiLqGY863mwq84SronfeVKVhgujY7C2Qsyxm30SZ296rRfQTg/CC2ZSuAOC
MgKtttlQp0wp6U1oydwRLhYj5dJUKU3nMtICZ9k12YJeb+i+SLsDzxdWihVnbrQHTGnpaDAqfgnu
TYNMQX4aVVHux+J+CyfO3B1omXUI43YZ7Q/ukvknOsdbquNXISpqUfisXhBGsMJncbtTqt+76DtL
iwkPmt9rmVXCXWjF/7QeZ3qTJHRjTimGUHLfVku10Z4jjaC7KqWsMPfts5uqsZRhi3WfrGRHgBBc
Nd9FWVwrY46RoK8hgs3wRS7ANd1xh9HcYeNLbhLjsks5j+xAAHWIbHlx2iNT7BbNs+dIxtYBIiKp
WInBr7qmjbwB8IbRYvYDCCCtDG3U/XQYPSpvlj4BC/oHaOoMLMEnr1IPo4oesL6Ary20GZThsivh
YXQwa1Dvzt9CjvczT02Eb0nD0MKIXUC4LPQjrTfb55nE0xz8joXOhklP8Ra4w8g2EyePzkZ1K8BM
76RRsEApEHxswAS8hx0/0OeT4RoyY0LrJfz6C6iTUbV4Wi7qYVTn5CtNREp5v3D6wUAqzQHDh9TE
2Oc3iw1kvhSLATxyblS+uqOIz1PiSjtrafnmNCy27eZM6/rStKrmUhQUL2VLT2qP5xh5FwzAt1ef
+Mq+zG+ks7nkC93pg/ODpDam+/aUbd611+iyyyetMYgmmSsTMBpOGOW47RbIqZ0XwKTpNo6WZDun
GcmN3tF6Txl723fMBWbvaiUYz5OpZomZgyfxyk/PYiaVYXAAfaXuK2LcxTbvKjItXF68PEHUGi4O
20fDxkeKCoOc3k8sf/Nn+0olBSFADfxR1oA2ecbDWK5vDRzvbl92Knv66xVt9D6uc1kFxYI2npvt
xVZ3+fQA+3HLjW8tBBqAdB81a05I1PLVCHqmk3tU5THTNYLyELrHyuxXjOCn7213pc55y5FOxyzB
aqRC9TrEtBUgT+WkZXayaRj4Cag4wn3DYWSnX8XHm+jH1Klru/83PWlvtsbJZil4oOW4/t2HF/Wl
9o1sN1s53HpNun7hXXbknyEvxhww5joBRqXfx7QjdI01KYACvP00IAplDYI0i6CCu9Y860pI8kji
VsuDy4kd9rO5q4tVzaOXnW4QV/dZhMMw1gN3O0mSlb9n6AiClxGn/gazOzo562lBVBZw0cMoeZtm
3w6hAuM14aQ91wf9NDbjFQ7XrGzCIb2JP0YKEjon/jiNF6eczoOGKSHq6tsLiecrpEJgyH0vh/vM
PBoGr/xNmRvx37PsMfQrPGWzq2HJxZpeW3TYrvuyvcwOgHMFf2iqRQIoLz0d77fyZJ1KmGGiOOk9
gcRIXxJ1X52lQGbGSeccbLJ692ho0Q57QeBeq4lVvoN4Z4ffqm3srNFwc4qVdIamHOH2hl5RGT0K
+cOnboXJGJxHGQntI6XXjGR6+ICnnJcOtzbwMjunVNjWD7hEDudxw9jXapLGALoHV6KlYawcPSBm
qy7t6/wveEl+k85K4DNimIOlFA8BVXtsY/bPklITA0OArLShe4xCfNkq8lBWixofDuPEUzC5oTgP
zBMc5og/63M2xHwFh/+aAi4xIYgjdQOCI7EtRFFAJjPaehQrwMHUlcMcoxBJBQ9a/SN/PtMBgRHI
7wOZ0WCzriek2wABLcZze3QRWSXT4YS682msMaUSQ61K+UFK16LnWCbfKY/R6cdcxL2euphpElua
UV0s0HSXQHJ5mRmoRZZeUBtt+mP8OinZg95CeYqpiYeuTGoxQldGNM4SGoDA3UowxcLGyL7ZTVD2
tFW5zmO/AEAy9VVJ7oqdvYeSv/NXmZCD5oNsNiElCcaywmAVxS7hFRs83otnc3nCzfFqlEIRYgFd
JXEaFKxI8fa54odhyeuDeCperXKtJ4prV1eqb0/tZQBiuci4S0RzwTj2bzzK7HyGTf2FWa/UBv5n
hPbSC23+T3VmvFF8cxMADakSNjpYVlG+jExcZiQqMFGEc4yqw6zgiMY1dMpnT0JKB0ulacLChiMs
Jz3Rn1whuvncWpREByRAwF4amlyTx58nncxKSnaFm/i7vuwyaevG+/OeniHKJmIzsStKbUQAU7Ry
fwkDHDTyWhKjrK0aMPbEyzyD0NXp6RhPm8UrGcTkiRRrgc2ds5DqMrjP1GcnWH4K64ifmvFljJJW
PJNgsNVSmVhElmcljgYeYb1AsTTwAH29umTZTKsZmNzcFC4KL1hTgL8Pi8idxPTiElyw2fjN1bZ1
4U9jvNeSt1CuVX/bJkgML/oCHPnW831Cuj8FsjTiFM2MOz5rdjG7E79sqrU2CZTqJPyRpGjWRJv3
O9WuvJWT/pyW08iXcF4gctqzorveNWh75ni/VVoFpMn7TG5bUpVaL5o8kJYtlOcb27A9Ag2Rq42x
TcTBHJTOpi5yo1vkQH+h83LaoJd0Ddzlov8LECSagSpvCqQ/kiS7Iu0xtKQJCgoPMqjUUISEVDmU
b1jCUu1gl22lT5V3nWT/syALWgwyn37Y/zzIwz8y7DxPeqSyE6f1vKd8RCnDdyBhreRqnWZyyW1p
dY4mGseteKh2bPgwN6z4dQMA4PguAm/WVuW3iyOXlkUmWLmn+8BFWODzztOS5fEabMtVtyivyHU3
dXLxleDL/MMsK9Wgse0mJtwfszjMmo2X2d8MEcNgFu9Q9Is+ouZV48JX3Ro5CcRHyr095TnOOTBO
ZKmUq3utO/Z6KyhpT7+7LRPiIx2UL99a+SbVQAp5YJnqcbfdt2m1nZK9C65hdqKpT6BVrk7JJpVO
ubWMeY8mham0Aht3msZ+3WglCojrzUH3CMKSgJHUaOzARORTujNAUHUXh/mQozVjfozi9dPlmUF+
6q0oZ0kE3+9i6O090WEgIdwkLjq5s84IRTWH9KVLgFPpKsWDMOcnl9MIsIVd9KCsdocUKhu1zPPq
n5o01qxO8eFKtob1IJgx4/YbBwrQlfE0yANQTZrApIaFfRa3ejbPImKEf0AKU3G0seZbJm61FKJq
NMgi42/fYNlUighF3agw8WfykoZSG6U6POWIsFgJxmM7gm5QPG522l93kRCNBt1GvTM/cihSXXip
VrNeFpxDnjOpe3yIn/0pMqIedQk5XkJCFViIEwMep9cXLlWaSwHmlyRR3p7/RaSr8TgKUa6w9shz
YgDPoSIws/0uj1SaEKkctS4+El95e54m34rMxzYenPyPbDTLX+m/nniR8X8wlsMWkiTOP5TzQJeN
J8qMhR3km2TmAmDGyld9tRrL3xzxZfZKsiolYhTxWvoQOW+aXoSD1U1HaoW5IfcLF3CqVhd0ccvi
biwg6si8W8HRAqiw7A9jffWvUNqGZ46/UGXcSXbcAPUNZYD+IzlfGPYA1UbqBNSFXgBDuMzqEr65
iuUVdcXOJNKMTH8VwsnKrAgJb5fn22noed1yi03RSW/Q+btbR7MOwwTu0G3MCa1NWZ1zInKhP8h3
MOs86WvJnAvnE0e6ISyNRSxtZEkZ+s4M+k+tsWJVCloeUceeySoF3zxpm3IiRQ3Iwcrmn3z/nShG
2USG+AEXPz4ntlvgbFxHKZEaqWPyfpZt4s6a1CcqABSq3iQNfegQcOf33S6QfFsGnhFB8gEWgTRs
ZXbHH/GBD8O6wz3FRqpMq2P+XoKwthJeViCk2nHeF+RgsPGOszJBIs+6Xebj1T+vbcap2lNKYL+l
nyMXKukKplaRHg5j0ycfdEVn4PnklP3oeF03+0Rg5MhrXh+lBI7l5ZgIY0oP3Kw+WHZK06tlcp9M
V+Jppo88kCREpq6JyWd5e7ynk7lFD0YcemfratGLAMEFtw6GuJaQ88G+AjcBGq7T3aB11ddK+j05
U5UDXG8aIxap8Dn2QAjCeCCEjNWiMJgwYWhnH3ROPiSvLv2rrGfnZs1D4sOnV1YvRjXRNyO/neIl
pZcTy+QkiML/oanN7y1Ha5LWBxPB28zYzu37QWQxwjw5CJBgXahF8SsEXxdHw2R5Dn9zHsyWnbkl
Fs5IxU4ZE0yEb2+VoNRph7RcB/ERP+KhUk+ADxfj6Fj70tnSBU8hFeiptD1O0XP83/n5U++mHVj/
cOa/4uYWKqCEQPr4ObPcP7oIdFs1Z6mhQaeAEbrdJxwtwU+BGFmSMF4TPH2QGIibvS37abFMYHBn
nq47CdNuALgmLWnHr1bbnVzSifLdi10KfTIgXtjHUtsc2CPV93YJj4zhpA/30kjHjgt7RX9svqM8
D5XTIssi1BJfmpeUD9gxFPrQhiBeFlwuKVA5zGRrn2ia7sczjqbBdkefLsDkCVQK9WHygAUdPdm3
ii24Svm2pFRyGXBHb1aBJykpmJhBXvAqLIurXj9pvj6heJCDIgtFjFG9nIvh37yK5e6/FNOMS/Dl
LdqhUDmzcvk3ZplDBVRZ6su/YL2YeKjCboP6RdmOlxrLR7JMbRgYiBfpzqRM1zd27ca47s9MR36U
fTnKYuHSb8xr+3Idn6CgraAIUIR5lILTLDqO3ahcS1RNoFRUx//LPuii1dF8DIIA8ccGXR/7L5gz
VulZR0QJqCPYlj4mRhAb1Gb5sLqpgYeUhlPAGO1QP49+Hr2mMOQV0ggYjL2oh9BNp87pg7g8Qfvg
8oL48ysPkBGu0+9z8HJGLrUz1QEG2HFNdSJfO+g/DGWRkxrsyeo6ZsmNEFU8BzbtySo6a/5wuPTI
W/mPwT3EToy/ByAZ4VWcC9h6YAABZMLss7BonnDPyrcy1HqoGJv2UWO5yMDGIS8MANdNdX852B99
dvDtkqEeWXbHBeUKixNoXHFPS6AvUDr48tkerO5yG2f+HlwAwqEKGJP3fD/MruSA72pYhyvqY7ZW
Jvi+QJKsUUWp0ARATtN5fVd6WA8GDskJBUWDG5Bl0UEh3r2J6XcWa0s/mNmMXgreNutWElg/iVvd
iSLgwYJBnS5Ani3QVDsuPB8bQRrjfRgP0VnLiZ6zuIyQW0k4b2NjjPV2SuFonEMuXjU2nOhO00Fn
cc+2ySdQD9vSCZQonPpvO+IseU4zVvRvR5A0ixss51luPulIOrTcft4Yb9lX7O5LncKc3CVnKa1U
5bBnDnSgU0Z+W62gGznQkd8ojjwTqIy5saQ9Q2hZgqeq+JclApupgIjcIA3u2hvsPXhcZzxmzPxq
RfGbNKvys4vGP9egxR3mDqV0g+m+rtOEPiYPktaQ6zt3hkdUbD3p4lG1lFnWg8kMF01Y1Q2+3zlp
n3tseK5YSSO8YX5wnIkM6g/TrPUVrSR3d1OVaMBa3yajbtOr8DisshWhjjauc3ztQXz+r5OnqIMZ
i3Wmdts4OAP+whHf5N57r4nmWZUVMUx6qKcynBBGB0oI5SYE6j4B+jF7w7PkMd+j+QSSYFgxfIh0
2Mq9c89IzWFuwSPqwpdFaOtpkVoYZDgxfy5UJ585Re2Ze6ZtIF44vvHs1Bfhhz75C15xDBcvJFsr
R5XTaqgAr52UJjLF4mF2FJB6xJPOPzOavqhXapS2TbrIVirzOecKfuUIKsioiXOXV4edY37mXOou
+PN/86kdIbRL4JNndDrpXMepMd2fkHBphstC6fM8m5aUtJAaWkzrlyKK5k3eFK1f6CJGxFI2XPMs
pHRfOmPknSTcaiNQEJXk3k7hEv1K9gRJBggpcQDmh2dJJTq7uoC/S7lH3V3KvhEbXcOdKaxPjlKa
TNKkje6pO4cNFVws92MCV8z+HjLCEl/Wkq0ckEIPT/1TwJ7m97x8RNzpeP73KcoXC6TwsOtDLy3q
BXwDlcvcFsbktnF5zzKt0NmdNeApzDLYnVRZPBodI1oxRNPZzZgAorbTC5CzCP6yjGh1A74c/OwY
y9TW88XIbwO2CAFEQVDpkJINUbT1kedzN1hi71dmMYUqUEb/hYgI4439WHchiKDqs9Ly6ds+lbkJ
9G6dzH3m1007q5m3413IwYsG10xFm9RzQSovKHUohfwoCvxkRK09FOQOA4kY3Lmf1IWA1Zfy/h5P
Dt7s8qE9nweaE52HPiPwd9n2P2pyXEGbSVUilbh17JrI46d9vjQi/JIBzHeGzlu+l8rR1CuIMfIy
C421g5TgzU/aJ0V6WI85SEw099D8vgpgPTD7WTct0TFz+qpuCf6jA/1Kq9tjgPbLAHXeAZzFhw7v
DpN2YzGOeUuThJ+qcTJ9dZcQwxP5pLsHVp/0h4aos6igYxNI72iRbLnGeYY2KLh3kwAmWKjj8el5
hxgDrLzGSeWt8FoR8zrgcTLH4/6aON+qNGekg6zTCHBgVhCJ+CKXXzkWPz4Hg1u5XlFnLePuJyNc
SCptE9gv/7y/Dk+PFZGAzwcv9okssAgnNhFoTmQYdBjHjjgIfyeQlaE029oRGKzChjOV3RPqyWBk
Wk7rmteglqhaab8GOR/t7ma/w7aI2UEf9LEbSTrYopLMT0tza+30/dOIfvPt8bjtJayopODjwvlr
VyewkRoKlnBJ7ad4xos4LHC18G97pRG2ZvQbFallN6UM2wOHN1TGeLlXHooffsw5TmPwDZFD7Qe8
97x4lwQnThN7uwsitTkTwLPx/IxtLH2icE6Ywi5XF/jvY+s7OZFdAhRWqCEh40gTmscg7ZNrwLop
xU0rGxL6Tf+PjgfdWEJNNJrAffeXfu23fo8OTokZ+7FnTbl6NApIadpSuOVOBCG0f3D74AX2kqL0
ffAAUcjsoAAknWLbjULD+Ti2j0c2c1exbCYBgoaJngc4ed0VQbhD74z8uFT6b0Onp5LYYGmm/EyP
JBViYnwMkCtARt2lei/WmO0jc7CiXm/MfO5CSOqQfBNELyTUciDm1RB6Z9+RQHd5T17Sh4InUMiP
qKbCV9jjwOZrJ4E7+HaNwK8zD7lukwZDd72ZdX68Unu5GIbo6SkPdxNAcXJwOlwnTQT7O91t94mk
lnfWW9svmoUs4J8/NMq6hM/4WqecNk8IsWKEl3gULroS5RbLnIXeb+pA6CLD4nmnZTORyr8Y9UrX
e+qhSYsO1lOotzVdOAT8ZZZn3HFt2YM5ryB0L+oI8iVVPOIlHL2QZtHwG80DaZm95baar03fqhR9
1gziX5wPoZWKtRiHHY+63IATsQ/AHFJeOMn8C3eBFXdD5XGIzrCbTGB3c37ErXHA7ld06xSRpD52
J8BdNlHFLTm5CLxIz+mLUTLLgqSNIpyAOH3YKuk6cVeCG7QC/cmNYj7U6XZE2JA+xHMAOT+179qk
9CvQnzHctVAK1duLl0YCLdqzJUt8CpNCjmilzkhxJhvws4HDJC5SRch26lDMUqh/VsAotEtnsLP4
DpRu/yhNh7CjXuprNpOor9vBhOIfEy0Dpymr+oRj0bKSNx/O1fzUswHXlHBM20EiiQiHcwzebeEG
TMgLGYDpRhZqFYNWPqhKHkt+H0DLR22clcRQUAhQs5anVx+UiEX3gOiAkFCJd/NZsQy/pLMKxDU8
V+ZnIId+e8tPgsK94mBbRpRyqONGcVdHFM7wExgU5Jr5ojCMN6cSe5H/haBzWMsIenGcT/CWXHzr
nad0lNJFsf7BK/ZOPAqY+8FV/ojJ8B+xcKlGFiJlVePlOC1fCOz6xMeLkfS51Odw69JAtTsM0W82
q/fVy9kYSiFPux9xtuozEd0J84gFkc5JlX/IU8dfiMNRcq4WMtHtz9To+F7K1b68FYfIvkX7WKMl
Ytct4/AvB/cO0ob/C+8LZRiSMrIdpguIEP87TwjPFCKRHJqvlKQ16qibuLUb1nZMt7WjlKPhLd/X
jjQljb5nkpFY3anh400k85iS4sW0tS3b6HpIHuVUp6gTO1jERXCuZyZy/CJl5+XoB+D9/uk5A14c
YbqQp2NZxpjRp9ATC2z+zXRv6lG2nYqMVOtAKClSygx3OuY79HaQ7E1BTL68SU8E4lPU+eo5PEHc
C8PhGmt3fXcUKyUdItKo48+nR2Mxz+c4fRN2xCA9bThcOVZipt+Hziq5KEsycqsuiUfT97nvpAFv
rxlmNYiJH8MFku1UsK0Y7HpflUrfRCuFE6Ia+H8XAXWSnAn+v8OZGY5qqy+HHePEhB43t7teW1ii
WY/WzdafexFHPLRia+LW+VWQpYDfzDdlfsD35t6hLQF8zRBWb/8P8T8kU8PMJfqAbPRuOQGcLCZG
yCw6oSe0NfWUJ6e/8WusW9HjA6KhUplyOdyGMfrdFO5vW2Qi9zGhXPztaRiD0DKHtSXiYdJFXI92
obutn0X59S3Q9jAiFhA/rj61z2+BEQvZ1qdzs7Y4dAD6S2J+Y9u2PCWapL6y3+M81PfvjxMxaYMo
JltJ2o1dy923/xnoepY3rqH1I7uxYCuAIJS/RygDuwbDbzAWbujL2He95CVL77CtL+KH76l4X0zq
HpVsOh8oHPJwPQn4hIbz0ZYvSXCOd7BQUaLPkfwdPzbp0uv0C7uhfhQNPJW2HWaRaQ5/Rp3wRc1E
Tyr4bLnzN9V0YW4PMOaieWmbbvAowYVM+10J8zJXV7pbJc+LvZpO/B7HkGXPd6XFm7L8rrodahGa
lZ1+aijFns8Y18A5VqfAVUSrNf/18pFiFPg9/fiMZp1qGHAIghbQQlx+IV/AeU41xBIqnsO2KSwP
JPio9wGmIK+rewMACiMcnxoMBOCFfxEABvjjZvfy0bRMXH+SLwLPIXHoUCEEhaqc/Tl8zsua9YCs
rzz1ZFRoJ09jJGXW6BnS3xR2rZnad7wei1NrVcqQrbm8e5avL4ARGHqYF7nB1u1Oe+0lP9tzuIdQ
NTmy5E6Eb3Xz1IMxKXZCrRbrzokmkMkptjgXohEoUhqerr2r8TpCLd4S0ry2goI6fKkMeDG1g2+6
CIX4sihxT9wI/a21bTVjXtH0m0p+KQ4GGC6MHSCok9eaCs8ya69xj5Mm15sYQXMB4v401fKpkrBj
npFtfMDzbT5fDa0gd+ZNYUy9AfBj7zWyc8mOaCPSPD3inCKU5p41QQXyIwk4DBDbYuq0h/X1oA3J
mRKpjNmzStMqud2xmNQw70gCK4qFVLGBdcavF703S5tMw2KEVfZyYJ6PC1f8MHg2K9kMmM29mHhW
/fl3iJvtH5noWqCIyxYjiCl1ttH51PNP+dPr6i2M8JnLhqCS6TEWFvA+Z0IpkmCKr8upApZ2KMlL
oVW7v14v+X3AcJFEIPKZuUwprrKURmvKgUe8dMAMsvWQ/YKfJ71xq1PcwTl+dIKF6jGZG1EfvLfH
k6hoAOO4A5Ige3FQMAtgrH2yL38LCN+GlNGaUtO7BTZ1bb7P07odD97Hi77IelZ/HpsdLikPPi5E
3qFH4fP01/MVTNbamovDk/vQ0AGfQOHeCgKnGMpaNt9xKpxFs6m3fgTZXk+HzbUGFvF0Xc4bOBYn
TkDHetQJvoSZpImL+hJvyUfB+e3QakK2jHocwGO24a4jAkyZMdO9TSAUKWMEaaDhEn9UqudHIrZe
81j9a6bKKFcigkc4fZKL8P9Nsup1xKtGBmII86nko6GEayNFcZiN2kOHGOwPu4+ZYzIEO24fWF3W
PF8brBA7PvDDEODs0mnWIjF1hqrrpPmqgUQRCJ2tUoxFFyd5xRWooowqiaq7UwMfrkvaPk+xUj/C
vkoRWwKLVOukKJ73kg3UBMs/YZiNyGZReqixetWTILQHckMwVuKkL+0ysp8HkRTh3WiX4pVgtAhz
j/B/z1R7eizaNqOxT6GhG9njyqYHJhUGVKGpeiAsA8CdYi3br2VhpRtYbJCFd7IkMfnuLHnuREWA
1w5QZOGp6yjh9jc7aeR/hqGBT2SF9tUAs+KJ+7T3m5iY2kOf7EQgEmPfltuBgGiv4TahZdz5Bs0H
Tqc1ZBFGmxcUmiUirfksAUkSJqMCyXvrBuBPQpw8xe1YQLC9QOq4OTsKX8DRMf58AYzfuslPJlaT
1uIudRvxBFj70K1RHC1HhHnYJEi5Uhy0H0ssA1CiJs+aAWAed6oVi2cxilb2u5L6gblYufPRzJLh
iKCDzk0UaglQc0fsMMRRk9AmBHk1UKzUEs1U0YXL/5m3+0zBZNCredU2lHLBe4mjseOFjcHIzcT2
U5i9vDu9V4eRRPEwcvne/Qc3wz9eVgGEwQkdF+NKyYWYJJ8indFeNuCC23uAUUTGxUiCxSSwOalp
LAicP0tzRS9ruirdsXoBsZoS9l9IOh98kG174rtxaSuo+X723YlwqwbXjaS9Ov3Ret3BWg6mTcff
cW+i9Xi6DpbyhLWHiK5g0TrV7FLXnKB7M0iRktz6mRItHVETJ4/0l3LbOc744EMEp9HytYqHBVSo
CKdE2uPaTmhGsKikxep7YZXArwUu2KrU9AheY06akW983rB86mfzFb9l03MKR8Xb7hrl5N5pOV42
tEU9NWxv8iMROVYaCvPxQTSHZ+toiaS2jJapRkrloTIhw9kp9z6K5IpYSafK3/qSb3qrt0cLeL4R
UUBlaBCZZWW3rH6SGyxtlEux4VLM0RkHOxOG8q4J0wBxl54kdOCcRGUK1WEEONFzFeTk/TsWUxyl
7JVh7f2X2PAwqkPSusLc68hTHP6e5kkbcV1Z2af665upzxq2dMDkXJWlV08aLOAfylvr8ayX8ovR
8a6tIxIyycZZ0Jd/dPCR9AdcDXH/3lD7keKqwVcCPdQpK9A/Jt3rIOLkIfO2/hCUO8VLFcNI4pMI
ML221vtwci7apL83mChmFLUjooqS7oBUYcKfq2VReNW/lASZLxqhMCofrOIlT8JJBq18jg6VgTNk
LxbsFhOPPcHAjDF5AFwArxxz3zV9AEKbBhWI1PnXh7Y63Ni+o0PkAO2bQKNdRjEUbI98iw7QhOnF
r7hJYRJHXTtd4x/zh/wiYGRtp3HtXlhfTkjPgFTp2/B7l/AR/WqgYxhPh4RNAf7wjY65oPgPIy8T
ut/bC1xQtXug12Mm822PZx0CQ4kixmrbqvbZ6yMaIZEaSyuUhQrDMALf2zmel1yMxkn0Ey/+0DOR
lpWqrQ/U0U2iflYXi+8pd6SpKEf/nbxt+EnM7hQhLqcJuX96qe2AK6qQ6k7yVhbWFQiq8qXF1+f/
JuquM9/zzHRvHQBNL5XAgGU6DkihZrRGZ3arr+rLpqj+MpjkrxhgpzjU3v5m8bZkbycXdek31afu
BhPdSIXwEcaJQs5sFFfjhYsJnIpL0EbabIqy8WW37kBdG5sJMrWH4t6v9fCVTxyi5bTERC66ADAU
i6XSHsglfLfVaWNIyRDy80Epl2/1Q/qSoeHDfTadIxzUw05jkLDz8TdtnvcMzPiVT/rY8d7W2Mxt
duVCcNP9zsk5y53UdMURWAT1rjPDfOGBalkjGj7S9JKIOjKslzLZh2X98oCW1B9bp1rjAM59ykLT
jfdfzwGbQY66UVuLI88AwlSKkpS3qUTMA2WkuJXUcQqgorEWbc+T7icnE05VW+SLmdzoGbWQ5Gil
QFXodMYdxTIVoMh8HuIo38jV3NJ0tt1P2zysAZMfkLfaLasAPiQ8AddD4RulVcdp9DJWd5rZyO06
l181T3FhWoDdK26e5zDfRr+XF60fqh1AjZbS3c/Fj0pelZSHwTP+uKoPyIQ3n1kP4Gh5VlLSuVb+
oEHx+7GtdQFx8fPsDVikR/NTZHNEwzNmK7Kuc0Exyp/9ZiTh4Fx4etX5Rl3hu4eJDDTGUpBbGjtY
F+/4ixMBJoEOrHpT94NzCXX9KEsVljstaTEPoDxtmfQJZsMvtRd2kq80+qdjfT6MvR06nqufiyAJ
Fneou8uYsZWMmjhW3UxdC6t5zBJl5WmCQP2UdmzmeuNJM/DlwtwrGh9xoaCbtZT3HahVfMjQSJ0o
eWFfnGEVGNPYBC5ptaOMGYhHgPNzLdS2Yvo+exMXCnyMg711se7nY9Z5ZL3fUt5uD8iS5Ga4fROk
Y186JktiCE/yaPQOawnSbEFE/3jSiFSZcPc4VNk3nePLGhAtRz9OVOTL4pr/YO8DNRDscps93Cru
RKPYsFeA5QiU/Fr3P9jkijD727uvi2ajCC4Auan/HqkUJEdYdmdNBnhPnUszIQZyTEQtwebrCkDG
MKNpxoH8DrBOD0UHqLZy7RjvuQSSX7B+NS1vZOzzOs8QxsjMMeD8gyWDZNM20yNOTagVuA9mayKf
xwAndwZYRVNBndNBK4KQCq0wDgDPszgvnN5A6+yZe2otiByy6dSsVxjdDtp/LLVMUqOxZLRUjJg0
gyFb8Gcn6NGEjcH995kNKELE3BiwJ5shooLfriM1en2TUuVabayK91KuQbzbWAbTYMjcdukMHiqD
SRmKsRosYsjpeqh/OKUhBLuIh2axcWDQ6UqF7pJylT4VYdMONhYrHlmdbvkULLTJ7FZPihoO5ux/
qWpRI0/sP3mas7x12B6vpIJqm7xM2YMXJAASVWvnH8tpH927PqVoizxOYpCNLaze7nN8oxDqYlus
3H42vkO39uGdpOEsEM1idXNLeiOO+SBgGSPyRD7Dwue3LPf6jyBPdy0ghZFrPDy7rbvzJQPb8wwS
1niFJt+C1chKBe1qK9FKaVUNrByY8/n5LmNkUlxY57hNyVkHtuAh84oAqgYM/L9KBkCWDzh6yS78
ZslNJABHcH+mq4HBULcxGscx2bWNlC/ONV030gdlQ8tUyi0zh3bnofkL9vsQd/0g3YMOaza0niYR
CifA2g0sXSTcRKej/epfstRCtRJLzlRj7wNLMjIr0s4/1dJZn3B27OTqxMLfYSwhrYKxpBrreZHp
u7QnYbobyX75ZhGLm5gLVQb0IS8tEiIhUfBpW/2Q+wln39gEf/Ssb/4nWtLpwuh9B5bJH71KCC/y
5M4f0R6Wvykmwqc9Oim2Yq1ho046zi5PtCovVYcWycHFywmpDND4LrspY2GxQ8Qn7GObP+E5DpzA
4ueeSt2T9mqtrQcDA39PCyoIZZBOOeBbflHPhbAAGqMCZY+UecmjAe0VanQZqGQqK3PaC2qSrxtt
6+CM9qam/kikdRi1k/sHIdu6FyHUcqFkdnMYWy24oqZIq9f8sNXweH93TixSQWNU9owlWUKKzV2V
H65T5mg3AWVVDQBf6XhEdMfCOMfUU3Qp3VsgqGsfLmu9J7wJAbbXMl6YXVhz6B0TzeHHt0Mr78E6
l9fHaaCIAzkUdLXw9qSArF6c6xp507/JIMZdanvIQ4La/Umb7gImR89tWJRtjGQWMYQZiWnX26CB
RWxKLGEIZKg/8h8C85j/s/SFBJOGew+zqcz6htlUhxvV1gdRwIfvHh7ub4mnxTgtJKSi6BwR02aJ
L0MoskEU00wgn+tjy+i78K8tcZBBahrnfJByVYkbd4Q6u3ZgsgBt/MCGGtNyzI5MQailjRkXpJoU
B+YS9T7zOBeG4U/PrpyxAe4jURzx78fwr5ZU0EyVcUZ3pHJLiyIxzAvOrMl0dp9zIt0Jv2Jdy//l
Ong1evh6+WvuQp6XfW9fxQT0f95yo6DQzXELwOQzSEp+ldXgx81slUWpmsu+j9AUQlnA7iT2Ww8M
MetDYkRL2yGG902LCggyoEDbopN7MD5W6P4nQcmSaJxjOIPIopTO69cLzMmnMqaDdnzuAYgwwy0+
/cQfDryU8EEtOFbhJ3AA5AytYsjrIAoq6Fh8DeldvO8MkVrnlY4xDF+7vjdYS2xYZ5KdqPtv4NU1
MFoQH880Qj4ulavf0tFMhnTnj0mAk3RM2C+IVBFaJThUkyM3p3nXZxWfHaEavBLdTHZ1krqmbJNM
Ml1Fs88XKA1ES0HDLvTfgV4ZUOyDxCTZMGcJGbkQG++MZH5rekfSD0olb0ARMqumyNcmioiWTND6
7xBQ1vshvFscSKpb7JYUOB6UbFkfDYeKwru1KPqT145aMYP0iKukO0A9OgHEbKFnzXV8mdgLovi8
FMxx0vcevOLTzyjXRieCgEzLqcBYO4zjmqAsjAT5m2I3toU/33BAQ9ihx15FYFnSLyMNznXv7WGS
ZdSMHpBHVZThUx3eKp6EbLXEV+1wiidV3vSgLvLpXvWeSIwnFGHl+KPoReJDxo6HUUZDch1DCexp
9T4UQ2928mzQ4IQp9hdp5swwcZdodVvZIqR5tHcTVcCEIIbiU7p6lAMQp1CkVUfSeVVLNJWRQJLR
lH38Teh7jPhCBGzR8K3wmlPl+7l80WWjMWbWjjL3Ii566Rm0PLJk8/ZT4N87Ax1Z6FcUSbg1LGW1
WEY56klzXj1XnDwp0qBco0p1iDXjb3IThjocts6MosbpUk2efuQbzFeQqNGAkXsszSFkEtg0HTlP
vxAw33/iUyYBIc+Yu9PlCeek++LmHUzENhTHX0e7KGWTCBC0kxeFITWn5MGDVakhKqLDvEgPjHLq
LOvhye9/IGHziiCqqRqtnL9uxOI/3R8fSXU6N1gegpcQajnzy5MatknPqiBlBArXRqcy1zI2NgF0
KH4TU5SjaDODsi4pWwGdTyAfp+n8wlqhYmRDJbPzeh3eGZnsYgTy3nNOawKdfLSKT2mKvEeku889
5+wumbnC2It6lLViOh0rlm2PRsSUWe8McZ1F0kra9mSEZm2aORlt+Uze2AnARIFLcKIFq/xRs/xK
bIXHC0rhk4r+0mN3oeBbou/JnNq2Mzjmkb13QqBeZZuyENrWZtOftJDJM/AhG3gw88WkIejvdsBz
0Qclk3ov3Z6PAG7ZG5r2178GmZeLwI+rjHKH5raZYNpINmyMEqrEuKlYEF1h5Fkd0/Y+dmNps/Q7
JuCPdvQLyPgrvje3K+f01k6IKar2y/CUX0socBx5VmzHjm4F1XPtzzWrmhXdI/BfZEYpd1HFmris
V5dIJPI5v62SKw59z7YMO2irjsvcPIgLFlocWi0bx5WPlkHbT4ZKSAz5I0Zy4oEoZ7MpajV+GmK7
yelIXEJuBB1Me5AwH72Yt5TynP6LZW5fWb/u9HiFrvhOYxk1bJDnHAxskTt8yfU7eG0L4RTH+9Pz
tUFMmfZoXpn8SCyfiUIvEgw//V4Kr4BJ4AQZd4rpaSsN/A38wsqoxFM35Jevwy25m/FdIWhXh9GI
WjYqEjVa3miuFrznEc2ZsJ9ruLwG+hA5SYTmP6UtU17a6IpmDoDBLprxHid3fSOIxR7W7kZSoxKj
MeNmEyFBeCK7k4UdAbuYS8kgBwKq6DEStmEbnetwhDRDJnn+CuWdVaICvvmLdHlTqhuRxancO/Wn
W/DyCMzBvtaI5IlskDqDoHLJqNtO9VXLaLH/Q8gO8zYxgRjwD5Z1mcJfmCv49Hpp7/7scihQguUc
CQK3RKjKAJ3GRCF6f+kagTqtqEY/z9JUCKjf7GGd9KV44qBBG6SQRtEVGVqMzRS6VG50N/G8nw7+
FMRksbw+I8/1iPePQtRIiKVZJ7ru9SF5Gkjl77+raHQsvrHBMX4NXkHJYoqDvzQegbFrSakdaD+4
9YScV2LuweYGI4zVVj2m5e/3LdfR3nhWiSAWn8IcvMyVwhVFtElPy63B4DqlA+mFxN2L9XIc6EXh
wIWm3Ht4jDlPxYMQ3CXVVmBHZcHkGBLHQOb/09sEyOJbMauIBjRudrTVFvEignDQNrHZjo6W5x7p
NKvOaZjtPqWwxiFxigLp7rQJqvvl1xEF/zsoB9D9oGgBLgeMw7AMqW24ztDNi8Ye32T7SuioEgM4
xkM8RG0RkB8a8ye47KpGNAnzStFOdYGBkfIclDZxazxaLjecSU7219aq8SZWx9pa+C6pmJR9qZnQ
HvxqfGq3ZFLfReYwzrWQ/dTxXs/dtK6851eypmAjKzvV+9mzIKqYUjcWBdHpgb3KT8ujFRvx85kg
hv5QO3cnCkSmmLaTYxEv1Y0pykZU+oK9L3o3oyk+C77pYC066eQLhaiGEYXcpREGVrg6U6vbIj3J
e05+jeHLBzmKpdkvgnaMR+/IItLOgKjzWSnnPEiDuDfiMBBvUqqoPOOZeIBar0zSE3XncYx5yIAz
vys2dqXGIHEH1An9OtfKwuCSPv9C0bfdRouhzoa26b0lESCiquRE9hZrx3MoNqWfZZKgRXJA+sNR
m0b5R0JTfp1AA5WkhFbDag7Sjn1QYzOCCfQFdM3E3O9OHnTWS5Pu5FBVYT32NZDYZ9O/c9pxYmKq
LbgnKCbTi0o354r1rRfpdxyGNq/gZ45oXfuKnNEDDU3+3dK8iy9OSI/GfZQyNiW8gth05Z95TSdn
u+n6nR2wWGRDyBP4oZEGz4uRWJmtAWCseWhd1wfh8SHEkgPrUDbrtaFcTsHZsPBM2lITl8L1iVuy
SXXRw0Sq6IkerbrbBai/p1sIMmelW7KciSxHW1HralB7Efdus1hXx+GDFFkLCH+7Pudt+7yS3eZE
eQ3sj53pEQzpk7281sKqGZC+IAGovVqBclX0qfQw38WKQQmGqYzL2yjAX9JqgDHc5J6FwtlRo8jg
wScOM8jPeJexQVzRZYwWWaDswUXiOIwbe1SUhLoVM/PgwuuZba7ssx1JJVgNCZRa1/wsIek20XZa
64W/5u3PXjAc6hVhHWsOoXVBwyBz3dNq9/EiJkgWRAEkGoIslZzic3bJWjraVOWmMgC1lw4ol3i/
CzYaIycThnsmRxqS5j9o25JydW+WI4zUVy2Up3WlsomlQ4HwAznhmx7Q40pGrZ8g6XBUBquyjaF0
ELJMb1ag0SvIgyGBaTGVXOuwnC32ZJEEFD4A4H3rzTyWyBcbWTTIhBDRqchg+hPUs0N/j9EnNezM
cYKMgHNdmZ8d4JdV3SDr4Zq+QwhDmalqyctufkonBrbN9KAnsy02olLZZXgdmbNtH7CNknAvIj7R
4gkoojXmw4g0iiSw2Bj02cWz++X0IdwEkCvLEJqLpVc8PYtdl1WIGBRYj3xEmCuJF9Y0m0POpMzM
k3N/RXkBRBR6FsBb0N4IrNQihvFtXBLEDcUZTqxfo06JONGB+O+cWMHJJttHORHBY73Be1l0Nbs0
luEjGo1SmfXMsux7eOsCAh/r6Cpk/N5O0ZAyO6s3ON8Wge3cLlO4d4JD77Aiv/Urwx4AbE1DBvlI
0PmNQ1/zTLiNaq/aN2NrY7srDAr4+CCGwu7yhQw0Sii2t+yBDNNsXZF4INCNTPvPSfs/Pi4Sve2N
AV711wB1YY9PLUMyxFo74RAvu6jR3DSxBTB7ba9CVZhL2cWuce2z0im/SrMnVbee41eNObmkE/sb
DhsIxsdcXj4TUP1hKWpdNWl3ZLAjoU0X5uJ0OPTCcWjsrmmmdhkD45KaathWHYwlndKVdoMlNW0t
ekXazLoIeAjy6v86hxPr7SO1aZKRl2KRvGXF5WhoIKXO0YR3j2lRKyzF9g04gJuXUPniWbzpx3a6
xGPMm54IDADYEwqTv+hPmbBqGRma2ClRZCyZb8z44izWe6ufUJftYq13ZWGj0xQT9pfsZWEzE9vX
xfpyHfgCLsK2pkrvg8ksBw7Cu/cijoIf+dbI8awV4JY7SKhnuy/FGFj3Vf8a9VzUPJTbPxQJ/iHX
COaWfb5ch51HfI2pSQuRWkHh6e/B6CEUJY6FSlYkUNeDonVIX4AvOc2AXhXCYD9IQW8JeU/D4n8E
r1XplN9rmgepEBwJM36MXi1WTn7nfCiWdwY87zEq3E18JUcdPSjyzW7sePTfDRDwXXiRwhTkXFJ2
zVW1/JDBwi9BM9QUb65jS5uw7mS6PVgh5BjWsrpvjirbCXCkRNTf5aZh5M1Ms8ySTKKbq7Y95H/d
fvq+mVf+aaEmEXEfgsktGCZcp1ZTd8/dUkwZj4TjaMhckdh7OI9zcgewfWnVssqk5IXBz3FF4RHe
H8EKmGe61eJepDqR2DuCOCRpF+mamBfc/DP/gW/3xofmRGVASnKO9HfPMu4JCOKazlGlnA6WizdA
nIlsK7jwDCU9a8l9dkXkUipoZ9QWpFj33gqlmRdjuEcTHvMxNOJro/MaJYtLA0j5jA1Ggf1m1QK1
9ndj14jKx8UyNpkPAWIPA7b12OFWdcKgat+O5uHvBaKGxNxDs1BKxg1ozyZhv0ZzMwCRWadiMwmC
eLHgxBuz6jdQ1d9yuKmcRLrBtf4iL2F3m5VKnRzoMPYEWPCelW72oHFotyUNlQI3YrD7nALkfRxS
M52rY+e94GQqwMfq7jtm40dDmeznOm/Yll1hEQwU/GK3Qi1TpZaqReH175rvS3wOvoY1r7gT6eQS
w5OVCAhBSvusLcK/4Cce+o3LxGYnLoEWP0TIjNx6b/Fir5IyoaMQdLYpdWtmATLOVxLVVMgAtig7
6FcAdg6a1cF+y/j8HHVc1tmPJQ9qPfHkQF9Hfu++I1bXtRcypvJysaNvaxgGQ1hp4KEVVsXEypMR
fMzeI//YjruF8OZRiaRIqNo6k1VNaVjcGVLG79YN5J/xjZPcbPq/Pp3Vh0RKTGGICAq+VzD6Zdi0
lGZr2SF1nFgZ0ojaCRIACiC8N1UZaSZuXVJ15RWbNYrf8fDwIIkBh7Z4YzMRDkLr66uSuS4TblhV
pyJzFGrJisxwcusHLUEdChSLHi9B4u0Z4AbhUYNFrIEJqUo4ni0orTy19mKMhXd6z7zq8LZXB+Kp
oXOHYwoa8022W9fQsl+k0TMwmpPeOam6tITa11VLFQQBRD0xW2+GrBYN24/EfLPaaXhYSE7zIZaR
ypRZm5eAtQVh/uvgESpQc4c0DiaOD30y4bzKoZzvDbpg8t9XG/3OiHANMCwmd+iBOhWreVUJ+nWI
I8orZgTqVRTCf4Ys+TXdOwYi6N5n0QKI9OgRm0ZXXy0xvOMXhwqYWNvpP1UXEgai3DWK2w7hQiq3
0XDVltX65eBWnYY9G2mbFMsRNO+yG3a7kD0qE+aML92WgoDe+M+OhECBJFdp/kxuCfnlfvV063A6
cY2wWrOnwa6ze7VSwozP9ILUi4ArltD6amtR9qC9o7An1k+C2rSnrIKYIN6nC90yf26lWEl9w2ki
7PZbn0UmhG7sYwYSyjCsiaG+17qaHbL6JKQTfizcDw2p9LNNVtOAHj6eiisK9kNnrGlftwEOg/0Z
TySobLlDb995MrQlkB24omnIwmvljf3z+/jg7NR0hDnKISWt0rCrzbM5fFo1bsU0B+GEJanRO5BT
mUOEHPwLA1Wmt2WOf3+7ZIJS5izyTUQgukX1ygNkvBAY0MBd8sn/00yfVukYwwha4arbZPaOUXRw
tnXS4mLOM2L9fcobC6sMB5r5oAedVuwqVg6+dNX6PUvJiRY405dzH81o4vD/zF3je9gBiHyNEM5s
ykEv39sNAq4L/iYSwPFXZ6SyC7/qfuDBrHkg+ipeODt3BTVbFvON0Clil9ynARAT9bYnyC8oSLbt
SlN6Wo8Wu95qK/Yd1UUs7KFx3yaA8Ai7lJt8UQXQAN2r6VeW5ueh82PhISpSBv4f18mDBxtIx01D
zSJ0TbCYNGLuG8GhlsjhBmzpgYN8V7Eiska2tttpNgjbbF1aQCACRnO4c81RoXZPoS6ZFKcpgJ+o
1ySiySCqdU7Ee8SoWN8MP8FQPyFxMVbiwkg1Hu6LTk+QiDu4WIhd093tmPGzF4oEY2xnSFRkpQo2
mfLTSmZComapX3Ii016a8GwV6BOccBCZYyL2n3NvYxRw7pYtcSo51OtGTmC/B1WQykTQoh1f0+hK
Ie0wSrJXD2VzENCarKxZZ90lfbVwQ8hg10PX8R1ARHhkzgPV/Hx3GFYmkl9FRWUSw0/qkJet4q/b
ov7tj2FLZEFsxp3zCeWJkFWAGIOUlx4AFwEWNA/XfWQbXHoz64RWRhTOiAgDV+sSWplXmr8MCvnF
IGs3DZYgxagkueSAq8QDHu7GOQh8nfvQye7NNqKdiyEYo8Xa6haATmnhyRMI3YGbQ2Y1xdmqpjw3
qP8c9hFaGGia4fILgdrnuMhaYxZ4+kd8tniM8FIvb8tHHX444GTknWBtcsRdRnllZGbBNeqZC6qj
5Q3XxYehXWTOeTJJEPiub8LK7WPot1YnFiIVnA3YxrFyjnR4lCMcoMlUQA6AMlQv4BQijMTqoTNb
b04LDXnjbacqPcVV6H+Ze0Sw8lwFricxQZD8yFP1Q3Qw73cfZN8kgn+qz1CdZuSXkpzXGOHmjFtB
ZFqrVntOX0qt+VIfHwhhkcK2bjnaGG0LekrJ5GLDjBak+EqZTN3hDeVtL+yrRi6XXjB/rc4wI7kB
4iH/DkDe7875CC2xjUN03PNfpWIRH9f3EcWjJRK3MG7fjEIyFD2sG4rzVo0/L4QrBJgjhfkYNIUf
0Q8lkxqIOJtReHtFT0VHRwZuEActPDLDbNVskMI1qtBznuEBEPfTSqdmwWRps/ZPt6EwVT9ccqgF
OfOw/vMPceJoI/MUdI/csuSKpXlzZtUNrcAV8+KkwptjatfxFJON/oT3EBQKPvTkYSBO25Pp8qa0
Z6aN8NGPuSDPwQb++1MgOI5+cwC/a5P5KrkcvkZc768nnJKUZJU2I6bPGP7Eks7RR0+VS24pZkU3
7w8Wt+cHw/LbHIdO5ogq3mxlOIVbhGz3rCgY8F6VlMMmK2KWlldImq8gnW+4cQ775zfWkQxcooQX
x6zx5evxFs8m1Egs3f10mg8bjs17VfVdHHhkihETsrLS0nvG2LSQdCSeOFBiEHIIx5cAXIA4HGOw
P4Kz7e45tTfGQJrMEmUEJ/jEkFbcI6Bq60FB52KZmoICy2H57JJiZbPtD7J2b7iE39m4qTcTf/jC
MfBfCJzX+NWoinyX0MI39cs7mfwhuaPY8miIsmVzPqihhD3rdqjVk425uRYT4wSfYYOoxHbDB6+K
nAkwItT0//ofom6MTo3Oz8unMEzuGqmz41XIujUM0yFB1kRvRSXh5B8C62iAr+or8muacSbvtvEY
uLMGzYeh09u9g6MIvCwRhhyLqiSlbcNCSzXoZCYA6LURKtWbIfBS/seEKPmosx1LCsnu+YCLlDa6
PjvaaC7ycFryF4UFrvf+NHfijxl7ulKH7XWLnm2bPboo1DJPwrEFhrm3zvgXmT/QtzSpLdy9VFKg
/DtHJQCe5ujmGSFXqnvvC/UFhc1CE5aPfmMB/SKsv6ecHkIo4fzVZPh0kKkZRPNlATYA4UYzuAxF
cDQ+KfZLFPcFzpackt5tQmwzdLpC1ZIbp94oN1ZM4gRVQNt6puSWPrZbIUFX9WtBN1JKwtQnKlB8
ivr9GhiqfrJdyO9mRa3e0uvTSb7OjJGYZ1S2Vh75sHVd+M+KlZIi5Y5XVXLXvHXXMS2MMHHmKkXH
QeaMHpSevRt2mTbXrdV7oJMyzYfPk/dYbIx92Zw/U2twKoj808RYsuj4U4b79X3o+bONSsK0LbVA
85iQmTZNFPG8vO/JiXgo9DzhlxdRKlYmWwZlDWHYR1ifpkKh/gySbpoSA41ZB/C8K0b4dEWeaOuH
PZJH6NxuSKJqWo/y+gKIqO3lpImyKUgKd05qWIvcEfAAbNTsSO+PoI0DfpwoBPjlyFtIY+l668UD
QMjro6LRPw2qKzbEa5mcRufo4Hp3ouV6rSytJoTZJpEdlxPM1pr79c75uaQ5KaxcCf2m6ZdJvGkt
M1sn1klT2xpc3BF5PdHqU0awSJQArEKDfHLE6mBUIKzb7GGPyBeqHBA5GdoqENZ2rzDgV7yTPNup
VzaAe09zWQpmWKG/t/HAH01FLU0BSvysxMEwhtJHSDCl/w3Kaz+8bTwVdK1EjY3spyHYweawBZL8
gUdaJHGQ7KRIuWdfZVr039Ihb2XULq4vqwvP5BjZPgKrnr+vp5hEUgczKM8xxgyBFE+B1MYN2tpO
N70zdYLeso5mxmG9jYQw4Rl1gHcjbUjdL9G55HtiutbsLbLifBMiuwwhjaKyoNgel9L6EDtDgIf+
JFEWZwufq5T/Co9rvmy+Tf/PdlAStZusBe6wbYY6MrY7pD3FXzEO9nksMBNi/xPrkfVNRFSC3vzG
u6wxRLKnwpXxLgMs5DwDZHkmWhY31sEzGr4Pn0mv0TYC74kjHAYM9BniOrTI5S9TpZ68fZuDmy7K
HiCmD+T1m0PRAiDHA26yy9MWR5tYvxUfelp1Bu2inCMaULnsmlyJPHxWGxTPQCY77NxBJiZh5Tl1
l3suIyrQ5o2z516mWpYxeIQ8FP/XpHqaTMQJzOHzEaoGJ3pbrzcNXHF5Povo+Cdy9UEnwPz6WfHg
1MkMqLFbQrt5FoMpGRuTSVxF5+Mk0CVywCwm5B9sLMcXNIYwL09jL87HWV08rbnMJ7vhAe75XArn
RvYPXILXNOoWsXRyvTsvBJ4c15aPNVeUj7k9DJewwF8VaQVZLYJ1xvAxjkXRmHOnJ8zKERPOvpnP
7WxgVMFTFtcjGBqMeIdE7TXfpHqwo7+vfC7iOHxqNwvA0/8wBDlgNdLog1yHkU5S+3MzvAqNUJb1
zMs1BYEyN3sIvI7p4HQCmnLDGU6WTZuyxK7AUVPjdbrNvhNVPjjPu1CmT5hKS/201IXELz9CQER2
jnjdH2iJ1mhbqnLSAxKiSGnirZsNScjed+WkQk8eoPujIvUqAowL8BDavGKSmX67wbciKTZeoiDr
EG7HWmMTQhrrm4CvCWJuSA3pELKeeVkrUSUWaJaiPitzvrMaU0lMw0I2X35KJMbq91H7Vq9orKm/
+ACXdWAWZ+wyu9mJeDZ0DiTbXytIXEE5mhkd/GN/EEJZemXkDCL+3LP28glid/U7NUpcptqmhXFv
9EnIeuSQXsytyQ6kfSIAT5FvdWTCVsc6k92sva5lJrR9jeIUAQaRE2wxJK0Rwa6BZ74sFXmp2OME
yQEqRjwurl8i8n94jmULk9wFf/PP2CQyQ3/lkCHRsa0xgu3Mc64Bgjwkx/zyy/WvpOuzuoAOyjJq
ie4mWaHyitwIagnMASHvqFyE2vIHwVAWg6qqIA126hz9QCPWbI1igul91XSypii6tBlF4OIyB8Pf
bogKVhfkCeVn4NZnlg7fhR6MRPmU36QbWProt0ew8T5ZOQrSd+G+s5yh8w6zr3Syzw2k0msTE3oY
/4wMsIBT4JL7dTBezfyJkDSOpQ3907CNDamPr1On63D6V3aJhC3rO91IyAdSEuECVnbVvQEtFm0W
oiySulu1POawdSj8TpzVFrwXcPF547hdh6z95SWDQkHD1hEQ5VUGa4i8P9CT5+XaFNU+qdHgotVY
xyXC6sVe42sIs+w8ooNGXNkSKfTfnQhNZHn0cxLz5XjjglHQBtG3O4vDwbbe4+3LSYx+9jf8x3QP
oEnYHtcFZ2bt/6ddwVK05wS41SAYxRCUoeI9ciiyr92/3TGR7sAKxqE4fyHaM7Pm4J6SULYOoO+f
WI4iQO93vj++reSPXc8pk/0qH7Y5sUBbh6eO0pUeKQeDqffP5pLMu+CCweiNs4AEED5ZSchA3Vlu
G8trC6yVK7YU03R767pswN7CzUM+Z+5VNK9E1QG37r38CnZhRKAtDDJvu1tWItZWXQbNeVLzAMf6
2zHReCqwRHVv149RIwi3/w96EGX9+AWU0Oxf/ss2B+rDgTeLY8o5WBG9pX61uIs39n+VjQRRD0A2
YXNHGI6/lhpu4xfMjroSMo9E8phAQba/PI7tTTsqmGJG7PW+Z9zmPg+rU3yePYcrNP9dw7+tocHN
0CCBIaq85g9Ul/McW/1TIs7uMLc79R4IEGYsELlH0/9vswxzZ1EVy/iZfkU9ZNdGwNSApC6RIAZX
gt6tYQTdSa0ZieuQcoP4gM8IaRvfe1/+/nvrOKN3AUmGxPIrU3yXoQkf52FGRUin6tQ21g0E/Y+w
DsMzNtb6BnlDyfdOSz3HYC4ofNe8zkamP0AmmuszdLniATa2HxioDHwuef59E/oEcAHe/tCxHOBN
O/oL8KUg/C6tuFoqYUOgVVusGOSQ3Ik5FWchYcWZ1Z9z0bi1krNNGuF+64OSA/G4XC6/06rxEbnF
+gjJks98T0Dl910ldLimSgLWqdmTDmPSf9Wxao7pNXecOo0wAhrQ1HhsW7Ilka/NDbwGPX6EUFT4
Ufv/CQtSz1T3ud92qgGKb6JECLYmMO3kRXh8XV6QNcb+vsp3wwSe5hXHAUiMf8F609zg8d4TnSx1
VF2jenmbHT2k5XMQgVsJCV+30SggGnCBevmuXIV3p83TtMt9aCICtFc5wdw/92DFzRyZ+0ntPDwc
Ju8KUbluYxx5vqOtSm+NWqgtOdN4LWFjPWuxTVQQ2SbDkGwJ8kgwEd/IIZ7WYDPYyll8tMU2ftcT
Bqx2FN1L5AFHwl/exnKeu8ot1JRhGjs3Qi/gEfnvTJz6q5DobxyiTzsjZWN0XAB1ZCi7jn5U8oEF
//KqQXuDbLe7cdqgPbVuUTtfY6J4x9cEhi9wDnUCmolRxBlyMShXcYNaD8ggK8SsylhP33lfVF7s
xWoJEpUH3KnfB2FlFilmGDt1PfQKmwGN/IdsYpuoizXNJQL2QerqzhUHUBDRTKjKeTvBw2w8VCn/
ngfmkpynBVXFieHcr1cSXOHH1OrF/RK+ruNBe/PccztP6sqtRakVaO+n4j67hvC8qOQEGBiDY9yn
XZwEplmgokxspZ9bUKw6g5wV4xsIm3pRy6EH564VwRos6fgKeFFbzfjXM0HLKM/xcY7i/fWB2RgN
bbE1mOJEHgf9oD4307gfbReXVaheIYtIJYXRhSrBkvmXp8AKTLg7EqrFgHoDZsc4qhJfJPgm/kuG
Pb8Zbu9CZJr+4GJQ+qP6C4jiZjTHuKdRrxs4wYMWnFaImxTca9etvMlq0w+uV7udrhWviG0pikXJ
weUnul3dFYbV/G6I9g3yP6pqDqEGDoP3mlejOz2a/XzE42YZcqX2T9fC5hG/GOqvcwqoeJYnY4NT
7iDT6PqZZfNgsKa7eyelyf5LKKHe3PLS8CujRgzldYGEfZ11MHe2luJpyu0nouCQ41v03p5Lq3iB
aCb1JJDjCu7iPbjjpVobWAE3/uJrracjhiYCo0WLYLQcjGxBv4Xw+JKJRMmZxdXLSy8UpCoKF0dg
VLicvg1v1da5/vRs87p1LLFddDadZmKgpO6DvBa4f2SYewhZ7cbLOi7H9slgG9slG7Infa5csJAr
7+Z5SkDC8ZtAWiz0U0ZpfUltzNFFLKuxhi4R85g9oruxVXqQkFg28nOEDDxCq/Sg2unj2eHmJHR8
UGdPdZ7gsMsla/dc3ldJG5Rzozvgr/9Csl5l0e6BHat0W3I2f165eM2BIox4YHguBMxaCWqEgQ6g
QcczvpyDCIrT/9KVhdjYvhm0ZVbjGY6bu1tZ9SYMUPzqNRhmvDSI+EzykQcJm8S6ijqyJ476G3+h
ul3neXVXFcyTyk8c59qD+DU/w/8PKfCzO1RSO+rO4KuW0+XV74befrfc7vE63QVIZkeu+rgC9plF
lbDJYMMt830uczgAPr2LEqYKGytyGyUQdDfQTKHTQRFJ4Wx3vBkEjt2Hnhs2/7Xn2r9wnOvuiW8k
oWdolf0/9qHNbLGg/L5juuw0tdj7k2/j4KxIb+RsjuhbyBff6fTEFuaTho26TtH7EcQ01tS+tOi6
bx4soENP3685lbiNXTGzkQEQZq0p+0S1RblYWd664VSJQCOMopK4gJIYPAGJNyVhSmNeTatiY0s0
zMHs2nxgB/WH55uuqbk3vg3BtCYQiIdxqMWHeamChpfU2ac2zzfvuZBNxSP0pKZxtB0m0Le5Hxls
GH3ycHz0VcEzC68o5nA9Gtml19dWV+59xJ01oPNJG7igrLd9XLgKOCn3VIT446cIQr4ffMEmqybA
nAKOz7mfBj9cD54Dj8xUN85N8YEqk6O8OHdlr761bkPGshw3KWiEyDIZGwgYfaVbOCf/4Pm6JI+t
tMNp9AxIqnWzKad8vFX8X2+cvOxdi1FGVk7GQuz9U8VJCqvIFVI2p08aRl0QDETzinr+SY0cOHtr
lbQMoMnFyox3mXe0OcQeNUgUeUvZMvx+InajYlFgNAka7nTGTfgISP8dpf2kRN75SX9BA9GmPJOD
qIgcOVYR61rV16m5GnJQJj0BARXfd8ZetCQh1pwC5m0aZhSJ0mdjL8xHFC21NrVM6G8duSSFMayX
PpTnUlid5nm0HCtbswkQXC7+5G3FWjvWWLEeIAGKfje2g8z62yH1V4gfZh8bJnFCR5vfdSDLkN4q
mE+FZ0CoL/i+Hva+rgcDDEXAYjw/Q8eGxsqsTVnbFEN2d3UE+9el3ZbNMCpI8gpZ2V9zpD/XbRi/
l4GQaOtVybW/CEXUMr9htolCPi5LSS0quHJoHWO2tbo/jT4HVGccu0tO8dgVmsfEQSxvFaHB4pDq
9z2HlXzmXwg4uBjq/ve5b1ePqyS1auIn3BxPQjzeTv7c29jhM8VLr/LHkKtv/dpvpi0Oie6iyTk8
tQH0jlEeP+D74nIsyRIxJDIuWBlO9oEagnqrBrl+3QabXxE4K3EkGwGDXrd02FL1ItFovJYFCCL2
OuKYurpJgdmT4Vw5fw0rBB9q8VJmJ64Dpb22sYC8bAdWxU7zeDbCaec/5cPo/fJHFAItZwwQLqnO
lycRC3iZZZLa+eJwAbZt9lp9ySTVLR8lTObuE7F2OEWtQUyX8HWl5WWklZXwKIrt0K9HfBqYBPWr
C38UraxtH3AT2vQTSd1IWfYKtws/g17spsH6SK75RnavvlgZ7LDSYllX+0pi0iSn8D4QuU0fBiBG
iqVVMyqdOwslV08dPelmo8yd/Q7lJDLb8Bjwavx1JZQhPijLOILYxdZuRsJB6x8takimEZmiKV+R
PM1t5JC5/alKExjPTodsEcly6fm+nRlMRnMipCGZo0f8dhJNpRUwqZtIG4Zd81CDtUrT6BafNPXt
ygyH+316Fy77MA7Cni73Y//5a+cAiHJDMdMTIcvUqqS/1qpcrobbVgstj2FNTRNEPPphY2bChwMC
am13NuQk2S/wxmOQ+Dg7tGEXQa8uO8A6dX319R1dB0RtpO651LR23oulEk+XsUcnJ72doaBLMTaw
lfdSuuueZuiIFRpHGwKYmjozocQimkyTg6PgAHfd4W6nzm+FZDovraQkg8pXPKFhgkgJDUK7zcn7
SYLr7GsgZhEmP+awGJjGnPwbOvWWqiwx8SQJMVMwJOmHLBMlML9z0v9Rmogv4aKXrQ9ME7hQ0NCR
Du+iMPNbwH6RNhuRLCxSQNTXxuoPHqyT2ZL0atRsod76IthFS/SUbL6Vr+0oZLMewGcOj4fGjoZG
5PXV9ralU1p/diIRT+RrC1T1aciSvfxvYzx5z0zuDGpwUimonjYaezY2ZNaK9KWPlTMnufyIwR6M
NFjuqVbhTDkTrBkonrKQ1JNx5kR8x6oSpFK7sKVBzPX9d2A7LowxkpCWKgbcGV5BKBj9qLFbBIkW
wqTLXLkeGJZNViRijCSpeg2gMAGevOB/CNjuGVigIdnqyogA2BEriADB4FqixTUOQkTdiuuuDSKV
wbJyWr67GtxqhXzBlhKPC49GRcNYLNF4j3Q1cKe6AigtXNrnTNjpfyy7GtTyg00cQqFTWbPGcSAO
5E/XoTGuChgk/MHztYQpvzFSgNqCCuMPyelDKyhesyumS2E9bqTU89mtAbXJxUKb3GgpBHJ97GRS
1QGCTRjzjEQDLXDx5YFgqpycFssGQcMxCXrbXCnr5x0dnolCFw86ij0E1lMAZAVXlkF0gO6wFeAj
sn1NSAa02++jhepL1PFBd/9ML5+3LnmTLLM/JuSHLZnPNXGUF4YTRtuMBwMFvcryps3dBkaaBBC/
yPm4be7IRsLG8bozhrNdyGp5qGLlq7aTmysUjThTHk7ZWhxdqQl2UpjmKt+ja3eZNvq2KgtygAoS
SxVegy1TRZkCdqqpQ7MEg7b5E8oxCx/7Guh6GHWwe9uta/p/IbKEeqnyilndD9Y9Zh6Jl2pfBY3v
PR7uHfFb+m9lvH4vi260XoYCnMlngUTwAIXoBv1wk5HHx+kwOnBmOY/R3Rq3KZ2SuQ2DVGglTi9H
FePKOWNXHb2FKU+Y19Zt1brcdB9QurOLETyzNHEw+PwQ55v9kdqx+Z+PscRJNauyNHb9cNV3EPe/
iBTy8SnTEXFyS10zgoOgPXxOR4z4g4e4E/8gJWzWyy/HicnsevkbBngr+TlypcUTn76wspx+8JlP
Spqr+XWc1Z7uRxcx8Kblbsaw50bjNLhLYQKW0rHx/FVdsEmhk8yRMnqNIqPp/pMrZUCtYBVnd5in
/dswPg1ejzYrMlIrwcYLhq6WyBRWSUMNLEHG2fMUHNgwg9YwYYIaMryng2Le7SpRPelc2cwZNUl+
ytiU8pYAyoCGA6pLy18lTqOXTLugBl1mU0fco2tK4J2Zy3Yr7wEZ+YwLYXi7NBdvevRZaM0HUDOm
cIQRItdNG8XKdAoRdDj4HhaPs/0BY38PdNvi5S5wSweO4T69E61IBgFXvTZx58YvGPsodiLwV9Aj
A/wiV3P9rO6f/WnuxHhp+fwx3IhkdxyEbsr+Wxq9FCmO4M7hy5L6DwU3luTEoQdGvXJKB+6+M+7z
r3/8Rhl9jUoXPR7bvDE2nFQRnH80/9tHaioktjxjt+JC5x6aPL+Yjtl+5FpMjmsV7P5nBFYW0N/p
2tAUX+wINwGu7bFTO1BM0qRhdn1765rK6vzvk62b3/byowoSgtIyBl0uYXaY1kgR3VN2aauroLu1
/qddQNv/2MhKUcXISyA04EhQgB5ydCXGylHB7/hxbGc7tS6y+df4E5YpOVAHGscf7XNjsN2UWSmd
59gnSL9Jf3glSOArXDKFYEvsUkdRG6OxCcXow4Sc1cliQ9w8JK54bKRxyL4gTWn3g7igCLWOZDTu
AralgKUC0LuMOH/ugTBeQs+GO70GhBpR051MxFKiD9M5A79RFMmcky0XtdKrJiKGGTVuxzlHL3Zh
Vd5D+EwDlMFYm9gQ3OpO7kb95R7S9UX+ncthlI0bhuFSJ61RbzJT2P+l9X6QPiEu2xg4UNnjCDx0
+cKBXImuIkzTjqZoIs6sM1+rBIJ5UuB9EMoX/fGybnulJmpWZ7E3XjPip/N51l5LsPxJ30uTcYcg
GrLnrRLCKzK7Ct1wT/Ead0wxH9Vop5opZSJdwxol1uOeyrxE0GjESPKP3Ll8LLHkClcDEAJk9KTb
Z/iFnB6Rq5EiiB47dwi/KBO2Hh+C6eYxFSnaIFI90zwSQwKZNgCCgJjCh/6cGQV7BpLoYfV7tXor
aHpkQUiP2QXdkLdIDwXrNyQwtLZsnlx4aATnpWLZfvNDt1UeJXBxc0nw7CRLCF9FdjsFu73Z4Jw4
RwZucuObRBw3cXngcWmhZMV3r77Xv2Eyafpk3U5Aq8TgRnNZONEaJBAe0PEVEerekCr+BaxnPRND
brdVdachcXt/FHdytyA//kbmevEd3fD1Duy01oO+6PWOGuVIJMYCrFjGRXdP+cGbavWNVoyKID4u
LeyWNUwqyLVjPzs/Aqzs4x21QJzD4SFZPmKG/NhMoDTR4U8DKw9ODV5UYCk43WZicZFv2H7ZsUcp
6JL70WxYz9vJZXD88BQHmibqb00oXUjm7tvC3IBwT2FLn661rtnEq5x6KliqIqbNWVHMalcTmcIX
fhdWJR0x1DlmplFkw0TyXWja4q2ORxSEScOERGHTtSNxM270A4RHlWE8SGqTu8Cb8ufVUoN/vdpu
PUQlnwMUAXNx7hFQI9ErQNdvpnSCXuie3t/HIJLyJU8DNKAM84dSIltlrufXspfKJ97KL83xy5Dr
OWEqou/fr83HejI0/MI+d0VApNxfRpbrSyiB3ZapM4fMMcVLuWBvCdfl95YHuIzbvQvqaIIb/9Hm
rrmKzJ87caRTf45A081XUU3Ad130zl0bZRjYL+T2sHpFE1Vt1r1bc69I8UEQtPEbKOc8f5J3T6Ag
d0Bp0VnwehJ3ohsoSuI+i9cFB46RKOpOWhTR/JIiMKxlGevDNfSg4Iujh3fm/c8D54cqq/9NVra0
nEkbjjIz3KLc954MrTfwQ94h2ySD1fOKC963v9Lk2puzLwXDkCONTbjDyYEOEkH3sz2Gq3XX57cD
wi7PbBMuwPmBBFqZrDWa66urcA9IVS5dWgEnM/9WE19gc6pNWuaLDUNV73ZeOBH6Wu4UE2xZWbzy
3s46tzVh/JD2rjWoABD8oc/P5mD67PqSxu9caZUS7hB/jsx9looOEWDNcYg8C/85EMBxPjhBSra9
HFwixFEP0GvUirzJpNt6Emw4O+QYVPNPHVCA+bgE4Wkikgh80zjLeUiM4RIG0Yvx1/CNmo1cdZQl
cOjV8tacVxfkZ/ET2mOj7qJ2prqgfimiWPE7nAcZmcGNz729Tm22ew74JtimxAuYRBlJPOECW+JQ
lbX7rY4sSQaKUL4xKAKrCSS24kixpTmEtStAK+vJSGLzGvsDqbm3r1zQ4bsgHlKtQLCjTLeXPckL
fWsZPS6vuM2eQGC7lxslFbOb4HqI90U7kbBa9etliWuJdlRiIgEySHYUCQES2ebhOmTp44tAXJhb
ckEfLrdk26yta5KBM5WEQSRt3rRbAsrKn7iB1D3idEwRe/Q3gsfXuiebIotCNc9jg6kV+juIJxwU
nzcC96Np3lMcdv0jFHngv2ZuXS1D1LtNsz24/EhQFwT0BRoSXkyd0XHlVIdkz3/tqUVk9LQG25yC
mZWN/kXrDEUHDK+afM2QAKGT/wlLZGPOJcGNbq2OEPay55t6dZqTC+DRAW2ZY9HryCLMpkfLGTLq
yC7gxSu9rq5qZFbnGcWJFoxwqT1roR6DIYA02KLZfBpr8b1OXGO6YAXdjhnzGY25BJkshDZQphLf
FEgIth7Cf/+C8x9qryFQsUj70+vAnyrJ6w3Haw3L43RxVeZPkJUUrW3mS7t4x1ZDi8HBFTWnaSiW
uji2T3Ul+RNrLJa9kBkog1cs7UhHbP4ydOC4h/9LRPEwMUf7zQ1YepiCmS+k9Y6CfkXB26c8va1X
OqAOzZnPYmCOJHwp90eXy73+p4BxwmsnWLf9P2w3Q7l6DFVlbW1L+5FADy+wc+7BrxHWAjsnX12F
AMRQ+SUdD5ctT/OjQEE3auoIYW6ZtVYsOJP3k2Y/zKfS8j7OmV8C62KEQradZc4hodwU/ED0d8cB
i70qWf2kcdGixwSQTW6NHqSvZKf/FSxy4P22ZqCt1noWk5In5dtAAuYpjlyGgAc1sf5zbo1HN01P
7k0CDRkzDR/b1+9wDOFGZEm9GW+S8ix4BOWmW3errBQ0NjVqja1uccnkLH6WugacwBVDiS8nQ2Pw
CstOOSTFur3E4s229e7eQRwGpad63UCyNs35Mc9ao3YkJqMNe0waMwcdLHU3oR1zdeoiHvf0Dg76
zKQ6P0kVJ52Efo9WCna8y5X3W7WUYoVrW+LaXFBZULuNe0Ddco7tWOqhW4TTiXvwnvgrYgslWpAf
uF2ncl2g1n4pu71PKBdirzAmStkxwbh/hQu7QONNi9i9TfxYuxWQXPkjfuPP8Br2jJb0afaRFHW+
+tNSG3A6+XfnJMRvluffoIkeOwFgl9IKDhbqOexNxc3PasZ5qjZ3yjNHKjhtr7MoWysseWo9aesa
Dv6Oned0xfbatDReuXXLclcp6d2gVyhSFl3pNCA6AceGVDhkaxZ9zkzuiX/15fSaxaHBsR/zHH3p
FDgM8jQmctTzTWGI5Rv++eZDjrVJrC/ZaJw4IzHgPRKqtCIAhuF+QUReTqKHCCgZf4UmxLc4wMz1
DAiOpGV4Pyd+2ygKKe0KKA37wyJ7rvwsdTWkQlE94vh0FFGtkmYYUR8UJc/iTlFV5KeW4efjagqV
EEHZ6ckiI4yhkve3z3UVTHQ92NggV2HMa4fiyttv2fT+R4FwdJAP+aV8lKw8TcoLGJVk/lRzxkEO
DOcFttt33RHtwoZ8NjqfAJ4b4+nvPy5kqmvT7OUTg1bydMqEwHxqq1GG6ZIP6Hf2Dt6DlzSAajdl
USfj6C88z7cMKZwUjwzogKaJQEqeCZ/lTi9faHU3n3L13KSGYj5Dx3hjUY/5AFzOTZ2NSqtqgnKO
hyi3c6MiTY3VoZ5LOtfDhVwGg2CSMkPjZ5JvEQKw3hYEfqAW01GMfFJVyiM0RAEjo1t1we9tkciq
75RNl3XkL6Y7kRMUy3zC525UY/UgPajNm0Fz1D69n+YZHcFKcHi0wradlqbzYnZHX8/ve0gpO8fS
3NakOKt312k2JALxdRSvQcCU5rIZWG5wJZ2KR4bmZOlgcEXu7w81A+sqGa5DOrfapxCTbWbhfsJs
Kzp3T9RbKtxhrteFEYB9XWfzbVdfn1eSPV/modt7ySkSCcL2jnCdTVzpqbwaTBmruicqcNAuSp3b
jcIvwHyG6VAYR/20VQhNV/SnimGhnd5Tm+0RFsIIpdJ9Di3l2yUfsweQrx4idqMRpCZIR5Fzw5fh
L4qYhkIdKBWmNnnexa6l/dPU7tAkGINs5kU6YDRiIKYf1I97yM36W012FtU+/ufWOrxQbZ/def2i
JCm+4dbzVTCat2tTzPTiFmpSMAra2abtD8XMw1mh/UNi7laeD9f11us8mxP/3Cmy5AgzPAuesStf
O0vw1cnj26eMkDAFLKIPuBw8arqSh3yl8bMeuQYFxoZ30INORchkiQLfTIH9yJTx9cRkJ9KA7Qv+
v7NjcbGLvxjLkJB5SdIbBnXxWclg5EMfyzYb2e+BWZjqgLDOVFfzv/JBHO6fKpC84/addalZTdMg
Y4dRts9Xp6vCTGWKnuCrF4EqoH5X+yjkUpvJC1VE2bqueNWcptPgZ57OwvFR63/DQo0HMf5FzLBl
s0Z9OS9EEBWySHJNihcd2I2XVh7kwmp2fx9ZqS2H/YirelJ6oeSqoTm1TpiECoa7Vc/tD9KztTvM
9qa9GJ1fmoDmtdHTJCtxqUu30qhuo6XxVwhcwDSq+6rv4P4T8vTAPBTkpGaf4rI+RBqm47xPo3E6
Ktz3z0UIMy6zVXwGVCj4mwJ8PnRR0nbySNsdUr8+svwuTkE2UignMKiD1MkIeWiSfkDXDwAbASUx
RvmE64iS/DBKOZ2ROY+fM2WOXzx+HdzvJ6N77iBg6QGpEzKFaSi/XF3zsz9mN2yLKadL39jNYXNS
B4LX1hvispfq+yBmCwSYiW2WSWnG0nKVGIzD9nxursHUz6fuDjmUY3vB6zg+haqnVr8OeAzZeC6N
cWHaZZW2KtL6FPB/5N9N0B3NCVTXdweicjY85Kzs0zoQzOwbJxVU7ve4GPnqQfyKUIJP+xQls4Rj
Hy7zxFBiWAJVBbDJH33t+0mG2jXHlR1U6enExdX8pVURP1WZCNYoubN0Jm9F9V9NZ0J4qSMcuqDD
FXaWqzbePpHt08TlYnVwufrj8MJ2tXpdI9WuUbKZUk2737+D2ALpIYwwE00AN4z72X5YLBZPXp4e
FOkmoU6SvlJRUlzAqwifbalbfl3TL4VbYRrAx4oQs5QL3LX3rBAe0QEPCieUlx+rW40lQyZR54AX
EwjDPlIWncWx0W7P94SueilljehFbUOm5yAgruBtc8oLZhNx8igGJ0LfECMyqrvVNxrykF3Fltrz
O9K6exEVUXBFUys0hYNOxOJC/9n59wSMmNtVGdoDhZMT1VynzjKq6cHsxr1gq4Fyd/AeibMdK0md
0NxZV06z/DouZn45wTbcZnoGDkhg+QGt6R/ZkUwblhhU7mzMygRfdVwXE2EP5x7z0VERzluYfgL1
Q09wIWUcH+KGMc0u4pX8+dOrPZtfPKgFjOAzgN9Acfu1xGZ7CgYghojlf4kvDIfhN/PGHjBiYVjz
0PkK2tTYRWccnwwO+GzWoLcMrbSr8WITEyY9pm5OfqkNlM3OHsESdrOJkCJlVw/5Wkoehsmd8cmJ
8of0K2lIUxPfYL5oDBgEVOLvOfCkfbsLe+xrSBVdzi47LY459RfFhxJAc+pX/+CfRRsfjpdilSmQ
/X3VmVSmRSW725ygbHmnqrWrbZuNLJ3pQvgbW6CH35B53/TnJbEK8MkH4TFc6x/UU3lYYfFs1tHU
Q0LA8tU1+CWfVMtWuha5Xce3mV9FfXfEiw5Ed1nLQSHOXrmIEnTuk4cDZ02ErQbf5XPTv9+FvFhU
18rmJuWUJeFZUmy8WRhqxLjtYRvQQ5Lu6Wh5YvUpUu+sNECNZ+q3wkMqQLCqarAAfZT7bN7lmNwW
dLDqvcgcsI3ORlfLQ+s8k55SgLvpfA//0diC0ElxX/iSydoUjDHK33e9wizu3SRJrhYX/fJPbNxV
gwSbHiUrOc6xYVO2zkLzikntpOCmjigxW6//OjgIcw1Ywqqa8mhmUTqt5Cz2ZPClcBFpQpWPITtL
0552Yb0AS36wZtk7Ce2dRZp5XqQHKPzisP1gcFZRAFRpty9jtvzRwLAHYGpl5qSUQEu1CQmgAf63
cjVud0Ax0VyMVbnqa9ww60/xVttF/+5buCC73U9y0ZFcE5YXYck8VEYDnlxMtJ0oQgay2QjPm5sG
Y6ZjVZakb4babCx4XGbo4p4wizob1h91sHHhG00pq796M7sV3SOmUZIrJqJxx9uPYUiuzZ5x5z9w
6PVJMQPO0KdCRk62H2Xxn1S6AYbxl4RflP9seZn3WA/yppWe1j1qjSs27R7qD5rMvKFyqF0xerUc
NGHbzoaX+7aMezfazKZ1Q9oMHIpa8975JwC6o7nVYwtSprzdPxKQMtGkFvRMiETfauI267QKMd2U
z2Shas/SIQHUIr2tfQgbHd2LrNMjH3bNUs9PyjMiCTfjUZj49cCR2dLH0Fc9Hd5bujX27mkmmEs1
k29OYCRhCT0Z8nfTyKUQsizlkxdMuAVb+udSyp03LlOzyyOHtRg5ivdl//z9uFCrb3B8A30FH3EI
Hu1ppSSbl/Zq56zEgegFrp4+T4ji9cMlK4Rgmao30wJgk42OaHXXFWLf5mRU/VieuqC5TqWbLxNS
ofGfgSwxbJhjAaWLH/vfTRDjAub+0qaJJa33kUsdg4SCYf9mXEiGh7QBd/D+9LRgfKX04tnzX5w1
EtcShr0n7U5ARWQ1sypVcnAYqAsv8dFiv9YLER8SNoDevTSnih0NkaWUNmwsh2bVxnJ1E9PBQLPb
R+bAVt5dGNMsnjT/r75c+vqME6Q2jPCufNffzF2Su1ALbTAj6/PWi9QbG3gOy91kWZ4lVLb5iITA
8k1qg3i2NwZA/i1D+r+Pq8MGq3VGkcc/vIkKxVSTgEMp3VMEzF+h8PwnoE05fbcYcS0oX1gX18aC
4Dxrn+VyG/kbzmMeCzlN92Br8LA6cQ9X6FZMEDITeI+Hyiupw2pljikRBAVs20DObAvsqpOyPYIx
eDMhOtRLzFaOUhN/8ZD3XffZ56IXs2X52Ivhsxy+kIAyQRtTEdlLx+LgyCXuTvsHeSU1xKEmYuwl
bc0/pPMgLYU7+Cq3cEEzuN77ALoC6nl86wWdclKDdBqylY3dIBoFM8vty2w+K9Zb1KwCz2Ik+Ynr
1w4BgZAOy7sCVT3G73hG4rCvICUbdnsKrQ/YPfgihP7SY/VI6dSkjmU7SnubQRPeyru2FqeQ9shu
zvbu8S60S3XRqBpue7v3oWpQA40iUcxgzXlxB3k2GwoZHRcb/FMCQUQYSjY1hQ08CwCY3oiW+r3c
R/SyaPe5cAKLqG+y7rxALglm6N2NFxZWHfX2C/b/ntQgtW0yxw+fvw2V8/wdY2s+RgCnHtUYWSM4
0O5KqXSdHQsRMJTTy5IuNv/iTy+X3qqS9yRCa1tqWbEt+IlvKh89jIwILanx8KQ1DWRTJ2SUeIkD
JEdIsUhTKqfMUTYI9wh7/kJq4rJPEOJUdOo2J+85WXV3dgBLS6C6YAAkDvwWx7RSNEQQfQWQGscA
a4ZTyMNMov4oPJPRZanQaL+QO7uIrv8dZuKktsfohqTjf/u4WYQmHS9CgmNc6ggzGIAQO0JY8a61
AWOIS9XN5dJZsApyFOZR/VJeJT5kGwo+Q3j95WPxxrSZJP9Y91XkWrdRGgbEBOeVjO0oZEeoxD89
8PfzacprUp0bLVX6nhEZn9M7iENJ4cnMs6PmzH/06gPaFFfBOQwcmBaA46sqS/3zMc33jucomAnl
mJ4BFEvoksE40Lz/HovqgQQAZ4voUk5KRK50HLe4G/k02VMSCQ/3xxYJPD3GJ6GQfIEhvX6xzrtO
4Rx2/VxZ+U8t0kzO6F/CaXnSbMy+gH14NzrtGSB41l3xujFJZQCD1GBPWpZsx9LftzV2PESG0BWY
aEP64W1NyzsQXCmkG+QPXFh6x/PcX9tASr7xdlcCGrSHpM0maRdRU49EyBisn/plbHdoa7HRbEbJ
dwu2ktxRfWKZE5fENbLj//wkXnfr/zwe26FZL+To9FXsKvnwTh39QaHzeYz32LV0kqZmtajvYMP8
5zfMEv56GsPeU+8r2rj2dRlw64muXtvM6XphGpv1Zu1fK4IA7kOJSycO2V+a/9ICjA1jdJ+tZOJT
npkFH/4n7MgmJE4yItqi9pVQE9KMfg94jgeXgDVF0yn/IQJkJztNj1ppLN5RKRz0ymWC66NjV4Vz
bYQMuJ5xYAbejn9gSkxtok0ns6HeAkFzAc1yDCivsyVmxbHKJfwNPGFAL2NNzoNwyD39OPGekud0
cuPZSsjy1B4Xsn5s3Jvm7+U3DT3M7g5r1DoqT2fD17SxXMpnNBBRFP7ocErK/VTXiFLf1tm+vpBB
160rlsZpfD7O0ZAII1NC9WMQLzHkkWOFFNDVcDi8UuwNmA8oLAvW2yQKBVVqJbuz3FrRM2G4Q/dx
pLLtUjQSvA9XLoyg3rrxc5B7mSzUzBBQc8TL2jvx8C1e4lhtnySm2TAPoJPt1ZhjqLIWOWEvjS6R
bgO0eruyUbsF7vRK2LsMVLjIIq2wFKLzVbpt4AeIozuJHc9Mho71JXLKd7eydQFGxtLYg7hEjVZo
IOyyKePl/Ov1exnNeHaszhS1ih1Dn8w0zoGGoVFZ3n0Hv/WG4FSndkdDavAVM3CEBB2Hj5MGv0gq
gFpewub7zbKl76m94NJDENQJoJHULsWfxghrItUu4ttSBDYVPPrFm3cOt1zSYzr7pQlxuP0SFUc5
V7Vi687iPdiYvEpBgHD+Dk3oNDHop7N7d+pgeSgjFcAbZwSUF+4g0gVKS5qX+ifZY7z1dD3HLkqW
NXqMobDLWbmumc7spXFvr9ivlx3yCmHomFDuao94BXEHNbGsb6t8tG8XeTWD21oDj9mZRU4r2241
txJCRxEt04yXbdoV6eROwNkp96878+BohagfcOVSIl28p6XFUAGcLituGJ3wcT8I0BPv2+ZKfhGz
e9YmmWV7k+PBHe4AoCUqT7Tw7yZt+/B4svGlFBXqjpWyoCGFAGN8AquYLMqzSqSHExcwXb2uCwST
9F4OskwTib0bC2Q2L35lwDtuC+pWIBxgyO2n5ZRN5xnWiGZ2z9qHoXMbyUvuFRXF8yUkpoQjFH8/
bG44D+cCfl4H/WDxq8mR3DTWzofHg6M0HhTqQjd2Cc/QhNSx9l4fz6wkwJmrl6rWuinlHKCqPVP6
kX8SMa4YmOAl0PDkwXGFmfSsjYitLtDhFP3C2FlCaBdpS8kQO5vKjffju/4U+FyA2o8AMdzVqKNc
teUTQ8zaoQh0+oHav/Co9MMJS2Xx3Tjus650nDAX359T3VxzHgVsq1xGfY7pAato4EAGiSXPlFK4
KWiRTVM74vQilDU+4ZGeWcIiEkRjnQwKeAIufd1ajBvZeESAuZBvFB2cb+0QVNEcx9FMwlOUhZoV
E4HVaiEFWo885vQG8UwN5MUNlr6FQlMhbZJsYEdNFZv5/BvabNCcMiYbe/1arUbM1rWZDG/29J2q
WNJave2aXBBl4pCX1UxQMXuxWjy2dGihPqqnuzscmDAPGJ0ttORcvd3CeCpYLZv+pbXLtP2dEvXv
xSt9L1YcwszhAOGkYY2WyhmdbthKLHX9wEMtljeccJut8l+ygKcsbnu9XyLJJsbJvRSCOunHXFBY
XnatIu5JiBzVXzbpeQvRWo2pEDEAC9C3/mswFntI+sCSEVv+dj7wfDkcAgAUcaFeQK4O9aO3R0N0
hfvanpCI+xrW6koK0QwUae7d5hK0QqFvtcWOmJbmtRrG3l6u91fjE2XVoNhut0AdJtJ0MSqYOL5W
zchRI4S3T5FP9jvHCDHu+1gPb67V+Uz17GdT5AluWFQ//VmvK9X6u3tWJ4QR3Kns9oeJn0EmXmij
5zpR6hIDxFAotlkrmXTuja3CX+NmW81vZZTes4zAECp+zewsRAqLZq+HGyXlpdaKWznU+0KJFe8W
Jj2cMlg/2rA2JV1MT+/EXxPxoRRunK7/zOm1E76umMJmgJTwpr+q6WgpiAV2aCUQF05u+Sziisil
TnJwQLi0EcoZ0KHjN4rRHvolLLgcXIcWx9zIR5aSGCw/nQRjiKn5i6Ql0OPmsvAhBvBnBSdNUEJA
C77aqoBBlhJJvFqXn3PaP/ZIFrHV02YKBD5Aj4M7plJ+X/bAzjWeAv1SopXHKhblK8PbvYGQ2A2/
v6vEVTWgRLAqfkDCV8UD0Gh9wAdZZhVRmXQgV6/gelLrntMQz5REAXnlcHluWY+qxNqd9rA6YFsT
qeg42aEYoIvfdZG0RI03pB6jyC7b043tGOnnJ5UT6X2ycFV819IV/V7NlFbc9PxcLjzGhqRN4rr4
61SVs9Qa/7Xg7R6AElvXRwBBQrN8rcIaUTHT59W5pkET8S36ZhUBgfObBpznwv67pdyA/34CUGJ7
VW/q9w9t/+FIq5iEtFIB2nzMld3pYLV4OIuiyurozjVG3dYexyby7ihIE2vo3P+ZmgxQvx9NXesh
4B3QHlDyLI6B/8EoxSU9HONIQjc7/X4cnhcA8QqEXjMhYaEr+HOMKn98xlRffGZ7nEXo/gJYLs2Y
95z/XRHviu1WbIJi+4DCxPq1m+R4cQs+2p7pNAMuVSbrSt6n7KUAl3WtKXR9HLASurh8XLkkyb1I
bPcF2XiVQ/uV1PHoWmWpVMQomPEJe4s7h+QcXOMI8HujlPjwJfoCXyCqfnB+Lw4dE3bEdlXXnsgT
Tt3I4dLo/iTuhcNJcT/caf9Dipiz7/iBafZMUkwvW/hlvRztEeHitY4iklVsjMNfZd4+el+3yrT2
Nf6D+fz/3zWXxdxVtmdwyYWZMl+V8Gb0tLRcIYhCBvOJw8lUeGeqO0LEcRRnS9iPAFAx9bLXqgY9
qs2SYulsW7td731B3+IFArwnY844vGXxXJXWWQUKzE2591jmhjD51drYOHmUrSwJkdl1JZ1gw536
j145Wm+qeZe2F5WRHHsCHbbIVRVWoyGE2AOm4W1rM85+AWzC3chC2shpoXVsn6Y3UQ4x0vB7ChDj
K94GhdaMELRCfWHBh2MDgOZ2qbXBP9vHPrLRIwDoae1Mtz9hAK/6y3hE4knCdPtKjFYjwEZsYvoA
LO5LwDd5aI7CKINiUr3OjsnKIy25BeUiF+wRo01BWw92kxWgi/t3d9E+jf3DrflvKxvvFFFQEN/Y
xXXcLTeCDmpiefe9wi+gqzJkzjy1aUAYmKqEZHrStCYskeDUXHrQqBDU3ey7v0o7DG7pJtiXd6BB
leRDNh2l8/L1HWmoMzMvhNkwtlw9gTWnq5mwrcQpT5Y32eR+QeYT4ydTUkLHbHOBtGNvZTut22Wf
LebsF7t2Gw3rqJL11RduR1+1eNxlkP5Pe3wIDjsa6keqWKczbKfdDffWuVqnKbpjLuSBndqtyqNx
fSVzx6S+zD9U5SIwo8T0dIA+gWFG+Rds6cYcO/qeD/IakKCSaoz5bV9DFipuytIUTeUoQ0r7E3ft
BGYjKLehMBB/m3/GqNglmtbuuXFJYDFiCDNO6micrSCqoS7EU8saO8Yf7wm9V+S7IYYmDz08FJRW
nxot4z4g7kFC5zdxFDAVTD2rSp9wxkSV1m8K6DeTjFzuTQrTvCItrg9iIdaNKHwYBpvDNGpDyrca
E2uUC9sWtTbAOKv6lp69ws02yXreM/CqyqV8Rv90TPap/Hsi9zSrqRW4u00KcbtbcfsFt+1Yt3Nx
eB9L6yv/fCek+ECHObONb5ih7kCMlo70BAx1MlkCDQUi3HO+9sOKlvPpEF8BtT2Ib1bPBKsEGN2v
0LNW/ZcA0yNAfHWNsw+jFx4BIlAUj1LR45HlNvW7gpHrDbBK8zCjSSvlaoZD8STZO+ssepZ3paRu
wtzEpbIA8cwjkfiTRz1HxHpwqpEfaiW5S0gSDvYavXj3zBtfAVSagsEyZ+qNUKJEjwJFMMxFa9HG
NWG5eh4C5owtCyoMEddh4N9o3pfEz7RRMBJnL/egmWyNyLlA/YFCYCeoAqxWUDxG7FK975cQ5Hmq
89EIQmZdW6ZOaxqVBh8Cd9v0qbCt4Zjqk24qcCogXC8IlWprcw5fycklMVPHCfVnqsC4vlH29Twu
MOmiPZpImE3eAFUGlgQHvi776hvRLl9MSYjgGDHIgXZ16XoS3vT8ZwGTS0In+2wmb5SnyaCDaC13
tVZ8gOdQkQZzwCF8/X/Rc1NZZ18Kv2eZTc6+Gg+AbosvOgmd/B/vrCKC6cOEh6wpGgK2/eicdrc6
i+Qx9UkLdTvCKR4nZZGu/5D2m8TC0MCfKHYJJZnv4iNPyzb75Wa9o77YfEfZMsZKQE+dPvPw+pE0
lfl9a6bqzFnXnBhbHepDJBpfcIIY3OdIIt5hX58Cw3x4RxJNm8nSyKTnHpq/vdawyPxNxHxl/DW+
pPXdx19+Xqe0TYy1Co4IXJmdxdWsZ3drtp93nuwD1bV1XV5IJKt0pzAQ8Y+g/62mkx7VRNzVBhP2
sQtDmVp8hBZsLaVD6n2oeZUDF5RNgLpURJR7HwOKpzjVJc2Pj/9P+6odR4F0b66N49CwfD2vnbCw
nuCoCSZlCHT0S1K891T1sv4uVj7kVJU13ShU1IkcnlUfAxjes2FIeSN0xTnunT+ValqDeRFWLCWM
84/MPBpNccm6TfQxzXNDo3aMeA1OpZOGmwXc7DX9Md6nFnJ+oMSWIcdA1Re8SaFly/VOKfvmtX4P
zEFnfElHMpCcJYR4ECJLgiZLcpgyZZ3WsgB/hHLDOk4ftUC43WHSxmmp0RxoU/w7jDv1+W1BlUhR
R5eFrg3VBGRlra8AZAVeLZDrzj7US7otOIC1ivWmp8kZXaWPRfw7WNYyAFmYTBck8PurZuH7Kejp
e0nEOpOaOnUmo6+FAdjxSt2acm3DwKFljgAm9CYCCRtzsFWUvoTeCHd7UXAga6ZRdflOc3FFiB7C
Q/vyqRKP5Zn/OYQjCQTpKZkkddFVfxEh5HWWAb9OwIvTPkAnfmzh8PRcY+oFoe/pzCc3jSakarpB
ujEi+AXvl4SddaKsGyvoWqNZUVNzvlhtXm4CiUATv4zjwnxCLvIzVDpayOvm0IC61b0fQ3P6XJL/
x5S8hggEtQ7srtW3BPMEYsKlthYfbp6J4XDPX+OKDmRNrbd/GLf61I52UnmPEpSSSVtCBMwGPHVG
dskrmtQaDQDO5z1nIXyCNH7aJ9jCRRhmZuMsAcusqOPnCf2vQfyhYArGsXG+RPNzepSkhF+DKFK7
YWpWRnTA4Qk0HDXlz2k5XADd6vVY34xrolqLxRcmLjG3CRhzAgHeF3eyhNKcf+TXb3/pqNYqJ1zk
gb/rETxjc0mwUicGIKBmB4Wiu7b6bGJYsRZTW9XEbdwU7dFFXu6EwTyJEzsEn0KUC9OOsYqreAEb
m7jZSB0ua6AdTPtF4ff2SrJ/tX/Ti1nuTWLCryiufPFmOkgbsXQQe1/dL6aq9DgJB1HKo5dkXbDp
vdQSwlklWNIlbYriqbeQ6zNaip3m+8PCkrAAjGIy1Hy6oMoMmMTUIwFKADp+uFZ5MHG+QxFLq626
n7PFK4QSgJmd8fByWXxCuLkIxlcAXSkFxnCsF5pt761wUU1VRcXnmpXOFBf+by24sUw+FELI9Hy+
qXyxk8gy6ofxdwegPBGb38G6oF81g9sQFztTILiZm2iwHy7pSsb3Cc0qBXRYp/bT3zTIm0fGypjy
Ow0hK2rtStP9qOj6d5/t+nLjxJmo0aOwSypWmdVUtPYKbSYiEKvgxBl6svxwTBMawy6jUFwQ7Hhr
NGAvmcYhKXFa17yCfyYvQgWKYQY13aCyTucpLtYCcZXSbo1+5dT174tsMUWP+7kueqVlpVzTWS9M
W6eEdyXxK7zDfSXwQC0hEq5KBcN7bnPrZtqkMJLpA6/AKRthJ2XUpklD+yGn3SD5kPYRgY5r+odi
596B30jz2iJnK5WHsSTH1i/E4oSHdOQqxz7GkuRo0KTuqAXSyVnaAsGW84ILH/epwqsWoLLoHPLk
CBPuqWLGBdVMJ0hILUgse2+esTVtTp7Rc0m3Jk5FS9uGppUUbfQuSLmWaDAHy5AH521G9mtdR7BQ
7vC4dG9B/YzAM7bSQvMNGs5E552Uy0v7zou8J9DD4/fqk/cyYWZFY1mDgWWdGX9Fyz2fppbHL12W
xYa54XPXDfv6hnzdvZMBTdU+UCxjiDcsDrl152G1orIUT0LT4SS40wBF5mX15s8PXHX+wXXJ7dMz
LL20gdcaMHL8oEfW5nW3hSaiwDu8kAetaOZ65Z3UE/bthivCpSg1U3PxqQ0D0eBVHt5FRX/51432
VWSYP8el4r/GnBZhi49AIWC8fRGCG7EzBpP1T1sAFnKWz9gEa07PbizuS+clAdGPfENJbi5abgqB
gxJGb1XSvqv4dpuPu1OYLDMNliZFjk+a5jPn7mV8xsXLp4eRFSYvEPR8uFV4rK7ZnikHrx1sB2fe
POz4ae44vzxGKfw4bLgm2d43slficB/kD96vboglC9Ko2Y9zMjrUOTp2dyPnJvTTdhghId9cs3va
O0ma6gTFn5Ux+hQ9AZbOtiQcvvSgqzkaYpKXp36gu/p3qCmYT9F447tFya4Q5VUesxjO8GU0+7QF
9k096iGmsjiv3i/QHgqK6O6TFffxXvG/tJtTvIgslN8QH3DFeQvuzPUhTMni+kyO8Ujf5JF6elri
pK80jVBJT86qZqUPaIOX4twhkuWaqPgyUGXBFDPsqmwlOBMQFLaz4mjgCnlJnrD55iSOUdT2uHDi
62zkcf3pBQYyMaAH3yFWD2b6Reisrei/wOKNbG/CELX8+ScujShJJGx+DYbkW33lHTkqvABnb1Yb
gl+fdR6mEaS2dl/tdr7AdvewBR/DbA5m/vwj6tk1pUDI/NSPLmeoYbJjYJdVOtghi1Z1IA+ZhAwN
S0rnLQ6IgCGW6ghYTfeFf5MzCFsC1sjJe5ZfISU62KQdJME+uIRFka+zCYOql9two0AbNcmkwVZL
9iPwLXItnObg9dXCx6uKdepSWAam1lqCiP0ZeLfa76lkwu+B4kYS2ogY6R5b7kpIxO29cmOjV/TT
9nBsaXSdqDZCQ+MPXDEdkK4t0sFZpaK/QjLOmc9hIza1u9zM7ITYw9z2S+u+I8csGbGAYmeiQgwr
Oy96kW9qEkISZAUiWSSTwFeOBLIOL5eWVUtNdnWx1BIJ6WEFrhGERQZZuvZqEJpGRktWTRBfU1gW
/1VHZFqW+08N33mFeXfOuPtyi2Kbn0jolKe7qmb21mu82gDLh5r9jVo9hQqG+NSWBh0UsA099HL6
+CxaKpo+NtVSFF7Hqu+oVG5U9tX/m+a3CaMvcslTyAeyntggF15c4i7Fu8xpV7Wg1RyvXZKpqPMz
2BuY4YcY7Plm89vD6Ji8bhCq54WqsECY7QAtDpIv3DrzZUGq5t9oApp2SfeleBx3ojyjNnrwldc3
Xj6t4JeKdXFeNOmRanVgyxsGQPYGa710XdttPCCq67ok4xA2WrV34xRi4+e193/SP7EnZmccvV5d
AMw1xtDy5d9X0nKFASSNqB0p8nc3/PpwguEAz7xqEo/1a+I99mo4U0NUorK7xnUxydGw1QAXnEsp
frg2iwOPAHHW8M6LOJAElDjR1nPpmW8dD1KqemAWdLFqeMLnmSJ//gAKb8tNFBiKZmK9Z8/yTb9H
ycpC2zxh0lgmEIi+/eHGLBWYtRoOyZzn79Pqgh2o7NDfg1FopcamqOGdjD1dJOAkAEF5bcDQEih3
OoL3NDtVwgtlVEvBqM54LX34uMyKXZL106JPj42KnGmgm8ABEaV35c0tDnM9ld0+zgWI017UXsLP
pcAH9AFyA9mm+o9jXvrcJEYkKWwM5yLGtfQOG9RIIq64+IN9bt/y+C2cHuAPyRk54V1ZgDA9zSiJ
PZdIQa55KfbBPZ9jTkaL/Bb3O/xXiPF3VxZB6H9x7TAIfRm4r6oto8GuRG95W1jsF2UsGJEvkxOO
KzHSqoenPZc1bTLA3hrGHsrKZ2s+af1jq7C7j9X6933ScPMlnVtzfdbEJKhFkJ9FDS8yxJ4XiqXe
pXOerDCpTcHB/sou2y79zRY1tC6O75X90XmYquixYM76dByOfRlQolrKJSV4SYcikFfvI3tKQRSb
zKzBTq9dWXJ2oJImbpEWQrkXOrmNUPfqXyzFnftws8ad/aLtn3IDMj6v6maW4RSmtMB/F9pUH4mH
E3ceHXKSoRmVeszG+x9Nksy+3YKzM7FoJoXp7AHG9pGmjP8J3c7iwdwE0V0Mm+ZXaCMLreJuHBsD
cO/P6Sl9qwJdrKAWdB8l15lAeF9+JjKVn5HPh2MOrysReFJglePMqLiT+z9g5Ar9N5C2lEn4abz/
VZOgTfmFYASiXJRd/mXZsTgHGSLIYUGfJ7SKsXCKXJbTGi83fl8t1hxdvgAosq7njw+T+OTPJZEZ
sbICdtJlVSHN+6iRZ+/J6aDyd85A/T1FWujV+ehIFkcYyuHfkrCtxM0DMe3MlVGDbBbfndjv3etA
QjDadfstNykBV6oc72+W7beEoHxC6TUBn0mCF0o3UaLrwTzjdPDIbpmt/SM1+ySkewgG8+Cnn0JX
XX0bgM61yR8Ima6Ez3fYgynNFNDBlbPDlaUkFKoghle/GZHIqFo7DVJxviuE57Jeoqkcaftuw5JC
gw5L8xoTT/EiT3MXyDIF1GyP+lREqk+7l99/QviiqRXJBrZx8AlRM7re/4+bPo+z0/L/OVC73Ufb
mXdBgnx2R8DAp4jJmOlD2XM+Tq3+fin/l/0bzI593OqPfshoSIo+FCspojnYuILsM1DI1tnetpzC
+BufwhukolxhbKeX5uirbvxMgG7wITlHOVv55dR8YNCILzlD8OtKrPnZp3JxVs3/weeR5GL027oO
1jO747T2gqgw5Ndrfzw1+DSeyBzkEq0I98rxdSz7MYkm7n0Hgv+07iJPdRhOh3tV1FBP7OvNdsR+
i0B1jzvMc6WtX9/B+yMHpSGUgZPUPiqlGVFZ/ZjN8sQ3IgQ8ZzyuWLrpL+sHlgiG/uqSqveEvnP6
uDV+fhAw8aKWuwPXwOxEQ5bgKfitnp6qKL8YkFWjCIjRkih4tlPAdIh5Av1lNGO17wh7jrfzVW1y
FDCk8lKFEhne6qc6Yl6mMAb5yfYmkS4qyWb+Aiao4WkckbmZ40x1Lav2v/wXIZ4/j6Z9HwFOM8K4
YpLzMK4tNf3CrcAeqsJ4WQdcZr3UQGpkVN/iU8ESkLnvB5eCjwsJIjFRjmC4/s97fhmH7jBhAoLn
9b79uotDw2ej1U7QBbhHSpNjNvqYd5xZQWGT4ybwWT0ShLG+OswzvB9GLiOUVzGoI4y/zwqnoyHU
eNw0r0UnHWg/awzHaLPGate2dzaRrGCZGMSLKUbnRUI8DZJnY9Fr8wftn1M89mrfC6PW4Ga7DiXW
3AWBGttYkFGag2CdnTPtyByoeDq4FyZy+r+bzNXUqpA/xs/dm4lSKMXXmikumsCs9yqz2Q/MYiEI
X8HainXoflcHjUNPVRkyBeMG+kbgEA/7AXLnNkM0x0jAcdMOntXRSGK+8DfyNvRKMV2jelpjTbYH
0EP1cwZrafoV9aqnKLSHV/Z6qQbYO23e+rKZWsFPAoAeqIjRaxe5n7mKR6CYFjH59o4nOI69zaJ3
C55AABR2nD21WtL7kor7LfVcQLQP8F2p5aetAcLGVi0qmpkpg7lRKBskJeUWr7BknI4c42VYYAW2
D3uKwPXp5sWu9719h1LjTiSGb9ymRepSF3mhqBrHvbC7FtBYNK4t7ktudwpsQ4Wy9cP2c2Ha2Aa0
KSWzKjif58m5sdXAtA6DyD96RKHvulGieTbn8/Z363XQEf7d9FpYf+2epI/Bhg59QgXWfTKI0q8Z
T5JB7z98eZjrqbBqdCdVoazSTSgUUhRCAR9So0v3TjdytQHVw+k1cSzNdRV4fejIh0wbDJUA2w9i
KW9DdGH64/DLsHE8wSLX6HKsgO2BjBp9s7PTkSRYULnx3U7uc24SNMBdrL1u8NPt1LlPWXKKn+w+
v1mh/oN6ef+iKT05PkoKtO3pGK1xnubYAAxZePnA19iM9poF7PuW5msycmvY3XnD37IU3kb37gCX
kzoLdXFcC5ubeiKxjwjmGT04Uf0sw2AkhMO+cITlwmbR1gGqMSXScfXP7MKIy0WAccvVjQG55vep
UAQ/JIBR14lzQO0jEwwpIJ9Hl9gNbVmmw1xmViWRSCt2nYHSxH8TSese4qaUYRXK3qYQqALsiL7n
lq/N+cfynvrGoPXyMO0IIp66o8wxbUWkp3MAm2+fOlqungK2bFfCuJ3dgZ35hSB7ygKbHe0pJsUq
dhxMvJ1pUQUqiob+vLXZoSNLk5D4e2d8KydVfZScrAkwEiCbDv3lWICra+Lm6kZpk5u8o5WbOc6x
9eEYeHRxumBB32219pS6tHT482BTcgJROwrLxBv0T0RoOZFZZ4PZNbB24936MnhomTkrIsaEJXmq
0tFhvGiiIVJV+5OeU4r7YUZPKrFEdycqrxMw+MLLJj5xDyOIvApN7EBt5BdJjDyQj+cmymNYUXGj
rxHD/ijts2QvKy0hhkkWfNnNTJBYbBajrhoOC858Lidz1uqKKlQ8BE2FQmrw6We52BRHMmbrLxRr
LOagLqKIyxBlApVpq/cWqhx4o6RjKhyv0ryTDGbWH5fZAzBGs2cKuhtOsGBz4ga927YZRA1yMmhn
Cem22cNel1UFlW0a5sGYRrx4pAAQSqhA3HNc7meNThYv6KUeQIEwdWGXnsl9xU0kagJQxIpFMi+P
Rf6UsSAB+my4NeT/yEk5HBxwaAhniOn+6XY72PWigzvsPROe+9YlEgZQQ/QCf387fFQ9U2E9IBCb
q0r3L/yT1sU+Z/WKgOKdfqOpyLnShYeM5tpk8oLSuCxilgg+hTMpWSOdcM3SLmBwkBL6wmeuSw2t
8PlejbN8uq3Bi4xw6qqpSG48mPKEhjru+mkI6z/3iNv1KwcCx9l7sHxE058DXe1JSeOWRDigGrRM
4GvH8kRNaa86izpBjtPVcNH9pgUHmMBt5lJdUcFufUutQS5u2FeUlSH2mm38PcDXKQXZUVyEwawt
LF3sM+hvl/rM5htAXK3Ye1WG3iWJ4FlWdtxuy2DAOZ72PNo+VRGw+SeZWiA8YdE1p9LIPsBvfDRy
feOlFpLB/gd6gPTsQRJ5KAJ7QLPUoSpnXrivxj3SjtVSRp86Xv+PbyxqSEC6pozzR1BE0wQtebNF
pmEWbV9yBPJXcta+2mBEz7wm1t8htxvxRb355mCvAGeU3itiYW8hT8DxfTcq8GyzAZZbU0m8u80c
+zmJE1CrYPXu+0uFtMhn3SoMep195ti6PjUjgs3cu3x87fmAGc7b1tvNOjNZhgLcDcJRRm5dCQ7m
hDqU6p1ftsk3KM5F3j+ugRnAACDisYoD+XHmMabKgWLvliEJGaWqnq7dklfSd+WrLVYCZLvprUHv
hNykRDo7T3fn1boYRFELKZJrUdSHnoOXomAF9y+zdUWTT1PnNs/UmYMjs+YWzYSi602wMBst0dcA
LV0rLRyqdJ3/DHoB92nGchFOzfRlRl09Sp2JGExevcVR9izAcbQu+fFfKWB6+gwqGmGvDaqyEY2G
/g88QH04aGNjsHzC4qa/6Kac9dovEa0UwO9mHuB+mzKZEVqu3SUTmxEKq4iMBOIEEZk4Io7I8en7
dawUbSeMWJve6vRax1CgixKCNvUNSB6pele+S3h6F2Uc12GjMYMkP3IEIwNa70xhQ8NKT0RnOXvd
5Cbzz8BLtaRzOIQ9mc+TQ/PDPi484/HztmN0yrb/Qwqx8xCsMiAFHgrKZPczKaTC4yPZCAHdrbcP
thKt1zz5jtqwyF46FQCXVOeUGGganQJAL3aYEIPegAaPK7Pv+/oKAKmR1rZTKFpNnCANfG/iuvUA
qYIObii0MByV7OmKiBTeKVdJitSt3XpH9VuZ6daonoqDwziF/lAfVztKaU0PMpgYMgknYxuLiVqq
eaLoW6Io8Y8KZTSTMlwNGeIojZoGDFt6Mv/lzyEeK/SJZ0hQhBcvz/uKMEDBgI0UHyy8gsKS4oKg
pR89h9xIVMmmGmKboc25d88C4rZ7MBvidaYiPRxYM9zgCXAKUV+p7iRGBUADQkPkbC0+hThaZUIn
2C8PaMrNyRE/OwjWnlNYBLmfgqwAfKHhhpHO9+yo0Nr5Oq4G/Tn62TwfkAefPanVkLg3LkNh1udD
sdI7Zwhb00+DriVjVbok9STJIcpGmuwAJgd/6cSTPgybEUfxmLkjU0C6/DI4XW7Du0tSoLUTJ9xM
Y6DfE2KLokpzAlIN7wI4ajfPHTJPxtXgd8NfJ7dlKcGe+AIQRUq8za9m4JCeOHdQQQ/+F3uQp0a6
KJpmfUIiVrTfX3YyRNxIOmeiKimcgMaZAnh1298g2iCgL51H1x7LwG1w989GQv4K1B/QHrA3WQmT
nqL5YALd89zrF6m9WOpSGDwq4FF7O21UzWLVmaDMIaS02h0R4bl2Ym7OMXYjYrMINFG2lGm/UYpM
pIbOTZSgPAe5d8WvSzox0S5c8pShrmNrk1kUiguh7/kcMKVCoGIVl4xYug4SL5xgx2ze+b8WRtYl
6kdcyssyIata+5lknu6NO/KRuuxF9EHt+H8j/LGI1jZd//ytwx8EOToBCa4Yaz2+o21tubCbPiBV
bFCF2EqZRJwbxzdgnpsJ468FSjiKA9Hwoz1lg7K4fvMaofhtxQklJV3OJx3TRM4Jdfb3lo4pG407
cfgn1TKIt2WLscCbATJ21K69K2uyP2oVUwY/cd6HHBbbCUBMglwBt3AQPuml7CV/ciYXaFACglgO
IVn6NZ/zV6LAzpAoFDBP/DLFauO6WDXP3RPkUIcz1SdOj5DmqIxHUOxolvEK3z71It/SxTFZvUtv
1mJYnlkXcvAuKL2EvoJgCGmEK3X8dbHg5xauD2j+isdHBymW9FMX6374cDQpgsf73iII8JLDLu+N
8Q3ZuRKrMTk59AjJhRRqzSOpHDF3QFmF39xFZsoF5Ro+GO+Tp/3J3YYTS4/xGdiWMbfuky6O+L97
EPRaQPv3zRU3sfdzYi62LP2rljR/m6qm1lCak0TN8ecrvs41YlxewJtD0zstJ3ijRw5Hp2xPhvCM
vzIflsBnWx3Dy7DZ9QmVQYnKtv/Qp0tdAxPdSApgV/qrSLTKO7C79TZ1D/prJt/irwu5WOksnQAc
Ti+CBMrRqM0BBpIGpTKo0XrawigXfc5FlJqmN5/QPyHGlX27wUfDcvvgKUjwLMe2yT75q88UFarK
wpwUsrFoNO74s+2PeHgkiqmcwzT9WJWkwutIpc8xTNcIJAUqKi/UaO2x7a4ximH9CrcQU7M67Jjy
nMkPlKYnXMVs4x3mInaHBDBSOLKAGzINeDIFAW6n0w+6rIMFtwKiAp+Z1a1WKAam91eUFcuQZ5bP
VC//fl+gA2ZqCbDQ/K2rT8oLahFfVQZlAZS2XdabFClP2fo3QNpJEkI0tdRQE+RReKCP2wIFO4IF
0CFeKjcd+oS4kUU3nYFB92gfPKWaxArAxvVwQq4rZXWCvjWYLwT2LilwPaDP6EibB8Qqph3667On
9V4yMW3++SMlmH9WTtCjhS85dzV0cavpmf89U6xXhcpJZ+lkmTnIPeyC/1odiihTGFWi8RNaA9Lr
M6OLB7uEJGcjfAYzEhtTf5vJ88MWgK7Et5O6Ra0EGSnfHxdcQu3Qy067WLqZdCDFRDg7DWcXsUEt
RJdTeu2o/erkS3sFMAs8aaCZu5EFtnJ6TQb7AUHyoBuQ59/YPtJ5vo5+5YOFgMWvWt7bpRdSV+SF
JSw5A6f8mmVcHDOwchWGKtD6aluQeC4DOLfZXA1LIm9eEp2YawoHfQrz6nZhrXRdsMQr22doWLgk
MwdZGGgo9IgarMWB0BZoa5l0ZclV03U01xYXHb/qJg71a3Uc23KZJC7MY/9bmCil8/2Bini+d1ns
ZjkLsGG6DfE9pTqLDPTX9mJK7UwNdiwZ6ze5tGc0IBfkjJlE1WtHcBKHRhbRpdl1VaX6lyyB+Knb
rjyRp5Xvs+7KoKv8ooGdmA1V4siVC/N1mjg+0l3YxyRPDzdgPqdUKTgrRevFygnx9yQMP2ynlASe
2H1fsJPb5GJVnpZOk3QER9A660VzWahJ9+mNVm4mnqNljdFuSsN+3TlgGM8euF0SnCfYBUaUG0jP
Z4R3nP2qZJ6dB835ytuP94ktB8+ms8A7ZH60qktoNpjwgg/o6U+XUzluPA+hbVbwP8kaqNN1JWju
ElkFkA6dHIKzhz6ZXiAhFt74RVh+nDNu0WvaiS+fSf2jZVa/GtFTb/biR7xsYwKEQ8qbIVs48Z3e
UThH+yliDg8Hir/6QeFw0jr89U96he5n6IRhfc9Sa5MGdYDYfzAaAwjuLTiin+rUhNJRSeiJ1Gpl
57AeKihHhEvuA2mS3RPwa1DP4IuBdd74HlL1ZZC9tA/iQbIEGxMEk0hFz7RWgFucbJoZON0jOA3r
26CSUnt5xwk2vqSWndwBAXXPlm2ArWqm317cDYr18PNBpeyZLldv+/AUlRZt3bPMBUsJx39m0I5Z
6G8tO84SB0eda0EG9B3C+0jA6TNKtVcJXlshFuan3XN3t1RS5lOGIeljs3WKzHYCg8wwrnEeGjnW
9SjU4xAo7NqdJ4DqH4Zmfvys9RHzb1Y82kF2QP+fc0/13w9HqN0iYFs9QbK30/b1c3m/KucKOwWO
CN3jxEaMMHE2QYEkseRRd5B/sP4kIYtc4DKjQTHTPXAJwJZJm4Akd8ik0tTnh1Pt1PjNr4/qBijg
0/eoFXFM7s+t2Adj+W/78PIVHUWd5uWnS/53iyNcoQ0f62ZFB74rTvd91rvxgVA64tiSV622dZBc
XyAc1iwJBkXdTdBK2CPH6RnHWj8eYkKfFVY/C1+ITpHZgU4MC8b0VCij4CGrwm9mq8S1cqnIM792
MACobN5A8UkuoD3b5h3O6cVs1LNoyEzOehAWVGd5tzUsB9/hDgWxOBYgxFJ9P0QA5WS6A278PPbe
a/M+osLOBgktBe7Gni3TQ0/Px9yZGgG7ihPW6QgzHN0eW4RyqRx9BJ+8Zy+bQIll/p2hJ+9BX3Bh
OJ624y3pKHe7jVilocAwQXuzyr9EMEEaRCTGePl8vvMJn3PYKZarr1RdKJWEosUsfvSbGmJ3WQuK
G175MRJwr2yvIc+XuvLjzaW3yze9BB8FZ67haYrgZweeMNZAlObQ+KMN4hccrqyd6Yun9lmJbFpb
dFgQfq9YDANF4qD1qi3N1i+UWxRixssD+o8BRlvTpHFV+kQwU99PRhAmiMEM4KFS2tKYgX2uFk24
t4OWwbHv7AxNyS7sEBnYu6EUW+to9DXicxDWMBRFIAlFCJ4e/PDvhFB3VU4dOtFfwHfKM5M3V6hk
4tVgDj+rlAWyX9A4mULVP8rVXaBGS9Ro+BdC/TLq8pJAv652m7zST99Ij70D97TVotLvi0brJ67M
Ihp2vMP3mqbvxWtAgcIpn73SE1JWFTVyMptldwWQt5jcTN7wl1ZHOksuzYFyjnQPNCxXaUD2mhd6
BZMPzhvVBFe4AZSDLBQm0UTqLWR5rpP+gj6PWGNul1mbqwIT7GgBvORVbH3+gdd3rfD96T65plQK
8eE2uCbE22HvIDiY2lnxpw7kv3KtAO6/ZcjL7y/eIK82GqPzOxfsXqw90g9JgkIySsLsn3ZiXbMm
qX8xQ0NKsxDpPCyGLKyQ/bu9OfUWQC9zHfdvuGi15rixOU30SQwg/Sm8BqcpkKF4W5o+kqcZi7Qs
DGDGcg5bnMqQAKTM7vTUFY2VBB5Nrvyn9rsC4bKmnuBDpKpiLAuw+KJyEaUyeNfSk7dmxqQcVVi0
Fgp3V+4boFVcYNkTUnJQUZT6qrHIe9kdL4lrAr9e8rK77naN+Sbb2rinqNwgbA4V9Z0Av7ivqoK9
XKqkJXhdLLsLyKxvd7lGR0ZbMfogDZi+sE7fTTkoeBQoJQ2zbjEFDde1H57j9FsRYPU9srG9OdPs
+dFjjcrtTCkUp/BhemaUO5+Aox5I8gfFf6I0ZEQISk0wBHX4F0l+4gaIRoiBcPpfLhQWHqAZvJRk
ZxRWukZ0DYV9h57vmMIi8woWfwOSmhTcRL7TewK35grCtJ5JKXM3qArYLXgJtXT5tfgWoLd6iKDU
D9j8ggXMBOybfPPGd6IkvuGFkLLwp5kMLBuSa/785P3h+9frEnW/Wk1hVN+7uCGKdXPL0wAanm1X
LWxxLUvRYRh5JTUUR5DciGHhwZJOrwwAUhS6r8MIMYTfMIirAmvM+Kd+jA98nvNYS4n/3IpJPGLG
EXsUg5v5Pws8tu7/Nyf3ltXEOrsY4YYpKiY5Jf1NpksoD3RFh4kL2/19mLX4hknbqcmOL8Db+J84
CTgvuUnBBXN1LJhzcsjq5U4izLoqArXFA3BAvPYWULV4Lrk3E1NxFCvZ4M0YpWIk8Y/04vH7sZRv
1yIcG2iD8qQdAuddfNzcTelOEK1zwjPbJb2xMXGNAFXhjNJ8vNwvXG2JyExE1qtRCe07C4nDCS8N
0Fv9aU2+LxPmzx8jM+Ts7Ow81sSS9aY0MzyNvq3xVGeJHWq0GiyN0Vhbd1SEkeu76ydubBE5KZkZ
HEzy9dEtCnTdzjqAy6PUIMRvVQ8XduizUUaEm7dNJuwHl4a69Osx6NrFovTXQz93yLETKXkxunk6
VDAakCmppjALPJ6g8kIm5e/vAJLSJaG1dV05iprr6B/aNut+IjwdmCnK8OckkL5beytWEsH6LHw/
1I1fAaaf/2upH2YQPSHNdSLjnF/V3No4MUJ1GhQDO22lhPYQ3c0wXtCqoG2L+stu67OEkTYWNSgr
oll5txLOQpVn08wH0ADrQoC8qv//nV0dC7U23kH3EpfXDjBukLxHTevrznBNEbRWgYETzsaLIA6T
mWiFujkK9QofGB+nriwI85KDsEgw8pHzuXtRvGagJV+mZ4euzPvtgN09e/NjIvl05TfsuDlyMDP9
eUP1YjsIkT+7N8V6LuEYPHPICpOIwuojCaOBjTD7cV91qZg48Rg1YNqq5ICj/gJRFUnJihfrQ49p
udaJwWQP3X6wxAQTu2D0gc3R9Q5GIs6sjM0uCvn33t4RCkkk9pAEiKUMk6DHAGtPbJjj+Y/fPU18
zY890eDn/N1+77QJKNtWDT4c9LO0msxrbe1KrmhW+uaMDE4FM6V6rsJNk3CCv3yeu5VohBIXNN+5
PSdAA6pK0H9mKGUJl7y4QXBR/oSPfauTZqNUJODyCBVer6XptSROK6rtzh0v1HzwlSe/4w3DOB3B
BZ6tMmWa0cPT872PbP/IafnFXVq2b5q98/C4xmR6/5kcdRkE+hrSYxMyKOJGAsLQiEMM/pVceAI+
tLQOOyicBBulDL2LnXOAOF1BvcrUoCyjP1pNDUWEfBUIknyTo0LCpjLFBq0Q73DQYQIajCIQzZhQ
YQQuADWCrOcqYfqIb2vxsfxF008DpwU3yoahj+Vs47w/VLahrkZZBp+NciDJn57aUusyJ5UYKBsF
AE73XpoubvIs0U59w6YdHxEBbKp51ylfhh9+gpuFtPDxQK8lCEKIue6cdOOayrgR8omJNeQUP/Gj
qrJa7HZmW8QsL510KmjNYBODxpLAR3FgYL3QusoAaX1NxSSxqkcdmvnL99nzQoYZb3iFhVf9XyWD
VS8VvnBH22d9UzMmcItL6FWSpRwOF2URne7PMJUNsZ0qOGVJhpMRmsCpHRZ5aOtBt7Esmt/utBN2
Pbuluu6woj864nlRKe1RoWYt2RrPkQwvZUKaQ15W1npnaVPE56BXq5T7mB9IE5z6EcGjG2rOxT+T
X5uOm2sIrbzuN5BqH+nd4nV9DPk8bmoyEWQoB9CLQGyTulM4MBUIftZRTvqjY5O/hDRfUSVYUZO5
BTRppfY2kXALG+qH+xyJBV/B/pftSFU2/YGz6XBbaoLmyzHt6dzla9OPdOaPYI7aT2lxlsY11MbW
NlIqA8zMrpSymInAcQEwc9jW3MbNI0o/wcJXhWiknaNCQlq8A0KHUw4gmOUvzL/DL84qekKglsph
nj/+gcIb8ggEWpmi9sAOd9diN5AfLaUK2pwRwOEasK66GawE758111j/ltQqWnxl7Fl62MOc3Wyi
IIK1Y9zrjXOEt+iwLTnybib7LbF8ooGcVI4ecZ2bYEVrXil4CLaFCxZvnhNcUWkbgh5SULCnn//h
oNE2cD1hVC53cURrCisn+PC2nS4u9xDESJCm/Xtcpky4UHdIX4BIHGZRz7dejH7ByDYFWajrU/Wb
qO+LsSsEAVmhIgeiGytIHhv8sIVsdXfFe5TfuHQSIh2AFtRltxzdCZf0kR3AIF3RrMkhKBQylio7
m/khFGH5NQjhucj7tGEsowoDAtksiRycGvuOnYASwwvjbpckgzCUZ7LV4c7TxVIeuogHd1xZQMy0
9BDfcMaWqzX2QEAAkswTjCprNk/IxGres1dCd6nmWUe7xFjEnV3r0zAQZJl+oO6Arz0Vi5M00oun
jH0WWPeb3EydoC/vIm6AOWUsP+zV4Eo4nkFwdGZ0F/ro2bvckcR6JZSso1GQPR3zXwhJ53HTOT0r
HSG3ye8QgetLuvc0ZoywYMzci6oXBbq6odQzyrgcxZCnMX4o1lK56fAapoBijcEi/wv60UToGDtB
Ll8OCdHLv+3bnxmwSWwpM0qtC6/hTXrn4R5K+hMuNSkXWT/o5XL4KZ+rY3U9rJOKJF6ZJgqDsB3s
OlUGBpkZmy8umcXOYVubu/JsdjI4D/KKYKWYPVDuGC8IirsUlipjfD9atcgRZWPh2xchr1O5byro
3Fs2nU7v2Y2NxBGVRHL4vVOAGjMig0xfmSfe8IdmIwO97RG7EmWx3Wjmlr0JmYN9/TZt6xxAL2St
KoLjk7RSLdxGBS9KWDpN+IrUD24xfTpfus+85f72XANYo9RcDoiOQNjAO6NlI11cb9TFF6fCiT+W
uqkNpApxRVyelL+mdnhlCH3keKWmwbJKAyoeB9joKygYEv1C4f38Cz7XIk+Vx5Hs8QqL5wLUNex9
SKVRZKUp6yqc24CjXmJFnqq4fxPBOz/3QmDcYXbRL5qbor/7dRcXZAUVj3HnOHpGk2lLRof0Dqrm
/RdwXIenVf3K/8uSqQU1XqiPDY7Ufvpol9bzZZ+KEQDLbYgeZeq62FQT3a8+32wCm9U618EAV9TQ
iYCsGjzxKGihrqMCV9zzk4PcE708wTsRcYZRZvLn1avsdmxTInUmslgHW0kRoKJN0PI4LHySoF5v
0vJ21hErwD8gp/fJce7OxmzmHP+lNqdprHJy6jQJTJXcGF9ywPJm7fX55vL4+7Y9tnAGQMpahRFd
TplveI3jCoBRgWvOgLB+WAvub0jZEEYdGoLOTf4hdltaHVDRwcdkHHAdm2TSU3JyZ45zptZdREUz
vCdRvEGc++mlkK0bAFb/CecApS0fun5bkn0eH8nfUZcrul2pKEl8TKWSCJpWf7Zmm0T7h1pS0adQ
whXLG8G/24hxaUtG8ABGMVqCGYrGH4cIYiD6ccXC4SRM5mI+7s2G3hW8y60o1Fu45bmYntRv5wD6
NicyTeIKgQCJ9FV3SP67erqU0NxBFo0uOcDwanFYnMp5wOV/WIlHiioThNFhf89M/jFCuL/u/Qwr
jujCtXgf5BMoW82afA6u3tUT9D1shypnQVzmKr6YIXhNHuWzNxRtpNWIIPy+BWPsMNfnz4xCx+9P
tBL9r3Nh9IzAZyVOBoNVuHDlXSvX5R+JQ/z8dpx4/tFs5sfEji4w/a9LcglfH1ektrPYfbvyvps7
RmE/vrtr7VoE/sFzJAS8kNva4jfml0aMokTcFWcZTWLh5Sr70+yKzjklx1qtDYYgM49wCU+9jb1G
VLN9c1Oe5XrwhDsnaXkKlIftXjjGyAQFe/oiMYqVaCUktS7ffmSjPTrEHoBrCUwk4aWEkdAfJR6D
w9PpXCEV3O+sXQJF370FurFteiQcleF92EGFR31JBt4SmvmoQflr0XMovLfSyac51HWo7jOGZVjb
tTRFyloHBejtm3y3nWSMCS3dW9LUkJXVtxtof0J7ywN3KQtctbxu11d2E881xk54DWc7GwRAmM55
RmMSTEmTJE6SqgpeGngbT0SMiUuwqpkT7wh7GeCStVP8ZML6crAnVJYLKy+aAJ+Ad7UZpsuXOKyV
21Z/hkREdvCLCBW4l27Xm/9RYT7FiIYM29aZn6iJ3S8x9tOGK63D6pWy0OanS8xgYrkhpAPVi07s
Ix/UlzJlj+lYUGUZd9yqkg0EKUPEuvIlaps6tjntsCjrnzpnocNtA1kP5+b8eOaWUaQ5FXsc5tWc
KXndpEfaqy7gCy6O9f8o9e4/FYiqL1Ji4mlPUghvRZSK/8uWms0+jlVY6JztTXWoo/yZ+QppUWtc
E/phmzeQDk32UrZ7WQsJ3luHaOykohcQvvuZsKmaBWjzVReP2c1B+Vbh7+1OnE4wza4IAl0bUHr2
CJbh6fIe63FjtX9XYUolJszQT6AO+nOrvGNZaWERxq4KLH6U5z8RZlLrUm1JHUceadv8cCLEpLRB
WoDC2GcloYSpKBuOyeQAFTl2WF6ARpd1AWwryhbNMFZ4OHgwJ6I8eQvo7wNt0N0a7UFRpU/ug96z
h17G4a8VeLAuGGyqjiHqk52UCYfIBqYdvquM0rXtkZnCSdH4BfE5xpwZ4f8NO4MvtTES5/cLu04w
IWSq50lIFvcCUmSAP0CLJJJuC3bKnVf+Ha6qs4Hq7NVGgzGzs0UjngzWGkkLhH4wJYyC7neN8ZFn
V9Tsq0d/ap5j8aWL/gEuyPtrroPjLlI/fWSQkzsGts2IAHxE4ME1UDJ77rf1M+22cRs7mrSWOifq
CJ8EYRe7F0DduVhOlTO3HzMLsdO/kTcyBxlMman7VW2KMNyaPIDqfahHO4SwekOjg7qfs6WHxzpT
uzlZQ5VJ+a5ga0VoiJMP3fHXeFcaaB6L/CEa3MBkbavYOzGdxmjiITlSSTP5zYMjDLTDmWF0Jxqm
hYbUMb/07VmdC9agP8NopNfWHzRGXlSqa9Wi+GCudTJlFgbkU/9DKVZ2Lr+sN0d1ZAqhtD/JjqMr
egQbSEF/3eAoTViS5BwQ9L7Wm218VeI6PlW8Q/ESn//3JVVEGl0CngD+30iedDFEKAzxZcuaEJBt
7JPIeczzHTNZmLk7+FrqaHpKGDSxheHTvXvKPUXvMZAb4KPiy7lAD4RQTdygyLUtqWdMImjjbYj5
v7GpvDtUx8tzN5HjXt2jwCkOLzInQPWwJ739RSrwm0ApdHFEa15hL8mtLJKvo5nEjpkPBt8WwAzq
4MLI20bHQnuYu567v12iokT/EhZrcDLp731HcgpUVBf0Ym3m2Nddx9ADFs2FIDN3pYlzq1Khj9Ej
m+wGG/a+iqBKY1WoaQzx9riqCXhaQy9xTFg8AuHqO+U47PPGKBaRE9BxYoHdBY8wgW6a+n7FYCuY
jWlVZPthAuyaGzjioMXwUuFV6sKCOvUzZZHQ9QYniJyELHFIThTbpPEnX8UjXO6o8qDeTLePgWqV
zoIAWZoTHrdj8XqzAiSFOgSzZW3f0XyUmMPJoqMbRw4UzDGkekKFpf7+jDH+AXjUu3XDXv+C1Re2
rjXryCQETpN8OuoTPLx5HWl4AqWvEQPsuLCTN8YG+Lz/GCz1Y6UULMSXQxsRg5db9YHvjeDfC4GF
E7yE242InR1/Ex06cB9pQbNYF5G1/F+BrELoSJAVvgWnfFHKXLZ3X6JOoRVM1oxfPGJ/wCVDHMa1
8j1J67K7iBdVMk/KKv0V9XhoTyf334a6eLMR7vNGwTajbIgz4n7z7Q3I8kF6ynQBUMqMii5Rs+/l
tXnTu3T+YzCTLiHZudLhLs+hcl6Q93//OVLScRslVm+AlI+FHjDK2p1H1sihhrzV/q1i+EtQvF+n
NJ/egFayHFV9IbcWXuOxkH1O2QRtqfdy7uzOpmOWI5GiD+4iwA6R5s7kbjCrv1JbhbFhwdiuStPE
KC7xGUN+Jb1aOdN2M9FZrIhEPTMYyb/VpAxqFsqmgKkQegT469eJnSu8YBqZ7WX0cGahfVhphImw
08MbNpNYzo7sgdqikwYo/zwfrSNqHbj1wKMfuNe9/nyXniDoToXkzmNI4BGArYZcGBYK+vyiKAws
PQJ7jI5pN5uAhLDs/xpLObJWbC5+IbYXiaJScuFlfZOtrPP1mSQkGoHheJGhG+vn+Pv9cxRqNKMY
B9nykY8eCpbusJvU3PHUH8xesmzy/Godzl9ER85D3BlAOzYiyZa8pJLfAax5qLtUdb6KwSrZoBdO
FMidLofkrNn52m9nuAbTiGRO+qBkbnHdrT/GY/fs3DTscFAOgq04wScB8hAd3tLnpZl9YQ70X5nm
L8QYz8IlcxxG4ZaqZ9n8vUxlMWJVO4ZiBnmVphSBQcMxTLFQleU/wYFkF2ZTUhnh1IWakr0MltpO
R9ALxHa5ATwi4T5B/NL/iNgcvbcioRxbwCJOyZQcqg7i6qHecMr0WOFX+cLd+jmOmR8pydC26+/I
/jEUGDoqua/ww9lPQR5HqYl25WPTfDs/1v6o7JOLLaF2yf86ZM9ChItYmHzK2GybgN9PiACf8T4S
usSH9gpuvWjYJLFUy+QBPVkgZxsszTMDsaQ5w8M98obPD7DYf6dHofTyvMqZvRZcASv48nF/UZyk
OiG+FzSsKJ1ggW+vgx6TMvqBoaZg0OWTnRpeqsD13PINcqKVV0jwgVpuzI5CqTRvhsP/cx14Fs7F
pTVgRcse1IpeUgGjwVi/bdtW4wzAKg/iML8VSr1pSX/gRLZByPHZfoUJ30je3K2DxbBPaAjAauAH
BSnyGEIAg3+Xgl4auQKaRj90gJ/slQrDvE1PezyPv3Sprf72n5zBFcCRPDSZFdjm5JAbtpcsW3qt
dFcCffa2Tc/siSTpXB/kbcfHqx8aQzU+sLR8TJaDY5Phdy9gef0ltCcz7yREegDbDJfYXEXqHSL9
O9AXHCkbLjphbh4ZRJK5l/zp2NBaEVpOPLJDaQ+Gpx+wNoNCW88pTU+N7F2iKlZAYYDMU5bFL3Q+
VSVLXgT2bcfaOPrkSF5X1Ff1Q0Us/wCB0MkQiFemM8g9uaxyXMRGBtmX7xDP3ySr0BoKrhORry5Z
jXNIUaxlxVRuA+ziyi/UBk+Hc2ORM4q+XDyRxoQmOhlihLaGW9ljtwU5TfR5wOVf4Z32zavebPEc
mTWkqWW7d96HvNhOnoWZ+UorcSpMuG89UvhAb4tuPeVaELkrNiaT3RPnwR6xWwd0herS7AyNLmUv
aX7bYKq/5FGW7VHPFc8tqIw9+neCAGjG/SGEBn0Tve3Qq0LGEFEj50BTaoQIZQtobsnvd+A+etOm
XWYZL2DOv1hzIy9Jtpb8aU1lJg13NOJfyhUfDtBGPLD6QVAlc61Bg7z/NHMxzxwVaC+yY9ULx8Hc
PkZ5XEc3HsHGtzpKzs+W3pwzY6saEZ2rR2NrKw7HkH5FBR8lIwE2C9eCiDzsG6GM2XBeRV/yh0Tz
kwm11D4ka65SlZRhogJb+PnOgx+nOUruXzA7sP2X5gILfWIIUmer0fLm8wqs6+airqJsFHjirlxo
hrZw/O+pLbYevCJlKLER94GjOxv27AyaIVhmgfkz102Mn8a4y8MCNRbO9AmFM66TpwkGqU08hS/J
V/i+q1UlXRc0Sqr2cpYYX+f7/4Kawit8I5FMeCGADP/06YddEBq85rfK+E/J1Kv3OEt2LataQQRP
mfhacpMM7BNChBIjs1cznKdP8Ptt75tJgmQQSV1vyPG7CrSS7Nv1rPFZULgzcr8BLCtEnh0ykjI9
xesiOiicvDkc/alfSTHp0dKkT01p380aryjYUOs7rMbVps9qHjLHsj1TvTIX50/MCa4R6qmjP6XZ
gc0HUgxzCCtybJuXbdhxFvynM+Owg3sRbRx0Y/uuJXkg1824W7WQYaOwNITxoMFcpePwIODXu1Ix
a3PkC2LEHVp7AR54c0nvGDPcNMA4ZkYe+X+fWi6/gXx3RndVPTk46j7XSkORvpsiGhEb3zP3Ew7d
ZhiLYZpvwETMIQYqxOLI/x5syfJeA/zEx+z9k3miXE4XSaWVhdMmc4ik8Zdid8+WJotr3+nq46VH
ggpJ6DlvnMsMauTcvQDj+26c/gg1QZVy/DP3bFYC8KYmmWRT2C/oKFvji7XOdY5mNUgl40vbfbMl
GLfzib1Y9a2C2V/tdsxZTq2djku38jG3zhdDJthKi6Ig0S3I/AZJb8Ra/JXt4AaRKjL5Z/yg3dQe
77fcscXuBZGD5Y7tjFAe+RwB2f1waCAbHD+PE5qWEYThLkKyP362EIVwi372O4YQ/xPyo3RIYE9I
0/qvZ5hDgm5jGepC1UeFXpRLETOxv986cjirQdvUboGZmW1wt7uglWuRKQPpVhyveTJSWyFUQz1k
bAHgb1CiCU61VwzvbUUEatoLjSviW5C+6bVXFCi2JQCxIo1NthMfrg4b/6RhUc73BpeCzV1bIHrG
y0AftOIHYr2Eczuz7kzK27BprPtmqgbtyFrSOJekVlH3z9cqS4PuCwb2m7ejqFOs5qVT6YGIEAyj
HfBCtr7rZcw1s8XgYp0K331SwznAm29uuLqKl1x+8ohrmbsOfPmKYu34EwzHmfP3LILQVJRwMfEj
Mu30TPZ+kP5h6q8mptA/JjoSTIWETzMDWd3nOgjOAH3hGzzp3LhhiNAKkDkQzFHMpPPklJ8n9cYA
pAmtMWTCkAjIFjK47L5KE+B20URCOms0kAO3o5Fv5/FOr4pcOudT5wXZJHXcYORm0Qx/gyidzOjA
9VWnwnvIerGHe9TbSQvtk70ZvVv920RbVsmGwsxCCsdxxNz2CCsl015FKjf6GuAt1mw9DLgpmZiZ
GhVkp2hWtAekb8RMyc0xakOflETJ2lo28sauGDi087ecoS6N0NvZqxL3khJGytFsTNVnr6XFWLRj
mld9s8LGyqmwfDOQX58pBhbO9jgI9yds5u4ckB9sCqFhThzmE/qEsYdnMZYYZ3DzDUrOFluq/q2+
bMBHj+Rc4FGZ997JtrykLaMbCvnpX+VzJqsXwPDtRVX0oTdJpZo+ppm/69/AG3gDrO9cDGFN2sWT
QBhCwt+C85Rdg0Bd/8d/PmI2Wer+ml+FAaRttMS7CsVDKNESN8D86IOQCUh6ENb45xLhdXcd7Xs4
ECVGRE6eEQq+edJJOagHif+ECTihorYy492+dmkOzMqLGCDy0hVjtVFDYghGAOmP/F3F2V/M0JFG
Vk1lSEUOR4tWxEDeFpSEoSEEkkHnC2LWuPEgEmKunE9OPKCH7T2F79iMYRnpKBe75/3pPZfynus7
1Rm8fd5Q9DagAOLxm0mDqu/0wNnZBc0vxnmXi5yhOP0twVfMw3eSmB+5wbRPnJ+2B+6HLqZ+RFn6
w0KsBA2RNXOrIM33ZsVELB0wwo02aywv3Ny77uOFDYQSoCkO8R9eFGwrzjn6gI3Nvq5b9HP/njnx
mW6/xfCAKctvctr/b74VlGXnHrMv946EyB6IjLSV96fRkifJHAuKqQU5p33Wxcl98kTd8t17IcVA
h9L27p5ZY8ix666CqA4hzbiZEDqhWZg4PCD9v+InZbKdeI8Av4Zxu3YFBzJUTqhvLnfNnJ9ie/uu
izbNoLcP6B8EDgP3oonL077iFr/fdOvRzkKQ+ka3PTec9biWKIAjo6Ud4XLos3CPVJxWL2NtT8R5
QrJfxwX9/RnlsbYsq5Y5CjkOMNThYeFTxovVZDtv4YdfEOdVK8dnO7QEWapZKuGGn4WNK2xYEAmw
oMwj9SpyCjSjJqHT7jP74tFlVDFM7cjaTu0tsOVbsVLTKwboFRMYaGJnMTsuwnndy8n+4QmwuC6a
8oyvWmSNAQ5yZ4w8nELlUurwkLvHYw4igleWPlPySHkuuD3N7ejv4U7lUw7jmXVkfgWMJNZB/zp2
HzvAYB2N0GbjLqqH2Ceyk9xuh5TMa7Rvh34Wlv6FlFN55oUV4yjDVDLzfCjAIiYIhUeLCjhYxhkp
3Nz0wodxwQutlIklpxeYOH6eOVKbfnYegltPwWITjedp+5VwtM3uuDdl3790Z+/8Rst37rbZz/gH
B0eM4/wTsAfM/gyz7EyiLACpAbYBqr1/v1Z0Q0AlgBUpBMJwvvQfW378uiSHmS2RGmRP/OiMb25O
ChnLS0OnKUnZFtVb75wZdls9wZNKIUMyoZDNX8jIm0dOw5+QZZNKeq1Xo6XeD1T5hyCwqHFGi5mv
75XSceGtPI3XMRm7gZMPzBJ9GyGDr9R05D1sY6X/rAu1y782WGleDXWNDnA36/3WH1n8A4d3eoQt
dS9QQq0BG4jf6MuUqVfvsA2R494QqsHL+H7Qn0IaBs3ioHRAQrRNQBrqWYqnvJFoRBf7TElKfm7L
yn1rv8ucLs8MW5I4zcH5Cj2Jl8jj1gj6PyaTb4B0Z2G4P9I/3380wPsCrQdtqnT+8yGEhX75yAtG
D2zoVXDBKkwwYqB7fh4qG/myaJG+TRwEkdbX6cxoMzsrZkJwlwt6vxARDTxccV2IOtxT1Uce0zoS
CkM9VVC6vc5uQy2Nt3jK3+Ak/7yA6zRlula9PKn9jTfNRuOgNT6JpzpStlPMgYDnwiHvowSlxzj6
+Qt528xebB0fGldg5v7YjiobsCEMzoI7lvPjM/2kK7iGW87+Bfn37YX1bpVHq2S7IkqoUnRu2ez9
JU2IzbJze9evvJrz1S+NepAkPAB5opy/UEOzYnGD6oAfLZe57Dtrd8uvQd5HxB7fiM9LYXMRdOVX
yIrKdWtidR045KqxxmnBeu9fCai0QVBZXuCpV3Pd+VnDxGl5fNk7NydX8y0DG5Ft6v8+9yOMnTrD
o5fqxJqVG9CcB5mD/I2xxcVstnC8HxoKVNsuWTOouNK25jKWtuUo+9MiRXB1oluOcJN/pYA4AcvT
rh6v7mRN9TI0MrQKZ6TzlB7Juw3UMhNnDHIDgSMmdGDxXV/RYpd8BamtXZ4e6XwcNV2NKIlS5PGQ
aA4w1zc/Xg1S0b4tTEKRXQe7eBFF4rCZDrYt6sCwtE8THUmI9YpWnDRN09X8TodDCaC9+P1D4qa/
g6puSCLqq4wJ1JXTUgO2pQDMMswqNbejrbl20zEaFM1fBVpH+58uxFackTO2pWI93diOYdGdPVtJ
xkuzzVTg346LbAVFKKya8s18xqSzxVspH9WYpJlMhu17zumAM1ETFjy4SH2XhCeX2mu2Ig+tdDvX
4tlSalCOaK+/QX9Uus1aTBoYM4LW6y1TloTcU3PQsJzBbpPGIeqmByKWwELSY2+GzzFdrPv20zZ3
Vm/0rmx1VjU3wvl55xgENhUdFJsl/hcToIRMGhZkatS434yQDzTUmSaNgzra4AhU1bOVk9kUbk2g
cQgB3/8IC4AmklO4FXDDIzR3RcThF3GoDV6Rj3nt1nO0XKnfK6Xl2Pck46YmZ8yZbwNhbqSLRLT9
JDF673cf+iwtmJ4O/HofFKqEFxoB5XmfCuUBO+v45GLUmJEA0OE20ZDJAxIH69/u6QHR1EDMwcGK
0r2Zb6J8L3XzmDyO6g08WSseNIzCC3XG2FdJbAejTjVuIY7mIvtZJvMhxXU7yfPdsekynmM/SNiH
1JbAQYKBp5oURjF2qZwL2oKbqSfHwDTrkSQ7MbvFNA1YzS5hKaRRdkZNdSXr2etOn/NIswMjRLT6
KLfwcRwSy56EP4L8yaVb8vblN2BqNBkxlqeRt7E1eQebToPaFo52mRTmxgMttJcs5ZEv32GZvufk
T3xUdGVqsPpyhQTcRAF1FWws/Ox80f58oCDSSgL6odBp2tfjwuHAFCd1YRVK/D6sFC+uht2bBI0v
hCllKBBRERNKRlcpIQ0iHPmzs/CbSshgoOcN7doXD1ALZbe8J9USGsi8ZPacCtCpgbC6jhq9rIYA
dZFwMhXNtTfK5y0Z/sz2gBbf2szqTXK/mt7EaoQPa2nIp0B8Lm+tqbUx7hyGpe1F9EwyVWValiOG
DFyLaRjKTrBLdt2Asjv/dAGEOXMxsl43pET0h/4D93CBURUMqUCreJDqeeCZ/nf2/CHA5sx41qZT
NvMjC45+s5OtIyohcTx3Yc5elo0pfDtR7hFyBOgEhzd008jZRyJbMUl+TqDjZZOspQwtd1v/5qqq
cQ/q8Fe++NQxdrF9/1wMWKREKEW6KB2aFucOKGh1NUExa2Xg3ekLMIii5m7apuZVxw1H7h1rjnDQ
tDJ7mrFJiUNu+61Om2xX/Nr6+ZzrV2Vn0K4LVlpda1hShitG3PYrdjExvxvtOeQcZ/5B+7aTbdu7
C1v+yjsb1l2TXak91yBALgVFxewjwyiwHkI7Ydly6zQVvZ54uBZQ+oCZA3VBsCxXFd5UpZdSvuwo
SkGeFcrRQ4HB0Z2Wlgf9NEm9RzMyG+fG71p+3ukDtzOR3lOkX6rUFaiBhk6Rj37ptOTxzH+PPm7M
ZHdAlnOqBQuCRZuGAcY3JJwIGUCQcPzSH+dmH73Ge+lCtWEfPVBBIBMSaxwZXb2CcROoIW3DyrEg
s2dMBUHFXfgp1AF0vi9OWcwgLJvRUZTSLvBDPASspBNyxc6jNyDaKVFV8VhWMuMNi+6KmXpOWDjm
zsQpH8dQBjf6dg1SJPcjmhkhTQ2h4HYfhOam3gAdRNVFxqqdLlOBccimoXJTjNXDJOnVcnSDNCI1
TksZB9enLRlF9QYcD0BCXoaOmLidDaQ+CR+Kze4xJ6hbPMbr/DT2Fhtn83zzyIsWUBBew0X9Ge03
+RgLCknoxD3SqypnFakCy2NkXLeDLe6PSy5cNmyGTeYDYSNfuq1DI5oBzzYm0g5ASfzD5Es7/3dz
tzHA15IV/U1oai30I7bDO4HbefjC7/3uRupN4pW1fbxIPlHIk/mWZXXfeApndb7tR/aYTVPqIdEG
9Il0WeZEsg9LOaBsjNGuxZn2V7VjX1o6uH91ouiC46YMmE7wZdX/hkffx2T5QgVRtmlDL12/RPLY
gyR2xVRYnjuqYYjIeydWea4s2aTschDdbvbF0J8w5zZx+wb1uCDtFLX3fQeiV1N9ahDJ8jzuDxZB
/5wWB/5ICTTL6Gu6WQRm6yjVo0+CgPytzpKT5DRZ8whjDyTzvCD09PRqS/TtswzlO4chKsniZ9lF
06MF48Oxgs6DnntERrQtyAutdZ7nAiMOkAdpRUB5H2OBwB7NYCKcmLHHnMbEbRT7KVmzOu7zYWdB
kUyfhmpUaU0i7FgSbB0UjIIPWLDVe9kMiAMwZimPdVDxckTiNltVvmPiVuNnOA3yEOSGJA5nUUI4
cjQrC8/HqXhxAb1qm1z+NihWzRi361ddaXRVc3IRrkY24K0TVDPDRlZdcUCArKP9a8G18UmdO7qN
bnGQhCFSpTo7i4RAo1V7zvRvQF66DgpBiUpPmHPNxnRGoVp7KZh7AHE9nqytTY9LqLzFLFbKzLwW
J/HjzxFFyXBH0AKsxWDzSLTOAPVMatH014W/+OLkLZqGT2CfWrdBuIYgEjhPQokkgeGhqNuWVFKH
6X6SPbXMbUaAX/T30Ot4VD/X1lAJwpzSAsZQos9z7mkuvbsGu/D+XRzypzUF6oH/KGW9vdG4ukq3
LxgRQ8/BVMrUYKVws1rYRJ5LvdIKFKVgg+BmdyIZcNRgro4YXNdAEwiVvNx4UFLmb300rHth6QZS
cUQT6aoQ+rT31wquN6dUopyP42+1vMBVm6XqknwGcMKmlh46WQBs92PxC2mlMrDJLAWDghHRFXEy
yGJZ5E+cI4y6Gy00jHVpCtBEoX5p3hVWHXDdlWrEn1ujeZSTnTFz4Ngq9HWsJL+ci3359DJRORCJ
kWBSx69QCDYxp+khmOTjKOGqHDoRm7acEECp4nVSJgdhL7/SY1HfSTDyJY2TSatUrX9aDnnvSSBN
8c8h1mggofp5CGfxCQ7Va20Nt0rmuIB+hKP0ZKzIFwBBxoSB1haRkcsJVkYm8Ts8RqsFOqbv8qT7
J64Nt/HkJJ1mdZUd9bLdJiGdvWje8ygY2gbP/9QWj6CfpSvJBtN4iRBt47epTXpzIOfHNykueNFW
5grofBG7s0hz+yrKpE6gjteELQ94UcQHrGHGYY92yVhl515sPmigU0mM1kYepZpPgZBSAVAVALWl
khvIeMM+PdehiBWk3NRFXuRZE0krH/COwzd86rprjZsB7d2Uj3WI+LYu6840RGckpDVYo3Lrl+8r
YSZtuc+1XduijzoNJ0OFEV3p/eufeWRGzGaEptusAZuwpVA05sJznGSUY+CTUpm4PWhUL+gluQy+
Ov11a7LnkDLmM7RKHrNn2RUb4oTnJJX3neAYcQ0Qi3KjaQTEIHc0GGmxsqC0LUIhxZ3kV+pOTS8C
uC8GsYww4D3xrNvnCOTYHrUxM7QGxmZ6puibyPGmRgckKdVr490Mekq9IuJAqqa/u7sFzCL/n7Uz
i+JwpFPpNiifHO3WG+GtWZwUmslhNe9lLAem2UQdiwVp8JBWvNPG3r7Ursr7mEAPdDp57J0cgxGW
rRfhyyZtpdSbXPyN0WnmFmaHqAeZtXdSUygyS92ux55K9vRLjJFtlAh/Qo9+IJ6sPQ0ovH1DcaEg
EJ9/RXXhbXH4lZ0x5v/tME4pF4g5Z53CZHFluyMdfcleKvXYZWWUXsHyiK7FLZiq9PkYfSAzPesU
UlRydth+GjLEbhnf3TOwA0mHIGhf2Ut3B+u6hcL3TyYfTi8phuPINOq3wSXg71uwPm896q2N8qkw
RdPXhhrE1l1kLf5otKmZmsGRysFU3QPofJ0w00PVcIdQ3y4Ed6A5CpzVq8qjbhQQVS4QcutMvxhl
AwS2eDM+xWmAkIJ8NKX/me+wwoxqGZ0P1C1cbLxyPCrDbWnh2o8RXcjX2Qs6PoRp8/kxp8PpQuEr
CX9C4BU7NDen3r4zqycpJvJ0alhAzH4tQ1R81DsYeyQN0egdj/maCZ3yzVomKEkVH7qeSLtErxw1
VXXIKZe3crrnxIHb+aii0Tdf67GwZLbny7IzfFGCpIdfNbpSa66ctQNkNXfOLYOogy27++qiCyJm
KGQbavRUg0sufuPyDYyiHd50ndm9OcKZwPjvp6Cm48hL5SJEUuHEjGrTfHVvZStzjPj14rBL5l9B
IFGdOK4E4QNJe9+KmLALmJDbi7XaQaidcdt2nFMbJh4ZvHLCtSuF5KmRo1h9kf1PuN5XcmcgeWg7
KB0qc+w10oHODtQHVKDpWR1UngzJ2tA0LVgQbWlu/dBNdbKUW8ICKaafiDuE7REswPqebWGrbk0k
UZyWgnimx8w99f5YSmdfQrtgjXXvjcuevdB8K5iRFP3moYM6rfpOE7moaSTH746VMl8lYHeNEjcd
2M1KWYQ2up61e7W2nr97W4JCOXzXUgFIjqE5qZWwQQoUt4SDHoVgKYnFVXc4QIKXZg43O2z8XbPH
Hw3BdpH43EvVuAZusI4bhntzG8BwOk0zRTFqGnuzueTI0uY7mVkNvDujUT+9+97svZ28Gdoc7iz5
nC7uagXgisPsZLoEQV75Dtt5eJlgV++Jk1r1F0ADUBdoMFEcmLtqp6xrZ4ye2oiu55vnu6z8DYzB
N1xJXqoL+Bo+SDdBdh4xyEZaFc7FdQGVGeH6ZfK61StyFldDmknHPfpzqZIclInQ1sD/4/KX6mUB
pej+GPh++mhrdGDOAwopZ8CzJ00p5TodycugloIKTH6ZK2jdgEBiVztXbaWBMkkmhmhWgjmDDFRB
IwGsCMe1FuWYDujQsibxSwLkAA0Z/V8VayiwwEtcrcG49RLLeiOLUGep6SGqsnYFpXcrhB9sDoVJ
tL7228o3wdwie2ZRlsclG/7ZHPM3RySIV4jtB4GrGt8h7yt6scdMn2HTfYSu9ZUPMzdS0NuGnHgm
Oz6hkgnbu2CQVeO7BfN7rTLN5EWu8YHVYU1iFehQsln6K45ks9FU4wN7YT+SCTDij8xMWPDpjtRG
9qAeQt6D/q7MLSLjqf5+CkLHULmKQNMsKVkF4OCFzsfHraVtZPJwCBABQ3uPd8Q4WWEAh3RAXHTD
he62Ako+ekWCsZ+9EUJZUFDDxmhECcq+9BjriJvi8qok+4uoU2ApIlavCA+Lk7UOylxRRfjB2rqO
852IhJxT732oUAdDWwYQYEAGiUO+wn3cPGR/LP3X4M8IMLcQG4BtPh260ZVNdkKq+/ibSN3YKweg
eqhXqHilglGFlmeFjJs8HbZHt/XUMmvDoE0S1Zc/+sJd0DfOn1ZxIUvH7s0nAoO3UmWRmirDjpVW
WjjXvkM/8isHzaMSjrpEmtjeO5TXgNqSSMP0NE/VwE/TQ10TANxzjfCePAML8WsENGKwpC3NaGLV
j3coT494jl5I7pWalv0Y+D354LuSi7dX64PJ2Flp6kUzmpWwqs7HSXS3FtRO+qTDfGxH157/DH1q
ce7mqYfVFE2Mvrry7PVLIlcG8Q6nIwl/Bcoi6PYnyZIYxAy7pD+1LQhVCnTElFxUDem+uhGUiw7H
M//2BHUju7I+A61p63YlCu6z22iQ2gZ6D8vNlRWQbAU+SlDchjhOyuGN25tfL84wOU3hbh+FwwjP
Av4nCQ0AijbG580tGmQvHXE41ElFdY9HIo+Y+JrQn/gstp33FG/iqzteOPaRMgtRrHlyv31AvaLl
SaCnmoFNP9ip3gaux64Z7zftAE5FHYISQvtIZlg4lk7nDeFMxNUeZ/JozZpwX7oMkC6vN7myON1+
NY9i2lCgn/WZofJM6SCs2upNi8h5WgGCcha8eeHtV02kilckGeewkp0Ykg0M6SpLfSv3qxiuxjre
HtkljmECtgF27m1rj6GNkc8lQXsUWhgCNavSRNx6KC1vCF9ntXrTrL17LrIQKsXb/ymB3w8Ga7HO
pQCeF15oR9z60aesWBmIk/Sr/dQbShTJADKjuwBwMPqmCNOLiDeEzHr5NcmqwmoWpF+jX0pcQbw5
HJCosK5AcY6RMi8aJkiRw6iyXy9VJmRIi3Fv59SZbu3UryG3hU9HFEtW1rt5z6e7jwfyV+8UJFac
mbf5gc2zOcwvqzQalFpufQfxnIg7dm0Hel8bAUVhhyFlOCEHJNZNrXXxubjMjpwNdrHbIpqi1og1
UsWN0gg+P5IdolcDJf45YMJIaXSYkc0JQGQBa6snuxvIq73LAqX0/4veNSw6FsBBWwwKUiSLNnZW
8cHA+tDiwVKLEWFbAv+NEcVV55utfM0FZ8OJEhMB3AToBcpYY4AnEAddFqYs0U1B2YPkf1jlyxN7
znBfVwZRa1XOZjxvJ+NndAFJrRqaHrKymFkLaKhzVko8Bq5PNUSRBjQ4aZPuiF1TvWrEKZ76RXjk
8vGQ21Ssrz7SztPjrnMvZ6U7BMx2XBxdoYcfSC40RHWQAlKKSUVvjkqvKbrUizq8EbKk5muw80ic
YPC2PZ0hMFpJCbXwUAvc0HAF4L0mD2Yl+EjQwn8Aa8UTap8C7BZAr0+982I6Id7U3y/9BswWlajG
tuSoMeG4/R2rX3QEz4OJpXgko9nOYXNuhmQJhwN/kGBGhn/zket0/nZH4AaHkfjMgnYL2gXDkOar
Oh9D4ogF7j/TLZonqP6LX3zrHAbN0InAXiR+ojUxI/w1RX+a2ZDF9Qhr4HqT/lb63Vr7LsoExFwK
whnpfdlYtQuATyreF4JKzzMI2+v5FZ47VBZOmJsCLdbz/ro4ku+yg/+3W77aWlPtYqwuZQDxv/Jl
NGTjWAhivXJ61QBdBNlk0dAoh0L9XPX3DRAbz9Cag8Rn1f1I+K/KnzPLZBPT45ZvpsWCsUJ1+4y9
f3axws3hsZ+P+VZeFGephUYvMwL+3POPlavgXfpkewV0crepDDH5xTIgZC3XX4/9daiJi8G+iopX
XvGtI9K8vf7IZa+EzqEMPJpGHwd2gE420HKesO3sWur7NKiVvVErA99SnZZPGbc2xDeQRfJsU5Sd
oYyDR+zJux+YdhrFTo1u+6gdFG5pJ/RYejZdyQbyB/shOYVu8bAAF7vAEOu3AgrWKMArvz6Y+2KW
i1pkoH8SBuS+RgUIvaQxK0NoMfwTjMeiCVnBG+ARiQs0Iptu4BWNwgMsOyzrK9fAsKIi/0hWJsh2
w7NnWF/jeKJVFI5fnbknzDRXu0mwmgbpH2Z8eY45DSmc9FE4coX8NQ3tJwroqREAiUCMTXtHuFWW
Fb7Xlom+KOl8ygmboCp6hqKI62GtLy3BHqa5AIVWl2qL9sQO0LAuqJOWWQ1QzQsIiyAV50ZvdTca
wS2x5MAtm7+zRQQR+I9WAlzKQ94WA8V2ag2+9c2f+fxlims4c/A60A4QRRe3/DUzvYre3ZOCMQWn
STJYZe2CTQZ8LWaSUVlZu++bQ1Pexmkg/kp7L67XWZhT6yEeHc0GVCUHZeOvtQensVaFHf4l+rPr
NsIvq35lxVV1jgPqSjjHVOrA2E4b2/G1fqJ0dxW/qSWitZyFJ5sxgVJUempJOaPzu3mqXgNo7YlX
37eYidpjhcEReemHVR7ctrl/krWmo8oEi8rXxosqXwSCt1LFTW0inB/E0WO4ZctScf/zBXkkA1g5
3PvZQhup752O2ZRD6SEErnNNF1pVGYWR3Ed1CD6I1inPfubLz5SUSIaEg1sd2KtEnol9rQxZ6aM7
j6wwH7V9Gpvj9eoC1IRTGeicwTniJgFWJEJxntU7FiFllxfuoEAPuNP7Oru0iGXphRSj2LhvWf7d
SeNZHq8+Hz6KuqtBQqzR9rAhjuErEE1ORqQuWelbntXDhCaGrXe42tsyr9Wg/rqbYcJ/o2AprO+1
/9HdKt2wHd0I/Pv683HqH2ml7aMPyYBh2gWYbii9PXHsEhaSI+z5+fbc3k6AsFXp5uyc4/YK/zLL
VN9H+W6acdXWo+ybeiRPEpgUDhmhEv6DJS6kZjVgYUJaT5e6d2lbrluQf+ej60e9ZaPgBVMJ9imj
J77hxZyVbA5IGnij4sG0d/ElqoTjhbMUaW+m8GwLL/sf+BR3KE6M7NP20N0zUj76rrN8k8uOAXyq
GH5RkFWjLqne9zEsIu5irACBh4g/4s8Kansii+C95I9HtKeRtuORBI8XJ603v+rm+QdwsjzRRyEz
dmKySmWs6rGsO5vFxEg3euJyIbBR2I3WxddnHjmKNnRi2UG/mHHX0xzwWx8qHW9emxdrj+dCEbRe
LN+wMdPMWSOFgrFHNUhSo51B4m9gscfCq5pXCqR6B9JvDmauI7z4kqGNKZoOC4AfxhlGunt2BwJ9
jjNLHnmqE7+LsZpqSC9hjHkmJGUyLMnkrUVXJzBzc//6zOMiq/1RhNsAE6S2fsQLffdqY/DUok9t
RhwKL7o/aKzt3kRp1uEI5Bi8GtuBZcCAD23c/Gm28UUnoZX6ddq6ZUlWiM1eGB593XvPHrXDDoO5
MquW2Bj61pEtDFmeuhX8o43iYQiEEQN5FbxLQNPH6Z6v+ilrJTvJwfxDGzPSxelHlR2/HWhczYEB
OPEwkU+pmLfuinsh//QfH37WXFnLXuX4VFsu3LtnY2lIc10VqgtQWIZ55BQyqKG+ELg4D1PoYcHV
mDMZg0Hein/YeVbrr8WzfCdGXoYH6E4XLpBllIle2mvcTAOSo418Agbpw12XW4IuAzjGYvpOO8B9
S8HmFWQC84Pa7fCENiPHBonqpY1sYN+FKcECi8k88beJhd+kgZT3UdnoNS80Nax9IU5fC9apOMQP
25IPoCVftZHYJFTzEbqQHrQcqhnKluS+CcwH2PGtZmXyPfonx8cFhrdYJ/PxbCrRTAv03fDoWJO2
/temGpKBbWed+7DPPPordihkVQ0W6cx7m2aWR8rGLYf6iMgIu+C5SwQ6QIM2njumtbUkwjaU5Njf
jjt+IuJWgXwlBS0SwAwJ09OtnKMkMUTlWqk+Jy57LNt88YjpiGb07JjJc+MSmdEBrictWLVciZWf
FSX0kzxEGuzf4HW1CdC9EsVHUQCInEO/QbkUnOAhrE4CTtq6gEX0toO8WzlxN9+9R9TvaaeZNbbn
3SXzstamU5vuKoJiqWfZzW/SdzWoyrKc7t+iYWhw17TJT6mL3g9yvHC08jSkth+7TkwCUWdUpToO
udHrmbk0/Mt+8FDePkVwOH/9F5yIGUbyxOvIPkoqYXn0DgUdAc+i/1/v4v5tIP8Wnnu2KBhYBMfK
QlFunhXlXl2Sww8IOdiJrD7mB4faGMSh49L2wf/Wxk+Us2Z17W7jcE6suAZThwx49gTOXXWiW0Fr
D7LpCP5wCloVAl/734aD+o1euWWSa7/HxjbhISXFVl8FgfkGZUrJc7sEvD9s1gRRdHLh5EQ4gF9H
0zTM2LQhT7AVqgdOrRaEDrbyvrKXymPhPPdbqLZM3oWew0553MPcngQjy9mUhQmNRKpw6uN7P/9g
lg5s398Y785FZKeEZbs8lwi11JpW759Imqb2G19SlgAw8h9mBSRJclUH1olwzch02lw+uM5NPcYW
/clpJzN1IyYa8CmRv3K5UW1NcULwT/+T7lC8mbHlixbSOy9u2HPF2WEtfyVunFuEMH0lF1/8BkkQ
bZSIdVKQbsbDK4tdMO3VE0vN6WulQolIHXNCrH7YgV7YhULcD5XxGFl8ma1MZ4no4GPRArFzLHKD
dWFhQjF8D0GvGKF34LOlvAJslHEJftmTI2kM9/5s8CxS+UQkoFI7gu7BnnyAUjMScv3CbjI+TziN
k7tipXVEuWy+NzGF0R6S0MZuAAcP+eH59whF3bmpK4rqchigPg9DrQC7+osYeixcubBpP91+SkDB
i2kgLg/kD02dYZrcPA5HLLUpDRrHGKH7d5XajmlIDvSR23zziQpKzFIJ/CDd2e49QSDAMLgL2pa4
1V1QRnj7lkZMwCjxOe0oHMrZENM1VMyXLyM/41weqGt9Sjhy63lfY5JiTkJOMRTWZ0pc7aWBG/xl
b23v+prOMl9MFFdqgb9PDkP7s333Up37gqqDAoddWw/RlB+YnD1aPSt+ep7GaNTSWLmoyd89kOf0
CeY/E462zfh7+gPlP1aUWWy3Rj1vhNJXO3xe6rsg7PfFasBWPg2U2EaAAh+e8MZbFl6dKSlcAcK9
K/jeXY6LfbZOZtwgyVgl1BStSF0Gqx5WzIzkUETsi9s6Y8jpFIktdKKhHjibzrin2hKqUuM1w/iv
qHneVyYqKoR6J7XBhEEkb0HjoHsUOP4/fVoFvB4ED4S7MqS6Ff3KbyYJKlYv9Qc4PLVEa2LZsGW7
BI6yE1HERwRLyj9S1w3uQY3/QEhl9bXPcSYukfanaRmZ/HrCBa6SdUxtJ26MIJdhPeUyyEEesg1S
95h+TRovQ/jA8sWtos4repJgEyI0CE4PM2/LIq95VsSnbYXNvihgg3DmMInAZ3KpqnQmQRNCQN7/
wYb7O1iZYOrvFllt6/kJLvk2hr8sczrwbxzK7s3p6f5doy608BhQyssCj5ukBiB4tAekFoKvFlYn
9d+pYX/28+c0jY+uueLz9E9zkUBnYZonhv47+ruOldcvkGrXNlmjeHeBQCnePkaSW2069qDFarlw
I6VBfXMkyO0DcHrEyug8vM67ECe7UoSNPiD1nIbLoXM0MnOSYF+eNAkKK+VfY3E3DuQLnzDV52Ff
6A5nQ6+Xe6eIj9fhiAvxONtwyT1pqq6l/sBW7VquP2sq5jlvHZsJRNmtjk9sZsCPhpYLfaZ3TCCH
u29CSxQ6KX/I0nYWHSyC0Q3jSwbPzIBVRYESL9bT0vDuEEj3I1P0QaVbEn5UrqhH4/VVRmnOlnqg
bBb4uSKIXXlOv8WZd0aMgnThgvrOnYrs5uASUPEvKWF3EXR8MM/h7bHXRaDw8laUkPUhzr6WpjDI
VFIf2BMhhKXQ5efut4WPtAdqIwO4YVW20F5uGyEgIMalv75/jJVDZgVJ1CjkOE22vBkFJhkQKYLI
NgcELbaRu+NqysWNiIV8ATQqJXtDnAzRi4WarOA8rIgmKtRje/x4bmp89A/tmBavbSRav3qlFIWu
cZCdPVkBkkZETdbExUQw43p+32TWLZKpTLwqO5Fu6Muo/iKcbssDsS3dmuGy1tb2lSBByF3+7Fl/
S4eU+FjDxVbZByaUQzbbXw0yxZ6eIED86j++QboA8+dRuCadZFGlMESvlEshbCsRhn0HtOdXYBKV
KkvISSJHUT18kIayrd7EzlHHEZYoLxB31/GCjovcHjffJ0xOHuzU6QW+eorJpuqQ103lj+6JfF7b
zs/bx9R404svQJoEXhU9d4+8RMvdfm7Z06FQT/Xia5XpsfB3O8SI3NjR2GXfGJ7i4YPNzp1Xcp5U
XGS3/itBdDqHdUOcc5cH6cg9h4qhBLlBnDCC4RbAYsGU+SYA44thZONIXZroEDeEDvmtuaj1IK5r
yMNVh1VCv4pTsDzT9B/n1Ynm9Gm9KaA5ABnqMXMRkamDu9/h4LLtOk88BcCrzQQQvBeTbHsciinj
PbqTPuB9hGsjeTxpM/SSLJIZX7cg3N1ueRAvwomWzCX3K+AfN0tEp6pDoVYIgoOIQNSdi3cgbdWk
I8WRdT9fxyPebFYZjdoGuVZevdqfUn21WIISnB7PLvFiZQDxj4HG3KwEYRdVQBapVWz/G3UHGJ6f
H7ReKQPJfnwHmQv/hIh0nzhuSxoIxgFl5xagka4ESuzsbD81eN2VNjeHIIMmdifz38R9STk0FNXO
OPH4aW6T99zKgkE4WeHp94xWsRxI9Fez0UWEAX1E0xUsOfL527VO9hxL9hCupk5y8FEb1Sj+ILLt
wR0AMcY4URM9Aix2tn08nkVSx6wK0ntjP/+6y3xoy4Iw3YZEY9RkNdeMdMA6SSa3kvtGS1sE+giL
WNsbAlBWwufTJt7Zp5Fdi64J3xD4CYoBTgNyk+ckSNRaRRXCdAu9PFgdnnHi9zHu+elnUhiqerwr
1mKsHmr3Gt1WgDs4MOl+IyfscquM3PErklCv5fsCGyLVlixUzqHrbtxbMvDpfgXqF6uhdo+/LhL+
iosV2x2fbImfPQ8WO73trtbWDlW2JAJ9c7TR07DQk5x+DzgxcfaGRKOwm6gebcs13CAFqMvJ1OWW
2e6pzn39TYYfYTXPPJ/2jO2nO6g6EyuG6IqeaGrBWqsd0mB7cfxTF7TQeKL/YrW6lMFrFlEnVAL1
TI68zdsvjJpZTXm0VKsQZrJVwm9Opv1TwWejkvJkUK9u3FPl3p+jdI3ed1SsCkUlAO3II4Xq9xUH
ZOo53/CwEBvZnYJpJkoBSdbnRdFdmnw7v+Ua9TYqEpjXaB30Jl5tur4hVTHr+Bk4tdFUFyuAguhX
dLbuHMyAvyCADGkilpTbRVobl5adcYOJ23NPLvk/cj3JYijE4hhiL59PBYLKQVecCq6ZR9i1l6ZV
lA/US2b3OJQSjblYxUA0iXaqWPfzvJ0xJ6Vn+HR4j8dgv6VWzCl9Z8DQuwd9K6UyOwlwYBkYv2Gq
aE7Ne1iuXoUZXAPvYexB8SpLHcoI4B99pH6TUEgMrYnO7fEG2ZYCvZRKZ9A/o4gY/8S+qacWGPqI
+rQICNT9QL+AJ/R910l3ZgSMyHUw+r3PJ+UldX2bAxGGSYzZjIlqFS44buXbFS6V1F0Jp84SmO7h
4s+c5in0qBjavhJf1+tXjtt/kMguk9+H3xj74H8bLCVKk05au3CIl3lT03fHdCN85Gl3zVVq88o7
K8Nd2VyxZH4tU0ILrCfDayeaxg/J3CbpvtIxmXiSmsKTRkgJwnIwHsZfZybUSxGuAJAzlOadwZvr
mqBUBA4gpvUU1fMFoCwDbeFhU8IIjurdmLcfrEQFpyAXUkVB7QLvW5URlVowm5b4k5zN9J8bmoRM
ubxEnlPohfWWn7IZ0jiF1D3dzMGWyif79sGg8OnCs3cTozKYOTdFMjM2kIAqbqNzMWJLmFwAqwk3
CjjryENmmq+kLFoNfLiK6mL2kKfGu9fNeTJGIld7RRObDKJUnJzWlDz+wNPQJ/Ug/0KS5RCbZ7lU
SIx+HY4VuS+bD48WId44N6olwk1dOkLIFj7MdkvxesqWhD0eJwZNjShtKryBv/3pCTmJqOcZvMF9
q4bqGeT4dR8rjiUT0OrfTcNPhr0ArefnsE7RhFt5uCkc3RgYntz4cMXMY3c08Vp3Px1WaAIp+Lle
vYKvM8tr1xmMOqv/Qv6Ty2PhzoDCvGRq+GEl4F4MChTJNSn5UeYKv7QMsfdkMR+ybIgjGDLhxLpY
JXWLUj+5C2y/HJNhXM/HWpz4ehr1BIZLhGRxIWPfmGJiUVWcr5uU2LtnyrAflXMrgY15jpxb6LHl
S52p02C17Erik6tK1wxPtL5ek+VvH4sKDGEzlUpCRSxuHYx2LxGXAFMrRRcazyrmt9NQ3O9ECw8F
Do9jAuzZDtpMsVKLQqWHYo4nXt5U4ppCTMuxDPcQGBwsnAP5Vq6Oh/AaN31L7PqX+sEgA2zojzRJ
Be6KiZuvAvxTwr4iv2VKjBzoWh9RJgiVZYM6vpRAffpk6Ge821M38EGVpMgDiqEuDkVUlTNSJzVa
EVTck/8CKw2KjFrW0dL7l0PSwmJ350DacrefUxhK6Q67SwQnsJox/yy6jYqN8fjDv5kcGUbgHByp
Ao87w4pGi6330nECYunBeBrT7yF5wymwptsodg1y1UqE9puE6KzWGVs6kvewFlUh1aSecFWP/y9t
xIK0EzqDV3hgRadB/w1QkpFzuMCvGYwFNg+WFDAD62QxfqJfuDy+X+hw1r/NxaMsTAMOMyjAE3h1
eLxPHpwMhHdFhX9uCZiADH3DEcC/IsjXK1Q7yGruNnjpL0WWzhQhn5/ftQGmEpkXYVxyHlIS/VkF
rKOEY4we0g3NO4lwS21m9rnjAajFMQq5Sdc7UkW4+7yHgT1v3RXaC0BgjgnCfcrjqucHUj9vAkw6
TO/QZDefWEjg78b9DVipDfW5qTsQUW1pkQPr5zGJ2vg+P8+KzfFe9ojvpxAMYyuEPMKKr5d8uRWs
qc6VJcFq51pOgUWz+mUceb1U+YVFtborsXXgyjc2mv+XtH/9lWYxBYpY13f8eTtjxn8xwmDc7pTp
qV9/eQkYHyfS1WESV+eMFO8d7vwpFDU82iLg/bKCpcJRzb1bbh5HbFbpfz7MiXs9C1xH/HvyEREy
P9Tw1WWYHpBUEsZyL5cO12U0ALxEm/dD+WugbYVn2V5J7L7uNBbf7+bC/rbAlC4lHUqP/8ybEXTH
IjKMSFeJcnEPyoC2y7ojy5OvdAwByOloYansIJFNIIJdwGOGm3K9THJM4WCCNP4lmnxOjsP4quy8
bo9Sf15u9YAMKX1coOkiJxYIOhEEte1TtMeQ96R7ujeqrU6N/tp8xn2hsJVPpi0YhZcUGnfiwfgT
bFUGdV3m6Lj18tVHbH44AD6zhzzedQqqB2aBKc2U/eQjDzS23KALfkiZHSTbCfMClF1U+fRBteq8
epgggOKVNA6ZyUs8upgZ+ojAnkJ9dtw25xsed+8ORvpXF1DV4F/oI88+HSBcXfghYU9+l5ytHqyR
ZeeKnMKN5Hczm5ame0UXYuRWXdgtmRCdm5AEFFn8FxMIZc1UZPPYM+jenMzuUakXfMyvIgOXSry9
H6zalDTNkBGyTyZY+kwRaIKhNITQi+t7VQD+sAROYP6nF+IGZFQPgHgAXBVSJt/RYfW0/igZCLLJ
jrH6pH9Yw7I5e7EtTfra6SyNbR+t5XGehqQy9C6ZjCh8+hmH4GQcdoURcJHXOurllcM6+JY7tGMw
YeI/dc93iNIfXNhzCjexoRAMPmhqiku6nmiN3HjSEJM1XRQTuegeyS1l6Nu3UJE1tCq46jALS8t4
jnw41Vl9Ka17r+Yv5uUPat3OJWlvOUmrMXDWUZ9zbGulA7003FL8Hm5fRinyCqRuUYlHQWpB7y51
t1hABEtrB2Zp28T/plMKdxwBetuItRcKHi4YkGwXw7+Qn2SzeQEOX7ANKeGNGh0lhea6p6gAhd+r
kkIa3v9DIypsY9BmIehsWOagl8wYJnoCp/nhjg3C327L8QoC7WqESM5oDHIQI53PqwCXP2C72ano
x2KFQRj5RU3SU+SmfhSiUxBL23IKg+2w5ndoHwnQM/L32ZixaBY1vFmp8weAoF4DtCbBU5L42tGu
K079vSZ6y9kZDAV8yHWC8FlLMS0X4ngDWvubJo8Ys9WHjDuttPfoZd4lzjIy6xShDTlwL51IwfBi
YXx+tnIJubBVj63XBAaKCC7hZVINSWcp1EXjwx805SonVpU0K/MTBXth18yvArCFVWr+srupJVjB
srqif7k9p7TUHD410XaP5aoCJlvWxWqKdFuvt0rwGHT4aui8g1rc+/7BS390Q3jPeHpI8Zea/y2n
B/jbFgAHje4SHPQXI1UIfmMo+dokSCGOVJ4ihRjyiQhS+k2+ZrZFxV4Z3d8elJjJuCMQqysMyqb8
1svhbhC/ha4r7OhVYLBzKTqhGLUAcwgpZXfZM3Mrf+mPu2kAZXh88BhRX6H8SPcZnLk1nnPhk9Yi
jqe+pBSaXuHQwQVvBjp1WiH0v8qa1wXWFWilPwR8f9CCqzKFuj/uNFpsH5BvnlpYMFefbK3m+/64
aI5G0+7lhgBD2DZrLAblO0GvUGK80H/9pSEd+ny83umOhQNz4cGnN/uZ6GH4963E+vzVOw+5MTCg
rH0qSqSllwAeRWU5FVQ41tUUkP3L+PL+2S0X6a6rBSoKJLXveodWd2wlXFmmPfhi97bCQ5xrVvhU
kHC+F+fVzYrq8TCMUshAjmTO0aU5uYSy/imJlmlCiO37Vb23cSv7hTVTGcwoysnP+M9M8+d+nsHS
7IICg+fhEt78t9PrFHEmePcp7LFU3XWLGfpMoufPI3gb+ytmob+acWqbx4kJdweoEgNAg8rA5G7K
rDdd4MtcD/rKibmOik7Hm+qNk67Qj52ZN8OzWZ3WZLRuzGBTDs3eDs33TZ2mooon+0E6/IjYMpVW
ZNA4TrH+GnRwVBD8HY2UiIGUxKzN3PCCGl5Kv7XxWWCB/IJDmvgHTcJexibNjZlrOLZ7TdTxCpq9
HxfUnCXUrF9MseG7gIpMQNjWpKxz+gtcK4x1eQnJtVAqquBmr8dICrqv+rPJJaGcqQqzYX2L8vjS
MBNaghgNRXL/QFHrano9EmDBiZmUZGGLUqsrnzEckipyeQD9h3Xm4sN8nlgVGEsG/5XMeJY3mZgi
Un6DTSWfnsGeLHxtzi5xlxKnGTkhNgf4nmnEYwVOHhG6vAmRNqL3modsIKuecW+0efMS+roZNNTn
/K9/tMmPZfMvb+bSYjKXVY14BHdTC4rf8Eo+TGzAhRxK9TkiK2yWvFuYwa5BLIJAp0V4/Wd58PLl
bZX8RzDkTkStlwvO9Ptb0MJwH4aZotet+EcYlzkJBaRS+eRbhqCOoaWiW0ODztsLGGj+NodjmSF9
7+xdv1WKxx6KX4yDNsdNdWu6pfUklNhekLaNz5Qf+x2Omvym3OB239WMQIb6Vz58Xft3IWuDBXW+
MC544fiXgwhdyXaGxs8D++lfnJ+4bXsukazNgsouXGe8XecVOHW/UCDiUMjTcml7B5jqCiDqnalX
+ibTsadZ5O535yDvokzJLd3yYpBH+ws68KRS0PVemo7MYe0q4V/nQH/ZaHrYzsf5aa1W5/P1oCUY
4o21k1pSYwNiHW8vfl3J+V+4fmifxATuzvt6bZet4Mw72Y07iTO5JL+xsZ+EVR9+PIMA48yxZ4+v
+SQC6wRD/PdoHqZXMOxphjzl+IxW6fQD0D1uiax1iXEWA/++x10e7jpzH7MYv+8kuhh3XGo5KTPv
zreyqNq08RMnqgsNCWX7bRrVVOpZjIbhqPIIApR5UPNHBc6yFhJUDCyf+VRAeysbygpH1mgkTRCl
17JZmSupxFRZS33J1m/hfnTfqUXAexPc/YhlSYWbnONNfedPJ3JmQSTalZym2wBR+zCNCAoCH2bj
KjfY6gSXs9qPwzJKfoQXvO7oBYk83K/n/hq5r+li2s3UOEbKwUJImrz27saetSBqSwYWJOJLcCxE
8WNtIRVvoJ7+eZe3mmIoymE3RFDo4XIdmK1HlkuxvGzIHATQYzNpTE0MCRtoGV/ypTufIEWOqesB
cdhm4KsFelBO1JWvmx41hHVZCVXypz+1QQiTqCrFbkzIkVvmTj6h80uKfI6RhlVH382cP7iiDbXu
9c+z0md+AVMhFndYUpD2q89j3HJ2ga9QXXd7EpiRVCkrX3bGqW/p+67hrYhIQjaRb7ACzAGJEJsM
ejfwHLXqwsdzU3RHbjOnQ7ZGE+UVncGuH3Aix3GAW/GGYqazk5ASSh6aHvPbc932xu9lmwyjdu2U
+y9NDdhIw/noki+GGYflhqUtNfrhSSvfssIfuuHiuEFRCcOTAWVlIPFNO90mBu/AP/1O8Sql8q0F
Pl7dUzxid1yQ+mN2GobadhsOmwy6FKbgbX5FBDNHWUn09uNJ4kMargTlswZ0bdWbsrPiEjXxV7A8
GDSFGcRmUGyUhMW2exQ6PxvgNSQ3k7vkFJgL5NsaYiqD3G4hmMTIi7ZuskMgiW5CHc4lxrFcp8mR
WNFQelwxbqmjhSOCf5GwDI/n1GLxyW7pEWxPmgIOrONKOzrZhmTMleewHTuig7BEynMQf8/F5WPA
CSZHoekR6XA9ds4yovcaU0EgC2IE1g/ZhGYBPPi3pRomNGK8h1nr6BufUMI7XIvCJoisd5xtZd7/
gdXr69EzgFc6G4HBb+b0X3MmhYRR4rqrKoCrmJ0uMZZJ4xIg1DC4477Jf0/fazNoN6qfs0lhdDkL
b4YJ/4sq+4qQ0e1TIZvZUqUUmKqduIGV97La1BOnTPZwwtxwhqesAhq4NZmkIsOMUhZnQW8uU6fK
FggU41LJRaQ9+n2JC1iYO+kAf8jwyA5BKtH7SHvI85a6rt+9W1TU5EObdil4/fFgY29iRCK2B/TF
rz8NUmxH6gjNcqY+FvQy4XQeqdHAnvBYeKinYgahGzPf7y7acb25P0waaHnwvwKaKNdFjjxAP1fz
R8choOSV/YeSRQEZ6xQvhpc96r+ETc+z0o6lTbJ9yBtDUPh1saQIU8MJDkpLG5N7306N6DdeRIj/
x8nq/Y6xMcUQj4stcY3PsPtiyeiVmkXJJFUCKSJ1YqK+cqZrEbNU2+Rw16p3JF35rac3cxnUp6kV
0Id+Rb/E9iuNAuYm5o1umeC21EKnp1KQIgvGAfjM+8yNqEDcGDxkyvj8z+obS+y4e9e8wjfYkQq8
Pev/LOYBzFsSYssBdcvNZmKF7bvYR0VYkWFFk1am9iZ5R5fFBMqbWTRCfS7QrWqUhP7Oi1XzSKai
HKouOM9raxNHkSy0ran+NP1HjP8tRH2sEd5tvfvaxqOWexLThEGH74LjdprNx+vaA0Px9dTR1oBC
1kwwa50Zw0OrXkqlBctf5MTYBL74vIVfNfS2UiABrLPVRxcUYehRyYGm+tZ1oIFqxXgup95srgwF
emJkE96O2uJpDJouovOb+7CNfHyShpBj4voSr19cNC5mwg1gkwoR+AZfAD2UZLpyoKdJ9Jur9I7d
0FrZC4oZmSZMRU7kmknms1UGgdzPh7JGzQbLxPXiPoZ20SdsDqW7HMv9l6SYNV/zEUfI3Pt9EyP/
UoDSk5eaVW99Bblmxqd5BeP8Uta27/r8s/49Xid/XiT1o/tzCutbLRhB8fPfyoURdtdvuJp6fG4Y
yzXiW3kFvUqYzki9vmFC/0XckooSD0dB2ckboDbGxIYQrribC1aKqAq3lMjxfmR59CzcsBq9f5ad
vswpQwPnZZaOD3YOsu+53iXp+nqaWmcR88DSrJuk8ZAZpUDHco0wNjcqJ1Q1O9rraRO2faQBu7Dh
7+atVDr+TDZaskXR73twvxqmlPUf2iyL5Koo/Sw7HWC2Bp0x1K1HOAgPtSyGtYcBc4HSLQRL7J5S
EgL+AO1QeIpLf9w+Qz43jQfDi5VyQdaG2v/VjcIN+105rxt4sp54bJvu31DsPXQWiKm+72HnuuD8
Srf3GdLeAkAI0770yPm6t9XBd2NTMmktHUJlfDTbuTDwYeJN5XVrRt+Wb0yEzE/lhioc25c1sZFG
CBfuHtsBcWSIVEmy4ORXShMqC4EcMz7Nv6NEMq/MSvkoAIjej0Yo62gwVcOoYbtf2isRfRejEO8d
JyqlWl73QKUmvhNlIF4hFJAmB/xQa5GjvHIv6tqshLlA/PfDuvxpg/rrQ0IrRPyzuCZTL3QT8Lo6
9pQCMfml3LjN1KbZ2mg1+IFExX+6pZhrswCX3qV3F7Pel6+IKlEwdkUrUNeyeJzTEF6pnfVHogOn
qlQOE54orzWBy9hQf/aSfTKHRUUNxzHT5CSaWI4AW3S+wij4qdxeWL4izRsRCcXQ+IE6BKLDF3yV
aJlN/hDyAkdrzijfWBQBXov1qK9CUWeKsuSfIHzHcQOvIBrDc7X11tPQsnn0Bj0HvALoGlfI4ZjW
LgS53ANqwXIol/BroFmIgXOyAYEYgqEemEz0uQWXMhJ+md9RnYnoGVVz3+z4jtUATJMk8wtwGluY
85aDpLiIJLXhPMBVEVuQtXXtVgV/wC20F1Vyz0+xpcOkqgzUQtCIefMq2XySxq4OBTzuG2+Vvimq
eR6wnQh7z3v62ZT0SsazFxdJfzRofuzihlUokm6AvI6OTlMwl/P2XzM1J76jlaFw/I6pmHG3cnBy
FMdxZ8QFU/7omuRILAqM/TdjCaUGtoh/Y2FJDSoK/+tPtd/W5T/Fhf9DA1g1v/WYjs7+DUHI//ZE
yH+2J7g3tAx31faiMAptNPLDD/uHNUJMoB8Q3NKXKEj5lTBVSQkNppAMqAWV99Muu81xve31d011
yVI5cS15Xaglz1p8r/+UqgR0+bHMAtaVlYwEKp/lc+T8p6zTQiM43fba6TYtdobORF2mjmbj2u3Y
zXJ3vX4EYh335Gf9yJf15JR4Oczbz/UlF8Cyd/0D69N1sHzex4iU1o+KJzqBjPVYRcrgcRWa0RFX
ZLkBkZpU/AGGj0pG33SfV4079IjGOxOsNjBLmFqStzpnljpb86TG3ynrnHWOQbhSHj+Gtt7s+ZIz
roMWFMpwhy+jpbuH7/uulYK6aZWy/mc8tWk2UOIzGpBBTW+e++sujE6Lz8lotqzc/HKthMdtsgGV
14wFcMhKKP7qyWflNeqrlOIBMKRDSgACzb1y+yoOG6DbOjR0Wm+qZN3/uG0FfiUk/4K81RLO+Z7H
9pcwCMQmo8RiC+Vr4MqEyf1zfsj4AFPz5s3dMN7xeOcWNYlEvjcbfq7sUqGJhIjvDeRLCWkKaYmj
rQjR/qN9L9fwPj60S6Jt/NQuzb9SPUrzgyxuzo8ZNorxoDLZFLg5HcLMbJdcA0o6RZw+iHYtoT+Y
425qE4+ouOFIM1t2FTciQ90KWuIwO7RuZLEyJapXxw2T5OOvQnAnS8ziGm5K3eoqBkzBSNzvIw7c
+I5hrC3RvQPkebrzKFyN99Q+XkNNLJmLf4g/IzpivrpPd2IGZZ5fpeX1WGey9Bq4+z+Rtj43Bevg
RSjhQYutF611gWzfcXQm4VAGHyfo25YjBbKP9fFCZ8gZqpqD9VSQoVZJTuo2nNOnoHoaHNOan1zF
TXzMbnnPaydT0qWhoQczQIRabFNC6J7+N+RWoNO8ONhHPvejMiGRN7lNZo5H0zj8X+bGOC/IsPqu
Wb3aqzL6I1bKlruVC7TEBbm8ZpclZhrDDnmoublOfwMIM6ywFO+V4um0AaojvBKbjwjMF3h6LymP
1dnlJaNWS9A+BdtveZnRhWTTizeGjh/s51W9iokiCiE74wnUDvuoWrj81RUppF9w2AU7p0i/pTTa
dkvUn5X0i7OvcgOnPuEG7sdhEwRm0z62O3v+HEwgiEjMHoy0m9OilcqwxImSBFddBRxHPw6BwzaI
cuOZe/ScD5DSeoubdtch/rnt9jqWDfk89KZrCW6roZuq37PbvUvGYcrvX+PFEchohAkt7n0H3yI2
24+ZlGR70X0AXLVUcvhfjYb2RqL6ZCCtYFBWCpqj6YsEpAhSxQnxVzsEW2rIkv9aYXrSA31VXWNE
QPlTH8svDOwq5K2Pnx4nQlxioL1ElNcXILBkPD+J/p6kHGjNDk5uKOfE/5jf83WT21NANiPTJ9NW
U5Jp4uc7pIgkVXAD9QHPpx5BqZB7umKZF9rB6B4CfVSs0gKJ7cWrGFX32zGhagz4jm83dgyowLXF
ZbAXQfm5aUSTjokbIvan9uEuvuvw+Q/cqVWwT+ayLPZB4yLmQU4hTSuHSTMCSdWX2kDmUKqjF679
7uNp7AfiSABbyExMXXVrtFFPAZHRHWazBUNc2dHSYtndOf5R/FZd+8dDgrmlJJnlbVSUYxgbSm0I
fgLBNFAaFLPivOvwzTiK25laQ3sGlf4oFFQWOtiU8KOOYcMtpMYrtgFImsKQIUwX6AYGGy2wuLbJ
xdu1hc2o9Q/ZH7kvQTUHKBPwa4z6IGKk5etX6jE0lTOXfRPazWp7KVjs+oFIRvD/o3RFkbQKRz0f
a4pUwqUURbyGaFF4TMA7C9WWbJ/0viUonYxjFP8nDFglXnot9s6759tHrMBzAWzYgVg47YzcI6PA
e0vHoY6u3jD4JH5GxZY2T+cgn2a4hC1FCZ4ApkvilSCGYoQhhE+shzZoBqPZXFmrgBWhl0qhlJnr
LbvbdwVGmfM2niinDUJFBrNAKh0pyUUuhRpOkqnyYYXpk/zQe9tC1Jvxvx1lYJQ3uwPJlbcu5QKG
lOTnvRNGjPTokm5b5qKMrGS6u9Y+MgUthgVvTqrADTQ1XhApFrD0F2QW+I1qULHcRzh1kvuLcKop
kW1lH+GuH2YEjfP5PkXOlibvpb2okWrZpb4i1+CP6xJqCtNEEknh1/oFXA15bOZM8RUayKhPXb0q
oY5ZKDvVyqoBRoN0iRoyZAC96IfYrbMF6Ru97A0X4HBygDCmqXKWopCaBMWmBGS0+hRxxY+1b028
nEzkDauv+kqN9dOwLZiOor+THM9CqL8bBK/7HJoqqPg4LIW4f/K+rLIXl65T+l8/mqexorlnEh5+
nIKUtFire4Hd/gdFuWo8JrLzkQoarAqt9O4fRRVgwQFQZygTYFXEnKXLBiKOqNy3qRdIS7HNSvHi
iajzk7BsPSK2QPyAShLdLqEq3n/2gTZztB+2QN+33yo07zjgkBa9UIzn6WllK2qpIPHx/VVdHMAG
iHA8+KbFPzI4E/3+MP1Gk/2jFqAyXukL4VR88zac43Cd78w7pxFc6yr6Ke+fwvM08hj2pJsXQtwE
ruqxiyxDeAs4Lc7RxyVOcIpfqCbP+cabB64MF2yYUCwxarR8FEviWhkxfS/HP7AZOB/eARdHaZ+p
1rCIL/oe15o+xM/xKQPgwVK/N6FgEoZQJTVROTgP2nWarpLH/U+oKPVkF5cUivsrdu79DAarGTWt
/V4QRtEObediilcLlwD5G+upzmdzZ/b597CfUpoCNZW5jbjJdmPDCmE5CN0YyyI8wJZFvUUM/q2k
jHvf+Q9GSAXVWmWxMmY8B3eVDvaNvpLTakGP7Lctnv6ymAmmTiPQ6jYnLLIkCTtVvqZKGFLoQ9tn
GbEdPZqdpqib+Feuzi02esATGCf0faQEtP57ZqFQH+1gohIylI/n+grAWMwXUZVf0ddgmMt9Pjf4
9gL2c1923/3ofnPxZPk3a1BkjGjLyc/JcYKtXPOlS+coPOSh51YpS8olWfTrjE/XrQ2LcsdUcGJB
L5MAA/HcJg3jVDLP4kz7v7ao7DuX8wQfTHRuHII1xV1yQmZuck7AM6KX6DIQGz0/EKhCcv4xkuQ+
ft1VvWmCPmnj1wV+l5hfjiBueAPS0zImmMXqqJ2qAeUiP1NJF0T48p9kEsI+RZI/kvD+lCSuhoxv
vU3UCaXme4d13AjQPDLIYCLCz2g/u9g5Fdl5W0D/JG8RET4gvRCh0njTDiZ+N9fxlpZR3om1NBSw
7Uhi1aBxDhI7c5zqzCmFE1xZvdXs3ssKR4nqEjbbRusu9Zq8J/hY7+uWV09bJBiTcGUUKqut7/C+
fHApUTwrfdLS12aw5/1Hgj5i1MNNJ1R4l0aJ4MHw5/6oxuw3oONKrYOi0p91qd8lizT0ORdBNiXb
wU+MhsebrFUAMeGQsJWnIKKmZD/CPc/eNo49WHVxWf4Cg8oh5VBhVt0JhiqePE1cYmAfDrZSrvMm
54xupBFCidXW7iMN+e65yNnYy0zrDLEOk2rVQ0/Ag5OxnjexjrwlTqLLZfmoptpIPQNR9MibRWX+
1UfLqpimloBBvNfSGvwOiX9U/y5ZZf4jSR4birorKtJiV1IWXgf6DxthlGYQeoGr7kYeWYkA2HqB
sgbXPkseKVAu9jmkyF/G9ycMN1iBVLCPxvKb6Uhw3pgMXz6UW+AZ1VtVSlGgWJvmsKNcuUeAWRYz
rghj/jWjfp5KBnWCN2SUl/6mL6fNhAm2L6zjshgGu/sxK+s6MIZdTrEL+/V4y95CtCTkpLiRLXg8
/gHChmuRanNQS0QHTxva/N6bqMteWj7L1FiMqknrDdIQQTIm/wGqRjAaqGXYqe8ucL27plx+kTXW
zIEfg1B8bxtRCQjFgX2WWUzmU9kG1zzQmejjGYuDxrurrQFdD+WtABnBy7HLW6pce+XwZaEt0Jl1
eIFw8/IDaWRRuSOgoz9Gcugmz737hBAJf/lUaZnI4VMjT/yVW4j5jlsM9nutWMdqcn+YYVki2s2N
dfz+CSLYZ9Dh7tIwHAjYS6TPauZfZL78+YpncymHbq9UBQodzxy5KEvnKGVkWc9xH6d9SOyPlDRT
3q7SzJX3wNCzbegc3DZUfk/AXcSjn6xWEvxSItMOnFM+yDZV7zx8qzo6PwjmxYusAVNHao13g/PW
QiFwDjA2rsBYTJgEJ/UI2wITzyGcpEfOfRAB9wzfoNPdzmdpmVPsOvcjeyI0lXhFFE6tv2At2MhJ
VinKelqhUneGKVrxM2bbwz+uZgZFD+Hh/5W14ERdSaZ4HSJLMbvuyoD7oTBr7/l/wB5a+zSNWBHY
PmfgXsNcsdzP0uo8Sg2tJAMo4uWLLrdTmNAEzOH7N5PKNTMCPvU9VbT4Q0sZZwfPbuYBLvSn5t1c
50tR5VywwMn35sZQvtguuLINUY8h2wRNrI3TaPgZ4zwQ4h9H11qf2NBCjQGoSpHN48Ul6U1ZrXMs
hRmVD8/g7wN8AVqkly40UfW4a/m2gLYmwZK/pDAcRMBvWcEjZOSWLamDOakZFvW39c7QAibF+Am3
P44kzUi+8IOkCrm2nTvOIa5Y56X+5+F4xFBzz5GFiAwOM/mFmyqq/+GehXo/rlLuHJbyG6oRIcOs
Fmw7rC7FyOd5EqvHiMKXhibEpKH1unhKP/EeLilesU3qRHx6OcbwATkU1BewMv1URPv4EB4K4OZu
fZlrOfeXJj8x1AWhiWDTaVhMvzUKSXaDR8aVEFu89sywXUwUP8kUg3l2nNiughqGBnAquVGWyZb5
+IKnPBN4iYkuBMUlZy1oymtSvwUevpueYeB36Oq3/KEtDIILieH8Conu2rsA3z99+USav8093Kqe
fDWxAO0c0cd4g7PgsimTFCxR88pcV1qzveka+jW7UoAM75+sfICs5AQKzIzY2SR8Yv89vJ3Q4vXF
lV8brw8l79Q7LC0H9SlWeT2aRgRVyk8GC5OnAU88ZxvLqnPa/krutcY3wpNg7y9fhSD2Gp0gtESv
SJlIuYae0QAUCuT4NXxwm2////wL2ZOoP/ccJ5JqjMzSG/IPTWmk2ui28PozvYDXTDVUv/uoLWZy
Mnpwg3qdOOsEOSMElmtqKJi9/7bAmYkg/Rj1Q4APMxtEJ+0Q/Xod9BSnVZTfsbVCPiBDrvKoyJRh
s3X03ps2+Y0Elc0wCbz0NeOpDLHW61T3EUnWZ1dxjKJp5A/rL10bmt0sTxbKvAhGvkTTEM1v/yRO
b7RaghSO/2VxyHo1oUBfv2zrzHIV2DyUTK07For0NYjiSXQcLt1pTNjIzNpkJ+mW8zmryypxHARw
RPqjhgA6i5r4DLvbESH29Jc+Uz9fScMAAAxQaHplYrY3ptPS4XPFNvT8A/DjxRM1ZLRX88IhUkQ0
E/nECQ9hHnuplkMepmESLZjOtR0Sw0sstS/vvfen1/kEcMfCJqYoowEA2g4O9BXmcbS4JF5598uF
O4KMh1HCStoxkKaBC0A9IFTovoO/o3t9cn3PR3ZY0v1GGxHhogjqItfDOhXZdAm7BZDozZuIS5WF
MES5QiGEsHnofIscgbKXQx8YBYGA6JrmIFrD+DbAEfrOnzoRMNxS+L8/FrFh5AIJFvyMZrlysmcb
WSbgZFzrNL8h+v4Nb3XgflqILOnEGPusfXnzEgpduu2NtLLwTERNlJ3reVfHGM/9jfH9SHzU7dbl
r3x69nkfAOuBfMPjQqPV7lF7uE5ctTINl5Xbs28mVCikC/HdfuaG9vjScC3CqI/U/4ogJOsSHgg+
TDHjRB/4jz7KQ5uDKCUwe8RWTpQMe3kOpMNbVLulsZ+faK5EMPSdKEycU/Lmytjg7rSivALyPqWQ
JiYKbdQWqOPAiHgV0TR+/kMDRWW4+RNZwO7O1CKxTqwWDawlagB91f0z94xd8zETecgSXLS/o/LR
UG0DRQeupXZ/nYma8Dk5HQk9d4YbobMb7zo3ce09ne+Ey/NE9uUCTCPWmv20EqVqz8fXq8tntKpv
lloue6Ev9eKdOVWmaT2oJfMlm9AvQhVX+ud2QzWKv9DUaT80ok2/5dHnXEI6Ski6iLZZ1SHnl5ro
RDKeO0R/JnLTg1KZce8H3K17xnb/s1as72ECPMICSUmGfSfXCcuuJ687QQfnpa9PMys1LJhOz8FJ
4abqS3s1drNcdUd9IUcCPMTFqN6aNKA2DUZfTU+snwtaGf+JCZN26ZCa8haIU5Pw6Kt8Dl+a0NRf
SSUqZOrLWQ7A7eH7FqNg3A7NFDoK+PP/Hxsc0n/cDTH/zlvqxuvvdBjo56c9Pnob6goHpAWq4PGv
sVVhUG7HtnhPl+2omJz0pywqm4JTxZvsQzoS3Vg0JPOS7Rh3lIQxxKvXraLCV+eTuY8zI4HbrW2t
42eVT07MTLLl5f8EvOrx3EBFYvDyyqaIdmVj+cvmQX7Yxe94/3JAeoGUEqpL5KZIDzoKEAiqjsAG
vCTc2grkhpUcstusg3aF0rBMXvHxjlc+XwZfI1714eSXIIuuwuGo8rdXo3ozpR9Hk09Z2VJ7cdXb
0MN/nqWIWzD8m9uupuBbbCqrD8of8YdmZjVLA3GlQEh1vv3jAC+kVj0sEDEQ8vKv2/A70YGco3Nv
o/v5/tSO2kKL8fg6wv6JLziJ71PYFev6bHC/1jNYZbXJ8CzH3wX3RFGsixsXo8Xz+lSZLuRASNus
2sDGV7N6oHbRKbZcaGuR6cGswNbaX++gzl6qD3qhpX8nRcHyBsJ7VFURQIsAVzd+8d0fO/oiHkh0
VFYZK0LXgYRMdJcYOAa/zKbkXa0CK1cZgozYZxu2lvWlPXw5IB0zbD8a+hml51y2qQ42lRnAVmoD
P5jd+IiP0d9oqReJ4u+f/3vsNiLmsvgJktgaqyEwx3SOUBirfRWzIlJ+NC8/Es1o2SoCsp8vccER
MHj+y8gkDTanAyKdiiK46EtDptgQg+gdmXPPZZcyK8lnSPwIZtpoWk5bafD0og1sVxp2oQVA2sUz
Ti0JSTtMK5gjjTnLzdNCEcwphCxRwHold2hG7JPbfk1u4A2gYhewp1hbrPxO8ea2++Aw1OGvuppW
GjwSvljIiHooR8fP0hJWx7UF7fSSIuH1ltmUxplsXHVeH0ZeIa+ScLBWALhIrbJNZQasgrBRaKtF
/48gEYmCzbtsH+KpBT0RolQUxTYA5Au4z1jqEcGk3SH0El95Nd6v5QAOesj8Hr+AxXG00aqUYGvG
fxYwmX5DBk3XS4COmiiizF0P++YC0QT/AmxMMh2PPqymJqsrhJ/HzyCSLrQyHhMJdPhE9g8DrEm3
BdixMR3HiAu9flCFGb/0hidpqbl+4a+CcPvDg1HwAEUzXE1gFZOac/ci3QDvQv57An5j08kpO+4b
OlYvmcOfGN3nvK3/192P36Lea2tiFMrAB2u7LiWi1xlI/4GtuNXMcL3iWwIZx27Fl5HVndVgufkI
MqVkJ1hVkhjB7dZwsuIe4FPIa5nvVssAZVB4byMnkFDepixYUqbH5a9gmkNxFIANJ2QhyAdwGBJg
6AcBwpoH0A5HUgGxnRNl5bfZs3YMxklC5BY2cc+eYGw0LCNVAXWzi+Di2B0Rx4zFqejNbuwQECa6
YfLYUKC5PPRl6MZWd/irPnejTyS681HsBPoUAjdyMwn3JMFPWMUIDXVXTDq1wi8fuylAplLHUEc4
WuKWOOAQjol0/bawMIzHSA/7nf/MGDKC9Iy2ujZ2/0oPfGA5xYAYE2ZqSKlsFSZbtQjdkxAzMaKR
YGcm19/+iH1ubv+vvfVrNhjNf67ZFK8hJXEe+LxwFGUN+pXYBWrwcfGDke1tzfjq4U6MqsPcAbvT
wKljw9UdF/Hf9dLvCZ+4xdmeiCFlSY6MnX5O6mKCcwjqngb3iUKDQtOL7NXzt7278DjW2W6cNFAn
k//aWedp7dyMDNW5Tkav4cSYgNsJTj7HCggxE6uD7YR/sfv+zP94EIBFdY064jSdoR+KM/xpMoRQ
jTvBjUisoApqEJkiF0K1juUy3TJlUdj466JIZOlSqUm8LRhnb7JWyVSbOS/tkydd7TYbY5+aAehO
xYQu7vq0mx9tjYzd5jvHED/ql3tC/xGa6JeZk5D9wIooKYkTVDzCu+MxTxkAFtj+j9vN0S/1PQIW
CKB99m+SJMQupDxvd8IOTQ3FnKQ/STRDOtDnb2HwFZkl5UiQv53yz/H0UV/6/TuAImKp5vW04Nyz
xOA5FTLIkYJcKDOo9nyB1zbH74aFjX5qvSGOTk1iHJorZjb5r5H5R5rda3PwLxWKIzXxjxxy7wLl
WOL9D4OBXK8GW//FkeYwkR8v5lqOnRfJqYvvX0En5GgQb64LS3m7VVUxtxqBgPFPTDcSfx2czqN9
i+zbYMTN9JqutC7kEjPvfrERLlBkHxubMLlJMNhvDom1kvneluv/u9IFQuKORpet4c1zj/cYI54w
oAIzIxWyvjYE6yVS/+NwTvH9k/ZyddgK7S+z0SobDILpvPwBmR3tZGh9pq2/fS3HJsnwrVuJUlQ7
HGictqItodxDgND4yO+h3giUbti1phnzPC0b9g1KqUeg6OyBeSBCouVxz13fjMiHcuokpvE9qSfB
ATgQbmQpoHirqZmGY1l+MJzEEhZr0MAqRAXdXhYx8EEfOK/ai+RcQswWLOOE6MNO09/28OeTsO31
Bvhm9bEMMnxQh7PDahXTx6bBgJ0v+VEJFSukToF1fQdplvddgORQUtwW96IPYHxPHNeAu6Y2hcXc
IIePjrLnVWh7R+Odq909khYQTuIBxMSGo9BGJnVI/v73sjVkBuXoGKpXHxLt7HLUCZSfJwCZBHKz
4x6IdRWFD78MCpcYmHxArZkTuG0M8QsdnYiwum1oBMeOy2ehJbn0PJGX3Rq0w3E/Wo5tWiKxbrWQ
TVl8pNwI3OXOTTtYFdHwVE8eBVZikbXfI9BuakXRoSsrwLtlqKnubMisiXtbmcPXoRg7YI0qpSVq
vfDcEJGzLl2Xk8Dk02EVIUKTj4RiA2Le9GSJfmTIHzWGHkODa2w/v2jAy3vvuBtBrXAm4hPq09PA
Y34zpxL7ZnSD8/4pxP3uhsOwuctlpP4+AQvBCl8G4FpQHWtonIC3wdu6YmNOidN965nbqUsxqSPf
bKNN2Rta1/jTtD+zwgaaIgyInfKHvUGVEMuEQxyzhv5zSOdlh33lG2DIWflXIuQhV+1rKmbIaVnt
FCEdDhhMTU/XUrbFqtOtp9mCZWYeQJSWC5qXlj5agwLcDVvPbuv7ZI5OUgrw38fRfnOR3FtlITd6
WMjSh6yk3a75bg+Qd5UPHxFyhhPGCup3fl6VcZTxNDY53JlPxR5mDKKkrx8gaZVFev1OBP//ZPLS
cgVZwUCpMA6Wfsgn05NVqJgZBy/V6GDB2pQSrTXeyGWryrlAL2eFXbF08kZvzzsyyNQ53nd4VoEc
bXwN++rto00Zd+36wtIugC7e4FI9EQBQIhvwx+uS7JVkOu4YG2/T28B+atf0U7y0kxiVyXupYput
201l4PeG1aBtZymYv5M7TjS0LJtI1koaVJuOSLkef5ytWK4frAoYyLylpFBOoZv7W/V4ZbUUS8dh
fhNeHRjmRNMV2h0BsffkMNVv2VOCBMTQpHbfmbzynumsKJ3uGBxbLuJc82M31KCRwgwhBKvzMxbx
HVpEAcgZAoqhvmFG+JPv1HbK2ZjxbD3aO8tvz3gXpbIHBOl1XfM0qWszzrN3mvcSOAYwo3VxwJbg
HvYBecS5m6ESvNaxkXi/OsAyF2SvpqTi69BNYeZn+Bqi2DMVE7XSGwSAK0+1gcsiUHwiWYsp9bzs
TdlbXK2DPnRutXh+2kQsV33tfpzLTAC296tbsOITwzi3EMfqe7/dkNYWYKq7wW7Q3SCV8+hk9x6M
iFexbY9ThyTAav/bMY8IFgeuub5UfQoEz2QycCpIBm0e57p+Bjs41lV7IIvYOcQ3YP81hZ5ljhSl
TpgdACZRJlf0NBjNE9I9YQZjEbJldummXLBC84lvqXVfCqGeB7FBIvph+hlZH+r46ec0GW86LlmF
2CIG12/js358qkxoqLuz9gQnpQD28SLasWc83BnJiNYMidTux5HX7y5noghzZyQunI8OR+AgN4LY
P2n1NsvMmFiCG2wDeWaGt6ejJERM8ik0cC/L4ad1WbdrS3Fl5xjAxTb8a9tECXWDOtlcsm5hubfh
0syU3xMi2wiuOceP80m6v3+YPed9QJ/nkKrejBegtNkV52vZTSHJrCLHbVEixTXsXS8DK1iXSIbI
PdTFeqZhP2QKXFni5LylBvo/n2jeoqlJPBH5tHNYM2ccEk09mb3CVmVeCbB1ROQc9Jek6ky9kT3V
Lv0UJRuaorlFHTdHxoB0qT1kKi2hZ5L1PHPArcWYB1jCLz3Tynngj6ZQmTtCuASRvNnnyrFxjY+F
zVF2JoY36fw5P7RsKxwnU5zYmZPL4De4+OL17VJNdxISj3WjS6ifEG7nBWXA3JS7Eb2RNEVTks6w
LayvKcUqGH0tY3gSHQ960Lu8uTuqQCIMDhMSEP5NCAG1v/sSHK4T8Gf7pj7AGyJfxayyhqwtWt+q
bNhLwjtTn9sdqj9+cZmp/nwBsRX8Ja1w0tibnnEQASU2snpPtbxEW0XYR0c6SBbLLdXuWar0/Vyw
tmF+pzKnooZY2By3P0YJVzN8xRihLotRPuCsNGa+AzvIB+2rKft8FwLewt0vc6vn9T/9yPdf8CGD
wLA6baOpEcRei/PgOXFqWapwveYdE7ti50Goc5OCyYK6TGM5ugdo65z5aEoV2tgCjGl9sD6eIZnO
luaKwJ6+X5axkgM0Lk2PWyc/2baqtitld30AREZYeJpVPlnXm8lAqtzoeLa8fYzSBPoNouglkD4k
LtNnSODkx1Qz5XRgqx3P9/0l9AHm7gmBf/TEkkuDAH0XbZWh/5UYTssFRVwXbsrIAxt5RIjW0eXN
GkX9+tuH0Bl4/NsGtx0IIwpV+U5JwGOATns9OFzBUagXqUCFO4kMUtu4ECRUTpO9Yc2Z39jGyj0G
aEacGXcCGEZVI4Cfjnt3MxvzXZVhI5Pya+JEGuTnwbo3B7eGuAnju/TeTNfsV47qsEDaIth/78Pc
Q7KGZsLjleEpWoIlRClqEkmBI8zAf7EYq3+ylm8r2e5AWudT0Ndu3xVBmLYXnkoRnFZUuFW26RUV
TeBV1SpKfawoRkU53XCmrcaSoEaj8cmShRRvC1veQ8GKyXqB+XRs36PYL4wt58b0AuVoSEsMMbq+
b+XNuzYK5f58TV5vuZV9Aa72LuhVDeFFyZ0UODWP/dV3qZvjd8WUn/jCS2KnroZOlq7SrBgZe8RX
yz1C3gf+5bXk8tE08VgOyJi+afxS7IJ7chTuwJXTwFXOsRn+tkM56QtZZWfhg10Y3mg7HjIX/It4
S+PIrAHjSGNe0sG2CSiT/Kq+Q0wtrAKmpPkEr+sv2qirfTK3+eF5PO3OI6mwOj/x3UJMvg2Fu26h
JelrhaRYyd6LO2YBY7ZlRyQsry+mK/FKo/ktpuvZT9oFSDtm7yLHTg515lqsheA8HytabM3Z0uWA
A3YI2YtAlZLSVaQpsfxsV4Vp3d2qqdIRRwB7WcPZXbsGx0KXhvE+Qe8cztCoBnmVlnFvk3iTYQAl
9dpogOSqDL7cnwyz33WDCQNC6yRs9V0V02cnjr170jgYOxmHvNqLwVp3SD6od028iXqjazyML6Cd
i2147qW6trupuvCwMvK8ZoJ+fhbOJAc+DraU5NiAD1M6y+HNScCEgMC4nOKazQ62DhrP6+O0bmX8
gevBlEct1uYUl5ybbVN6tWlTKyMKgLE085rqZhMaoz0QGPmprzXBezmI4KKusyytwF1k4pLh2YkR
g16rEExjHXOziAU0xO9XEhvrwkB/VTgiA/JhhVMpXh4QA02aLvlelrX7EncUG2N2jS7e3hXNsoBx
fnnjErUF50R/Lxs/t5x+N0p1CF4VoTaShpKFVLsIVShrEq9BRNfd1OekjYgxEitS60hLJqLNjQBY
NbRPrgmKnoFsKEvTBYEwZoLkjPwXg6KYQDkJ+yqj7aDaaJTKF/46wU5hhnMOzQFQdRw804iWwK9G
2himUhfHsuqCdE/bESUWZv4bgOPS9cW1bjAH7f2hAZv9U5lKl+Hd7DVb/JuHDo5OelQrmdtbzB5C
MUCwrBEwhumzd9sM21uuu+oRgcfXWaDXp/nP/Z8nHEJKHPL1WONurb9fjIyr+zguyYb1JBuxjrgl
l717ICTPWOzuXdSNqv4mUsAMyXT+IYbp6FFotDbxPfDxkEJn3cHRZF/rkw8omqelhbIs7Mdgm5Eo
ffKCBb/L/vCjg2m/9vg7cDb699IR1kOKKBhGnPFenLUC2AxypxFAiSu4P7UyOmEYvA2U8NmzbeC+
xKQFImSJ5RlQy0ACD1UW6KWtrfyWus1TwdDk5IY1ckUe6/OjYVOTvau2PvORRjvo0Z1/aNANtBaR
Yi2XSpdFrhZGMAKgJsed7XDg9S89nyTeXp+dnTimqGu1gNApL5CUNJwb2DPDOqg3B3VaG8Dtvygf
ZQsDPzU02ShC2Lz0wNqwdWfGzZGOJz0QECmFoZZdqaUrLHAi/jEAYyMf4gjCEFNjjTqrcb4SlvsG
6rNZnBHfrGhXiAyal/Fd1n3VHj47U/h7CZJfPeY6cP9fehnWL/bxffR4aGoik2fkchwSWfm4vl3R
CPYotehxs+oYpMVXUzbmqE/vclZ1yIjcc/T6ZMp92AHn+Ad36xTsDicg3wmTdU/j+wmYs6/6hUW9
yz/koMKFjp8aEmkkSU3HpqB7raMTnfFhBnunXkuTKgfQ8pyRmKTV7xvH9PpDHw4bvHA2IxSggc1O
KAjcSGLGp2q2Q4jGM4T6CVkpyDqmPnnRZKBpoETpgNYLde4Esu1K2sXshduXb5PO/BL5F15VWYMR
ykPMG/zbTcZLbfOG2RVzs2gVw0EjYyFqUodx5p17Yry504KmxJx5eGuLB488z48vL/WhaOu4jSSR
UEMUKwlioFhrY2IW3NT8yL/lhRzEdkC6I9XKfV5e8vf+mx8iVkzSFmVWfHeEO2rcNIVXmcltqWE2
nPxbzIFj81EAFdg3V8i4XbhbT2n50F2/63p12CE21eZzKDDIdVesniURs4DwkqgR8uucc6LqbzFg
zlMF7x/PUYOSmK9QU5PRXGFelPxzVwHIGS1p89zm0FvkSlud1DxNquEBnHxG9HmqTpZPhQIsD0Qe
h4qugojzUElHgjkF3Ts5No+m8NjAquAbt3Z6aDLyup4cAqc1Bd61XYJIxJpcPynE2/sN2Hyjjc/E
O5O3+4SNvYyYrPSbpiFNy93s/cdseY5g6/3BBP2XRUaXAPJsq2shQkXMXTwJEzVtB+4WoyIUXu90
LCS6FIoPXcT2Ivgu18FaH9desQCbTI2sPL3vCfiPcwKKN2cagi18I3Ws2vXLl6NvIl+O42cWNOIJ
Yw4gpbwcv529gfjkbdU2Wdcjn7M19qLyenL5aSdyG+cEmtHks22gDfva7HlnISoe6y4KEL+OGeps
MfD3CDFlqZjaVN8Og0B2pHqx3NUU71cVIti3wLpnVC8cwos5wwUXoWHkxdUfycWf4vSt6xltrwiB
NJOO7PygRqXSSUcNCilj6Lx9GDHLid/OSN1/HzxcPd2kEkQauHw1HLZh//03oMgDXAcRQt6O27YR
kX6Qxl9U5awaa+O5aiBxG/oakDl8hED2ohuDGH9FyhrG8C4kupTdwQWSIIJUjO8KLeSIfh0Glumv
7NiN7rLYGlwdjdDgBpK+MdLQ22HrkNCosgYNAj4TFtENnWuupbiRdwo0sZrfePVaoIJNGJ9zTif2
xUprZBCRjqEUdX8xq/Y99lq5ocdCo6wp50CWvZbsPT39zPVLUNIx2UsMN9e+ip7zOD8dYDir+x/T
dauefJbuDAjNptbtOmJWibIA/SKaKv80sQFiLUEik6p9FuT8cByUjOfgAWb/h1WcbVic/jSkAoZC
1HaIv1wUbuELZwxaZgRr7r5rSjeww7Q9F8DWn3m1lmE92YOQIv95qSpFvL9Sg4VLICc7I8JHhLqY
KhUf7HzxyU+aPi706fxqvii3lFf1cFM9IP3+J+xjH1NHrMnGZDqIYkPp/P7XMrZYNTUD8KiqmtVy
Dlh8KmigifnJX05oo8rL02GE88qwqN+yL4MGCOIDICb+7maElSUnPAoax9au90sb4LVooktxlk4m
GfRbz+6uoRUR00mE8ZhdWD6jYt3gAgqvy3mNqtRlmawAYp4XF5yQeFhMzUW78D5wOf8DYxuz0hew
jWhUUbcJfMcAEwFAFT5l20/YOwxYL3jqWKVGz52DRa2akdutKQYd7kHJHniP1YO/V0Nr1jsR3A0m
TGx8J8AVqLJjtHPSXaasx1vJKiqKCahTmE3GlEQ2mzyKnVij7wG6sVevGiAVzR0NKNUa7XePaCxE
bXouEAtx/9XJUKkrPj1EtUww3tTRR0ij6GGrdfuVyy/ZkTTdfpkP6ItsoWDVpIbLrPXOEhdnKZtD
gs4O/tYFYJ19lNoKRkH/7BGduu6CKE76evUUSG6bx8gczC97o1jDfQEOLk6Cfd6muNbkBwZm/yF/
SHSyonGlSCy4YH8ok1Lh76eXdA5IPi5rWmWk1yE+gd+BEGJhLPEK85qsUCMVXKCkJeEe5il/LxXk
SaY/wPxZuR8go6RcOYE+ybdgYg/g4NoZcj8l8sRb43OW7Mg+CUCpMugzluUnBQZ+OF7mjVB+MvwD
erYrLZrZr/D74FgY2pjIdXME6ZzV8EbweLbcuujw6qw0h00injqJjVBvmHgIcj12canm/EtZ89r7
fMb9P3kzROQ2Bfy1VFSIZ6i4yFz6hy499XdjzQ1+H0dNyhDzljcrr7h4c1U6gPO056IpVsJPmZpn
fSBg20GSL+a4t7Ed3meUq8sV0dBaCdDnT4+Q0FTo4ieUExZGvANCsZWaxDkrTWG0zXVmnK2ePG3y
Z4glvt+tre2hDEFLuOH62dG90aL9OuIy/60qtwC32Icj/062ZBgCymFETwzEVN5DnWtIaluKlOck
9D+8iGo/pvD862L8z/8ZIx2G5XYD5fH1MGGyxi+PFCS5isGGeHC/PnNOvPH2G0HYvoN/nHkdKGXv
X+NAz71pywoywiJkWtUzzJBKlEuOyuZJQ1bEnnh0PzMymBRj+IKddCpli31fyMVawlyLhZj10ABC
Z0pmHDcoXrwNs5JDyV7juA8WuSrsXb9GC41TM3JIxkM5F/Tkrf0mI10MVCAizrVYzu9ijRwb7cfU
iku3p7OP/nCDJNFyx0Jom/60B1kbz83Svkcp2q6b752WCs1UGKQuehrcKiRiQLI7xv8FveP9YVuw
Jp+QFqzKuMLTprVP/WY9wGxoBT51f/LzrPLnTkhEwqMNIbRvbVF4vbzLwRGWUWrByGuGVZwTWtqd
3dq3nQO5zAEvsiv2fGkLPwjiXMYBUirXg3IczE4eRNdjHUStkfp0Bc1bhWgfBNxTwfG/1VQGYHfE
VjfLysqHc1KA2W1vsU8naBDG9zboaQ4XEwidlwFXOohkxu0dDmqLIcHg55NAFZ8nvch4Y/SnI610
oeKSLQzCt2c9+Q1qUBI496ch7R+WUvlIDwAx0quoCf5kl+KxMeftwugo/7PuEcFRytbTAXgnVnG4
eNpuT9GoqJZqXF4TnEUNIv47Qp1DAQWV0CfHn8YgyLBcag8bYtCf/c8qDFknC5xDsHC1hQq/hYLy
I0J6BA6fy7kbom3Y0uzxaOsDnIIOe3up4AgF9qN49morsce3JK4EyT3g0TfztkY+XBGuPETatHgg
Qvnctu4HXTsPB6EK6yjO/sM707JJnjyli0YQfA3006zRcLAWJGnZzIYkWtQQFpfIp36VzTuLlowi
8AwaV/YhbG/tG1HbPlMfZvyDmU3QgxABAj65LtxZgZYHin1Uw3OX7z9qaWbZI6NyUUJZGBfDVHiq
cQZGVI0QPDbYNKE/Ok/t/74FQ3XRbSJ8SdVHtaezB+p7g/3Ti5B7BWu+5eagAkEoy6X1UBW+t5kW
R4YoIa5oTZFbvCNYb1goYoPXcydYvJQiQmUlwTClZo3pUopiDjmtR3tq/GrYLDY0FhqwKjQwmryw
9ojrFw0rZ/oq2Py3B8gBrtXnTlhqzZ56mLHQjncOOXbAvJcJBDThizEKItSExvt7+xkNSZU5pRs9
Ksoo5MJDWJk1mq3+3kYccUa3E/L15nL0vwhDFf1HRE5lKu4ySpi6dd0HOntz8UFhRqUdA0a+jnoy
Y98YAveJf9NW/PV7m4pDc5vhg/hbPATvrpnue569hoi//CbJa1aAbOCFZqwqIC9xgOETxD3ayBub
68xNPUjNmqAY8YSGRyiKPV/yT5qzlY/jsRfHB+JslyZ8UAAqIOZs7hl6b8lqm7dIDA5/BsRPC0+q
PLEMJAGRk7UtAphLaddt3rUY4bH4+e9cbkAQlzsKqf0dkDrukJ/gnDEOwKxSkcz4NlA7+ULUzvqA
U9mlMLmPbs5A/lewA0I8MjXfMd20ejdqmlqnYhU/n1tJvO4wGtJCpBsi+wfU77X8nlMNvtL9rjOj
0X19cCx1SXhV+vdAowFTlRh2pJUFT7zW/gB8UCmUd6UL7NSwfO3eab4hB8HFxOplyWBz1xG3jjbC
cyOj9wwJUoYl/O0yGz1eIo0ctgllTtYPq3ClCP5f+f2ec+2JWgGchuIFh7t0rqTvkRkwCGlTIj48
/XdUtRomyyMaYhW8PFpED51RdfdMrhsAV7N8dw16vc8krf9+h9MaHf0w9fXOtsh71t8HCSszQqCR
wxaLDPB1bE89eC6DrJMlyyeQboy9fe6yLbLh5y7mt7JTIge1f2edQptukmAY6Z/q3cvf8R1Rdq9n
RPGIEtXbffkNU5BnFT7+kFbPIrmQO8FatquEsWbwufERlvixDvj756NQq03VghHyL+ibr/+jvFxy
eZy4Z2bzWSr9Na0WFN5LaaCZmlB1BsspUcbNSHfxIHJY6Kv+pMgRzF1GTejZhGmicX1vTPbtcznf
5kg1hCIK8tSnhulDu+Y4JbH1lAZaQh+TrZwzlUEEom6n6fB9sRg9GG4iUF7RvJX3/1vSSVqkaEd0
CLupyaxm84YmXIgfo1UrA7RHIYjb8gZ22kNUjg37Fjubc1lNCK3hYJhbvs9dgqre918X9lEjcL/m
gYrcgtAn9fr+v0AZi24rLNVLzXfMZfRv/g42w5nCrbAOnD3U3aN4CyBDa1QjRj5M7GosbJ4XqZwn
vC9A8wkjByMONuCD7tNvowD1CxKxt62OGz9DIs5hVfDHzqkWOihfXUmyDtfG5UAIY6cjaRAm9c06
WYxz4S4T2dDe2hljegU9iNlnk+JOOp1jK3ctXzP/shiZ4bXmX7ppDbbE1JnknAdh9rEgcURed7E/
N36xVizBMGvf0eWeGb8bAbYl2zkhhfneGJwuErEOQb85tIkhys40dvM4nV/icXZhxvc8NoTSp7+I
0kN4nWLwNXLPPFwfr8nLflFSHYgVBuH1BuwwlAthNoN9wJL4L0/hjymn4AnorXkjtb+sLaQuvOYX
sFf+be5W+TELTjYgkom79RvF3kSia9Fvn2g3qKihgRwmHqnaIMKybxaHV065KrUhpkxpWQmwop+F
kitCOwBynQ0gVQn/f2utnIzC7WGYIhBgSSScX+TNItrcappDmsnkIOJpOqKAuoi1SdF1s6Ei19S5
jCLMBzO8SrQoP0WxR2cXe1WgnnPB+wOyYKRTVVwIsZOTDj1qN6WrYJedzr6N6brQOCYcXoTEYYun
r1cZmxgCtVRvCggMojcAvRh/PBR/RXcn4hZojNG9fsXHN7jD1AuRnpjbjYWV+JlKogunk9UWo5bO
5rZWIuoH0osY42NW0ZPP43DIgzkPdk92gGuwj4QdRx4+zXXUYcEka71kJjCQelh5JvowsgkMX2nL
Fpu+xIM8aEA1RnlTA6vsah58Pkn9qy0zuJ9zfcikbptF84pFvOMasteal7/P/lvbE5FVE90GJHlI
y+vB9hn4XQasj3J3nEK38RLWPWOus0Ji6sYbz2PB4vLXTKuXVYQk7NHaZb7D9GRFX2F9sfVKKddO
9cOTW4yUc8tTMzYtNL1ERyS1idxXVsFc7spUdqXx0fJW3O5sFA8nELH57dFbk8NdQCBThokex1jk
TyMddVP7mCu+1xLiJgisLtdKtD/clayFSxPxPcEuJHzaNmadCNpSFLvc4liRDSPvfju6pJVc2Ao1
Cxe+Sygzh/JEMcApCu+dcYsAW+8zgeub0STs2YxGA9Hg5WI8p7dJ45lMNi/mAVoUwo/7LMVKv40h
rLtC8hnYe6+/cY77UskropRmS76y31lQ7OpTAOwziSunmC35NMnrD9zeWgo0r9a4wCEjOr84Oe0k
Xcl6W/O4Syx7iauduTBt08LrmIXbcILfTwZDYrpjao9AtgSk0OwB83bnLEIYN7v7f8mqHyQA4VVs
ATkDVpxVssQa2lo7fOrIDrtT94DGATQKHBCpaUtZn6gIsUa5V4lJwNVP5z6Ak/375pAqeUxRbEev
5B3dCKmmHFHRLelisIhF51+MqpHPf1lrXOIt+UOn5dt5KWdzqeIWtoyr6cpxO5z/WWqwXBE8h/OO
3sHHO0IpCNr69xu5kv8L1ZBATDVIFpOs7lC78oJ1h63fIf71oRmkbTgDeLs3yVpb201NMIUK35n4
1egjZCdpev+H5jxZiWm+1GoAvLal/QBihH4VUQ3yQUUB7yqX0Vi5hF5mTU2QInJ3mBpmoCck4ONN
pp+KL3CUcrY8gH/8fs586LO0WTFl6CFuwS6GpNH3HTxbV3lluCDneBwEaYCmtw1XN3vbX+l8ykDp
nGWtJ3IBDnFqJuqlASqO0NoKaBPhVTHzGV6N9eC5ucijKh4UnsUeCsWZxTBQ99tOpQvuXngRVJQ4
MESOQbHa1zRrudPgkuyWZdY4jImntJOtnDvs5nm8PlrM2cwdHhm89GFmYWgNYFqZ2oSVSiRmyjCo
7T/Zs7u/Dw45VB8MkmpdsfyUG760zCrXjCouS47px1mP/Xj0PyVY5K4+kaVdo4M62t0GPR6a65lf
Zr87P9uOvHBYSSqHFwyU8rvniB+RJy2gcndQWSFpbu27j0jn/g1W+pyLVp+V82Il7w17eMkLJExJ
yfwVU3hFV7r6Qc/GSehGTLb4LFkm+v1d06CyyX5VyQqowQLKgwpGy0NbOIwYhcLetuzkqgCABDiN
fCcx8x35bYHGRqnpTHRJAp5ns81MsFt+7YodrViCXf2gVnLJhCaztqmsVtE/d8+PMLzvlVOZRc5m
NecIua8/E2hZAVgFaQIOdO7bm16+cYiuZ4mclJSVotaerQEtyIe9AYrEKyJcxxGPvU01oGtwcoJU
VqimLjVpEVutTwoWxpm6XdfBoT/ngqkHp5mvjjCrPTX5hFpayVd7dEtJAeBGyOcvbM2BckBJhUmH
EHSVbj42m4ryIg9yMAIB/JbauobeKiupwnrf3wtQN28Zf47imLRT4Jf1YJj2MoWVuFHESy6vWjkG
L07Fw+aNKVQ374+N89REc3ghsQtwT4VgqXKI5H9rvYAqWaMtsnpewulLf7vSJ9kgR9iz4wEEcIct
6dJOQwiMonMaXY3wryHR8frJiPIdVNsePGPjVqnxBQnR8IYKvv4rPBdykuVHcARm8dKabZqnlRc9
gXtRQQ4nCf46Ghw02vJJm6qY52CmVUVh6Pcm4iPVG3slXrKtiNdm4fQUQMN2Zx0RBW97hUS4a9Ka
C70x4bZcBCIJ5SXfM6YpNTwsdDndTbgykzvHZb2a8oY2VvLtSgnOHF70fBnHjGOEJHYe41wCi+nw
v1cLSenC8VYjKy3h2HuiwWR/XZqgPPWF/m4R7Dp79XR5KMM5ejVcjXF8rl4/qwvBKfUDz/D7yBJZ
dAa1uqlQaWjX7HzjU+uro8D0E8t3wnZT6nuphDbf7r7bTR8xJ76Y2gbPjSqcA4ZZAn7iEl8ToLKI
HaCS/MPn87O2+uiyUYM5phpsdRavyxWPEoc0mYRkF3RXSUjgZST+AEjq/iq4rFedda4X/OWOVCJI
+VcUDu8xpBEgL582njNDgdVRl7Jl6F1wr7Z4IkxLcOilimvA6QvpaMJssHNVBfNvFxfRN5jItqKE
RSubDZLI++OSYGQYE0Bp+5+9V/qZXmINehFBdLLAmmaONwlLdsMmxBkfGYnNFVCb+rs0iLJaUQm+
XrQhEMYWtSPXKw1BqgFS7owZYtNMpC3t/vE8LtoTILU8V2cNoaB9kgVg39qSpQ3+aLx9NTWw+I3/
W1gXnMLkf7Zp+MTjBl80sXZZ0wJTXCLeQ8/N2bB0VhppzwGIfZBopjiI9PB+L2sX6fUZZtwQNq4k
oCgxNE1k4Fmc1PlG0Y9CfxhZIan1obAbgtm77YQepTMS8Z1NZjIBUvfsq6a+fCsfPDeANmeuP6TD
9MM1D6eZc0ffPURCYdk7CPoAwkPcu9i9DhHlhejVPtxiBT+CUxCs5rrwlAKncJxcWn9pXHX9xGsg
2/bG0EMXsYdb373kFyG+lSKci1xFqy7VQqgEfx4gY5S4sAxOJLnSYF8uYL6HsfJCds0kFd8DIPHw
+EqONIX0rYz6cUsR6iM4yAAxBEp8Yd9Q2noJJej4A1BAcoFfuXHrFU8pqoojWHm5EPhxYddYDUW3
GL20W9O81CZDQmA+U/HBn+7vfb5oAvLM/LHfk4l6Q56z7THwnPvq0NEu7HCyd83nnsMz6FujWLeJ
XtCTOvOVCJyW6BhNinSm30h7VOahu0MgNSDCjVSL+CWPhmxxXPY2WPc4uoY1OrWSb92/BJuECSEf
OVYDQwn7nyxpLJSjdDrz/uxBEfkgRIyc/vyO2+UB9g368rgQtLlC5hxkOUCkYHLCljdxWOA4Goml
GddHalHanMsq3npdsRu3i0R8Zd72uqyzdcBYa3Z/vRDiugJjmdvMoe9aphxD9d27RYfFeCHdIUJa
b2+rbbNelDHpO/8irxhMC67XOZXPRkqgR1+8vllBaU4e61BWiX02i+au9mNjx3EQr2Z0BFb/k3q1
Kz8PQjjTghv+59shzzDxCWhOfRUFLAkbqNtkv0a5I27uFuF+jCdOm81EeYoomA7vqsLhrzXekZbD
Rm1s2aQTSxsB10hQEAq2j6g910w7FwznUnPuMrOyz1kED5s20Uq7cYGeqO7lN0g9LeJlkAKmqtE/
O4koT1u0khMCWb4h3IXyLHagdZlxPv/dpF4/kPKrVR4wszikloPiXaARzOrXQ5EIUfxIspdQ3rDM
FHtq7YnCMQLEF8GGz8yb49kTTEHJSnblqD0MuXS3mBTLc7WiQpkIshalDmZAanOiEsD/TxKTFhJd
k0JB4mWEYeNh+78CXhvKJkFu1LrKw3vvjOHa8xZ1w2Fjq+lFX9rZi0SqRuezbP0FZ26eQfjOWaB/
coSrbSS5hGRzUCgxAGWnSJ8aQA4URSt32W9IxZ8935QCb0NDeJXb2p9+iSEJnVJB9IAzBPE33aFN
h6OursFI8nnhB65+aPdpTXTmZ8YTJhyj/O4kMPaNARlv9isMM5QZt+OXfJkyz/dV4qVMgzN4qhVB
nsWJOpB0J+KMqofLFoZ78dr7A0jZ0Vds8k7qVDtv1ElsnwnaNmjk2t5IqVgZ+f/Q+dKhPGEbUQSV
8zNLzheSTA4iz+uCBBMI/ruPq7VpM7dLcJEhknsc6Jc4SiRBUr7Eeju0anu6fJbENWSdDD1l4vkQ
YeR4xZulEjbWF3GagZw8bo/XHOCrNyS1FSVLmvPqu3nGK88jBhEgF102kDQhKjOolcbjBg85cD6T
vfxd7Tw1pT+veWY63bWu9kM4QVPj40MaZUIicK/9dPJYExyMVD8FkUbmPNd5z4hDfEcvSrA28sLf
b3cPjsde9nmNPNWXQCskM9ZBh98sKetFavusF8qtecKMEm2DjBAnCatzAN9cHv4ujdQrZ6suMy9F
5GI4Qg8yzi81HCsVrXFesU+CXFWzxPl+ZWM9bQT2K55+50k3H8VQBo6dqxujcWsWWAtvaySuuVIy
yyel1pIDnAvC0M/zPMMiHg0yX4wM8xnKuj5V+ltfnqJSMKkG7hgg4CPSys6Ma+5h/0KKw90EIuLk
ec02hzmLM2ubRt2h47yBBoeQanO19pNrDSBTXQTKRnmqYmXIcYJZObBoOnQOYWmNyGMCrCPxLjKN
iseBecHrbNUc2dFHEnX951OoqiHIhXz8JgYFL+jbPbWDpAFUxu8QnccDD6Q1SaCmmmuYXmUUO+Qp
Aw1nEVW2uigcWKOU+k+kgNpPdVkuPBQfRib6qVYq5P9FyIqu2XH12va6OqyYidj7Bj1kVA46JkV+
Yz4aNwIAE+KFPdVb8XL8pz/Wx/Ym01Kl3FoNsmHNAJ1wNajzGeVUFfOJ4rAjEMZSbDpa5CQ0wMRF
F3kqXItAlTu/u2po2V36+rZk3AJIoS/yGHheVs/xU6ZUnz0Z4AYr0RpTtOLNin1Re14jpPfOVSyy
Ka9zTJ9fMGzchUgg1va6d8/x+WQ8ZW3d+Bhl7t0rWDtWz1VKrclhR1WvcURquykf1uxRwz3ZJMjJ
1bIFI3c53A2i+qCn9jONKeLqCXUASc0lihY9RGU3VOkAL3+L4Ee4GxNSyVovijFlwGzKzU1nUD/7
KGi9YMSoZCrosogPWbkwrDmdWrp9AIRJbRpxSNFPKTrdwPBLNY1zlO35WKNlGvrMnh+YSNanrHc7
q0F68lbDMNl3RetcoWSQxJPnFKNqI2Ch7QxHolxIRr1EUsBSiOIp0yTSZNhS1NBlP0sADW7Z/37V
Bv7/EHRPUxRvWJszkxurK0q6tzhve4/De2Vou0swbxJ/fOfnR/xzWnC3WKt1Jh2JyV2UH/II3TI+
CmoN1K5s0lTjDbpfYbLkrlVlpoUxPXteymYeHFryG+zuH6XFF74k9Rmwd7Myzwgeas/0N8wcueJR
lU/7TN0Nu5zhfWJfygYGyJVstNoNZuLPx27iiCCEX+hjHJ9TKc6Tjea8imHalIacxrpKhrglvPH3
hyqhzWqTXY2TsAACm8N+2V+yFogN6OgZFP33oyGRKhRk9yCq51ejUgAViQGC0ldE1UGaUEioboMi
08NUC7tTkdaqBdHvVJyaRPjqqSKxpPIsNQlARXqwO1Ekmva9os1ajrEAGUxIVDMGNmpeniHiUyJ5
GMABIXTPdV+LeW39D6vW987UtTG91o5BZ5ji+WBCVThYGTBC5b7UabfidHKNv/POXP6Wp4kTiQBA
8PvCk1m5E9qNGuq8RMG9efXEy7RzSjyFxDa5RxA0lfPOEGtxvAjqbWTBzXmCSG7GQ8djNU91QMce
7N0Z9c2ziaDRqutXDO6NU4TmR8CpGfKJb0lEmpG9oYBkZoYGBQosmSs13RwBnUogVcYxcsWmAZtj
EUGH0lAK7+8vPJBRo0BBVN3sKsGzRi/WP9wdw5VOl+1m52/m/OEKqdzyEVBvsR/jTG1Cl7wI94dC
tJsZsshnQIPKDI89wISl1JhjutFlZp9jv7Ebb9EjtgqP3CDWm7eqUzcnJVyUzpJAWx3PQhSTYY4y
yZ/K1X0AexdsnyWgMrHcBz3m/gSuelLnTjzEFOW60K3/ICurSwTvX3WtpbunGSb+3vq8gkhAb694
4siN5Nk4M51CEypZFmnDfYbx+Lf65MrZGDEqKZIxpowP+5a4zdGThrHXFX0YYNdIuMuct4HBaROU
USX+lTYeF4X2qS+StJzXNN//mgX5PVblOKWlTPU/H/Cm6PuiSh3D11I3USZtuV9fS3vndAutQL7x
M/AAcx737giMcb8YaJqsMDAfqV5u0jazVKy4+NW2KiS3E+8DvoyYwgGvL4AAt0/uDhbAaJi1w4fL
r7raBi14k1DPkun/7jYlXjWBvoNLTtX5+yukbS0Ar4oiyd9rHMgpr9e0CHOn1LJm2VhU2Y+uyxai
Y8dwbIHIuhQgKy0pCNEOvKPXCs8+G15YuwcJw042GwkLBagjuG+PYCtmFz/pmzvM1qJgKDnhdmpl
AwNSZa7xJRCP/ngn12KAqECHpCzEjpf+jCChRmV91VcBlfF5Xpl/ciNqCQue5Rh2gk0AG34mv8+J
2b+IqrzM2LDd6O3WrHTW0o6pUp8SJYaEJPcOQW+y4UiywkAFEILnMc4WQ3I2FBT68Qe6mwOB6+bH
vrPo6yhtzJ0UXXz9ZKPM0HeOk7JM9I2DYh++E9687fms9l9+c4GGxLR13UEY2SdQi8HCueg0VWob
RUOHBBydveoPmSUCL8T8KYqGvcjAI8HzxoNkEqNzgpJSoC/M/l7wH66QsQapL9p2FsvK0S9IJL7f
VRkCheDR3vwmNcroY6UJQsatBzpo2WY0DaSWh4Cd1gkqFbMbJql6eJ/ccSYSSTpC5+paTXnGLyWx
u2W2weuhDtkdnGpOMa4sjC5SLPbm5yqMzLsdy7fw154kCd2EZHf+OaW6Esh5jPWMTJ+rysmDFLWy
tMDIGTpETF7OTe/016eWzy1w/u7iHJ6XBAf8x9+iN1bUt6/zroFOa2sKAtpFi+kpNsuhLEJg4aFY
qhC/9rWECZ+GZbQeorqIodF90MjEYS6/CodeaG94Jc6dwNk3JKtvsLfydtqRP3OB26cp8OEdqt3n
yY4TXFx8m6ReFFh7QeVHh/5IFGdY9o3+2SW3iscPUjX9kvVWyUKymYsp3rd6lmeSTL+ZJ06ZcGV5
8KVvDgfB9wJj4G5KP9HqoRCVFsdwNDSCLOfbObEday3NdiYQb4wru2bnBhABTc3phELrf1lzlR23
KIKK3NJAEAXZbHk5KwLHMaGEqmIZdJGClDETs0zWJQyGhzzelDQXlH8dNmUdA2VOqR1vdd7NC5ru
AGoQl9t/lj1B26uPywoQ/a4JGl7Stz3gCAb95ATTgCrpE1WWRfYqCu2PoIFuQWGU5nuVW7vFwIBA
oPGNV7DuS1NXiDbjTx6TKMWMrqH6aDRzxSVlhWwT7Sib5ogsKMhJ4YVcFCSl1EVnq5QoR1nbV71L
NwzV0IdI2cKh3R1kE9rLrRg8mWhytrw3wdud/OlKPZx0yUUpOGXeL9q4uNEZUoRJjzJD28QyJPnS
yh3e7uI68EwZwLP2ZtwKA0XyLozHvCIg2KkHirqM09ICXSXJp/Hc6OgPxAbPBZlXMjt+iRBKLm54
FcYmLrMrxj1oRWXDmWVRHiK5JoTmVEnwZkuHX9aYD/3A1+EPOObBdcZ8OWfedhLXXtmVdW11+rf+
r4zkm3qRfKdrRABaEa8wMYKIcPaLLQUaLJI4wmfqvHq+a9n3MzuqJr1pBdQEoQ7gdg9b7FA2Hinc
zrwYcRUhgBfiFM7MrRL3MvoKfNfhhqISLFVaXhra8wrI1K8nTnJ8IyS8GdctS8uVtx3ncfWlvzRN
Qz1lUjYQSpJdVNoCJfTTnRYp9UeHPbThpP4H3DdmAgIwmAv2sdsBd/qOU0laUmfX+ruVi2XXxl21
T8FFlVgoC6pMqyReRat0NPefiVngJG9Y9dSDJZvgZVsgb+5sjNC71vA1agL3eQXZq6HQDfoByPmm
x7vGnGrRXQCZyAuUNJjXa6Sz/enlzQBGcvlOJmr5oxo+2T8/XiJo7jvonLLXpyNWIRQUpHK0O4bD
lEYhPDmmFDrj3GDJcRqMEMZjrXttDhVmYrMlLbnVahXiiBZAPXYRUiqkSz60Qvt++AM3PcyodoQK
2zo6mkup3NZUoPDNKa2CwPz6RQIwyq5eQ+C4LSHNxp4++C20InFLsyvoOuCa954weoxDKM9VGJUa
wTllLXw6Wd3TkLJ40AtIJgcXu6SiLfdFc/KyxCmr7FjBbnLAJwZjQxZohvgGjBhZJMd3iFE8HUQL
ddCy5PumQl0Y22cAfeww3fwZ4oDWBDLr48iE/UUn9MdnsCy1iNOvK/AV5rNn/0h6e7Or5v1vSO3s
A5PWw61kXAasqwxRZ2z7fjQgeU3YqMUF9mvvHzbkUvGX54Tlne+1uMeH9VSwb8kq+RJju5fLdwlk
SFsynmrkqXXhI3lsi7WTf2RplmIiH9vpo8DiQM84cuPkkGpwfm75xaWYGSaVccPPQT/SiUaHDhsk
rM12nTOx11QzFSiNbuHOh4HACylmjLyycfiFyceZUn/GJ7ZmYbGpwsSe7aq3dqBd9ofRgIO24dXh
GQXrz5xgrttDp3ygFiWl6s96fhsRUQ0Ftopwu9CH5Rye7HmZTcwB/t+iR4gpgnOUpWD6iUUumxvo
WFT37XHU7XD3a/N1eu5rrTBOB/2wiECmjecWqIb8HM7vCTAk2ZUkKQvX0sgX181wc4Wwi3AKyVxG
8RTNAUKs5tv/HjUdqnZavqkSLGh1S491ni7UrNiO9P458vBFNzPf4Cmu32GLR2HuTZRLPSB6EbHY
/BhhCnDKDdvCkTNeG4qxPkTSUFllykbUIzC294IOFerC2GLuhJqqzLaszvaGjltCcXEyqQo8/A0t
rZMzNuAxj+MtcyteAbUOjI9zJOa4lVO2H+JwnsBFbTUpyIZbcJWRuoMJDC6dfd+B0b4BfQw6Hnvx
gV4nG3Yt29I0794fRXg8O27FbD3XXC3GTDxe6Nybqa2kRgfPXTzets263exiw80ejcWfWx0pB8bM
6kj/5eagKPskXIG/0CvbcphyqIH7oT9vqb3jZmPFcdCxzRRIL7HfLOulMPiNjQGf2jU9D67YLBg0
Jtm0TjT2TMLfgRFImVZ1se203ep0xIby6N3Ft0/E6tTKpQR4ZH3aWczPulyyavlmWTuBqmtLBiSx
DR+Ccj+OrxRVvD+ojmivImmAR6P5K2xlOIgUgWXm6rY8kB4elGGXnCnwpvaHkSQMy7zfbW9xpzEo
6kgZUnRar+XDXONgS2zfGl4QJdzQvdQXh4mJ8GbeiTUCyJR4pR0eVMoGhzf0Af01OK31e4yK80Kw
wGpXG1+JoXpN3Ec8mdQurP0aX3NCAwjsMf7kG5/I0X/gKgBxX3xN9B3j66k1qJwgs+FuuopauW/z
SAP9wiT3jTd2dZN5NZg3pCwn7mmewnRBbH1FC96cIFwN807vRrNSk8aBp9Ys9pQSpL1gWaNt6DWB
LKNjhF46zFmZqGbXIbdx3gI53BLFRlKWB9IefpaCkZS7ztoi1JZAjGY/X0vYqyAytsFMxaRKUSb7
QWOIjXP+jIYwZMTO//gNIHZXORurAl3RQ58bKBFVrXFXVoyL0fXHULpa3iq5PrrTjyKcAsFvgEdu
ykSgxmtYW1Ar5BgUTT7GcewXUGQqWyOyup/5spH1KTQPeZ4LTbo8Gus8HIJrEHMibod2VspxdzK0
85zlQxOrwkk3dkwNQOZArlO3fmC3l0sJf2bACMp8JcMDlbFz/u82fm1gYjB0H00BocYh+TK1FmOA
MgbPWKSKMVv5DOnwhaXQbWjKiyPQOlTDmHmFXpA3xWb2SoBSILQMcIEItTiqDpOmXS2WljyhWbk7
RCcqJG+gGbUAlGiT8BYj9vaUjTNxs+rphyqEVyGdK5Qs7ZlyZBWG6k0Ca3yd1lIo5VQ/gSx1u/B1
p63KQU2IbLmS8NQKxFl2e7hVnxiu7ZoTk6mSd44KVYWQ68Fbo/KVLIdMT/+Nr9/sy4/7wUrd9dcG
qFgNdbeaaB4M6NIKgAN45PWoUXzCFM4lwupBvC950s1hqZXHKUQJhjIE6vMTpf1h6rUoIxnTUt0W
pSJ6zPCb2yWD7C1vm1PeEV+upFik7V6JEPcAqC1Ep/Z7shTotYM7ku73PQolef69hx1IFFswxFAd
SCKNNBpO2vwid2JqtxUYXYKERZrWs8yHC9JDTFR/IeGoRGAAfTeLU1SgcALMPSI1BWkkJVyYEP6L
nYliLbn41UHqYGqZpbP9qkWILJ/xS9DSwB9zP91onJuDy33QCbjMuDhGZ6zdZMDr6HDI++p2qu7e
c5a9abGi9EomMzAYNp7QNCtwGXsvoAbS0a4gwOc5UjmrtiSvCVdgqxo0vYrjcjo6KYUZwDJYhuiu
DyB1szn18Zi6ccWnm5f1bAGZRQsjdZOJLdSI6V3yiQ0mz7Nw/u9+ONpDPUnUs0Ix35soS1QQQrr4
YAJctcCrOqjujXPOgwC59w8As43tfyJGEPu+ssRsOdE3YEGc7XQCnXBtcvPvULkHdGH0rkYhC2lj
T6FO1UsuTlGQFoYnZNn2HwvikqlOwOQlDVp73ozzSoVCQCqUxrw2BffXINUKPaMq3zZJWgbcGW+o
QsAYjkZlp5ojwMR0ruY0PcNwopwZhv2OHBdCSTdIvhapPjW3ufRpmgyhgiXjFV4Wr1mk8JUCgDXG
5w7RYy53I3dbCG4SF6ey9+gbWLhktXelg4dNNNx1luhpJzdWcNo+6tK4lt75pa0x2rcL/3/a8MlE
3uyWM6NoP2/v2LdIUb4eS97cvm4m2HQHg0Dv2nkE/7PxnZEUx8T7dU668T8a6mxGJ3XBzmOezVDr
OMfe5ANRWNwcCcRybKKV8a10gAC0tA0homY92ojp8FwVNNCDnp0IQZhnAVT91BXHq5t0KxKfjMrh
fH7YTCS6GYzS1xXVjF1QkiIOCeGXYsiEKLd3EIpEqjwtuaUxaFQsT+pqDw0y2FHbCbrRy/RQXIRl
Fy0E6sPtxUI7je3GrootXrE1K1E7/sgizQUkFEpDyQRaXPrT2MOxHCJ+xR87vm+Xf1iqfCvumLtG
6v5tHhAbQSKAnSYCU80kOLHyDt6vI/SaqzTrrvVXHt8Y4GizuUOCOTeK+hK5lo6KRA+PYZyOdYdn
pe3lHLepK4+7sonAumtSSomvG0bmo07UI1vAfghAAK9XnntD9Z4Zq1/T5u4D5+QMgLexNyaJEwmA
gCcF/1l1MzkcydYewGzRtT43usdF1syUFPY3VdJhMfsjIBCB9pRbUGPpMLO20pipH7fcFD1jfqvA
g3CDeEHS60duV50hqJ2oJB+ITG6g+2pwD8AbVQGEfzUPEWkCoHM3Uu8xo1zWfSOtOGwwv2iTXqo4
bn4BMzK+K2ABwJgW7MAj+Iour4c3D+bt1WVKVDl/pobuJp5Z2SGWXwPa0KoMmdH0bbW3+pJOYX1e
g4CtEJ7q9aIs5Xi0KKlFx+EKZPogG3bR6Cvb4YRlb2VhdK5ucBXViFc483qMn0KonzT3QQgHfpV2
2uKEXVk/iGKt2X+qXxMYByqHAKFWK50Y4AaDvDJhEqXuoriiH6We/N3YtBLEnFml5eqD+vvBFZYG
Q8RfDMnz6wCYx8LGf09AEADHDKqjrof5ZvYIXFSLNGf0CXSVbTOXG//DQAtveDnDbGZ3DWGcAj3M
7jXvnCieKEZpiNNoJoeFOjoJH5SF4pEV/zXES2wqMTQ9IbscT3yyJwtDwec6Abi1jgpyPlM5u/4Q
cKjUKhqtexuiSs+u8OalGEZykml9Ms4YMEPx3H+1iG6wamhP5YGMlKJhRzelGE9kXKkMM701/F8z
q5vlrygiJwJq29K5DaYHxlBdCaqfBAW5FhsVIeloMCqrEUXdHkyT/N3Ryafuzq7VkoV1xA4NeXiO
94IvmHY4TDGS2TzEdVDsr4dIjm+8yzO8yeRZFJDC/L+hF68oSccv5R59cG9iJfsOjhPzgcdXxh+r
wbRwyrgrJ5wYfrlm1mfSXSXHS/Z0wWD0DrlTd372yiAEf8WB82q6eMUOmWi0qiaroFDBe/WxBi2p
1I3wfk8MFV9jNgZZODxfPigoNBvEoMrrEx5dkuGseSg+dRTt1piv6qQTz1RAQvknEqHPyk9iFe8I
dDiNwDaT53LgE61gn12K70tkOVTNcfmI58/ot04FRzLDgPyyjSERzaLlltLAf8ifgUX+EBuKe1g5
UCeAclY20FLY2CBcfKdS3NI+sD7p/I1J3OxTFkZXFevdRFswq4j/xXrnZlP8rFMat/Pme+LUh+0z
tRhHckPbKnCQx+HHsWcaRWszXD5rmC5RPkDMiWis1w5ZIKFNcUOrEJZf1uUUcgNrW86UPNBeRKhh
SgjNzyLTmzml5KtGrZpLO7EP8msV2uG0k7gEWzWz/I3g2EWbxYWo79EJ5Rp6yq5GLuJyGBqrxTFA
k1fg3ptaFFlQ0R0fw8nLtZefABrHNTO8cI8Op6xVZSVpkuBa/voGvBSOz1ju+iz3d7F9R03xZBeM
LEb7PIl8zQQFT45q1x0hosWtqmeEzLuQ8BJw8KQ5BcE1oQUmCARG0T2dArHsFv6N8+2gLZklKshq
y2dHrpE9qOjsk1SCV8PCu8Ob3WSWYJvoQZNNN08xdudphpRTA5SMp9iR3gbqWwI1suhznA9IiESg
YCYeQFIMMWd0lc+uikQF7gxuSGPtv+3ecEx6D6l0nOTTApgjNB9x67d7wrqrZdDi8vPFMXzfzFh2
8tjOxztnCQfYHA12iOVsaK5v0E7CEIpvY82C3rluKK1AcA1iQXmrEoS8trApgzow2VDv/wsPO66p
4/1fr+M0RBaWdI4KXE/O36WOXiSB2RUUNsFiIy3n1SIBn4MWuC8/qR4+/ugXDsvgQBZArfzrxqp1
0mxV787Qo7R3ITzK0dZ++YdlermYQQUWN30wnpRCgHtZFVaG3gr3V/AfJw0GhdlBsqwTDebW53up
CI5PY7dSV2ca4uumq+KNHuAc0FW1LiAO7KRsxDrzFgGjWISj9jY7uk11PjEwlMf+EkoMjbQJgr/j
grzcJdj1AAET0J9K1xF7U5q8CKW1f1q6ZwjHCOPA3sUvWfyA9gIZKbcUTWzLHq83+WZ/rEvTCs4R
ODvxqY3sSIfYhK7Ly6K4E7WkI3VZNtgvmVJRlTdCE/uryXhlNmju52WjykDZj4xLmn0n3VxF/3UO
u+7W/7WU/eZGhkF/oIg+P2UdM1IyjLvH2rAQCRpFrqYexd2HikIHxddJ9X/K1M60JDeBcknmAfFu
oTbjWt6frR678duyRp3GmdN84+RJ/AbAsKqUA9pQVqGQjWd53szG0IZlG3BmL0+eCvki7DARgP2E
kGqTrhJNfszgr+NqXXy8f5zMuPwgzWczo76YpzCf1cE705a1E+2/v718GeFd51jGNS5wiVvu4GP0
trKPFj0ctB78jPAOPdsCmV0NfZkL/4Fxgx6qZWvBu5fmx3NFNo3ZnfdC6OZSku+lUafshYkfMvVv
1jYP0GD8twIM99v7YCZY0ltOQ12+Z8RcBpkz+nc+2pEj6bDTmGP4aDBEpfF7R0agIEW5aOEQteka
FiehsBiOS2SbVubuDIYiaH+0xdWM3BgiVKfzn/iX3bjzTRkp99JMnbUfNwzzYNtnsuyISbLVMI3Z
jKc1MiM8fzJeegxpYSCloRnxAeQF8czhbkHtRhm/LMyL91yumbpwcEEVChP4EjuHDsrdhgAB7X6r
eZHoCavfg9nRMsf5pTEcicCrTapPBHx+MJC3gckl3ptaYIG21LOYIMIBNxw6M3WxshyvAmftnjdO
WDQ4Wj3UKU3X7C9cOfd4oeBN03mIqS3McupTiJhw/I8DwLgVmMdTzwunQzPRo+S7XvwX4uUjSp1n
l7jgGBym4qFo9gWd2k+Zb8ZMF4OjgNKu1EUjK2gOxU4Gw/t+Ox4FAkjgJQMsPqh1qWK5a8Iy9hz/
By9HTrS0uwGlxnng+OQlgLP6E64ScbphYU+4WRWLaUZgT8GcIbCx1l0tT23a/37kIYdV+vETxGay
RA5RtpiC8aMlE2mEk3xyatQEDclZirTaXzqatMUHQ2pViHusPTQ07DBOl29Fw44quZeM3IVHvUQ8
E+mDOPS11K+INHpGqkOyMyfpHZCl/0g/sv9BfsJYhPIgiSXZ6ETKNsm56XHvKQ2H3NktkHjQpGmH
7U4namfvd+KHs9IAtlqxx4EWQRfCPSZCgZ8vMWRe83RGwVH5NNQTKcOeu9m/kar0JgakMi3chhq+
Z7nEdj/AWixh7/UWC+cJzXFUNWhZDlEexkI/JSg8cIiU6yxLgqTtSANVhLZSFeo5ujTRwWtnE4yu
KZUZuZoripUeWngOAfEO7W+3ZMNQ1tyX3MMhFocCYyPuva3c/5TLDD5nk+JgFIK/amM2qTQUb5S7
zFZnZdWsfX23nO6KC6B7tOAZ8MOSpVOeoHx2eWQAyZ0evR+lcPiBTylAyeWGJ7pQjdxSZf3MKuJy
rDRgwOo5RHLq1NQ5a7NvE+xlCWlg/ZBr+H2i997zbwLvISlsHVNQ2TKHrYM4MjJ9q/+aIimVuaD1
+ysisCRmRdbiyUN2Sf9xYXruxU4VtOYlvY1l5YAL4J2iBaIfGbftzuUsA7QKG4bd6Zp6YH3GHGUe
6YodDJdTtha+nZ+kNQzshkWQtt6AipY5+RLH1gg38oXEyjTn9KTW/AWWdDJx9uEZ2fpY7oMOzGSX
JrwEoYKwihP85ocMKAIiN1sL8MFKjLIivZxDkvZ5qIg9A8tvO2Dc85xqZu4iJwejys7ctSvNPNCq
JyHcdSPrMk7n1pQ5EMDfPyiUXmLPqiY2XAyvgyk7j7k6meqm45/UGjpoYPDrznTlekvCmTzBY/DI
Ub4hbShifU+wkHpY/FrSB7eDHga9r8rSKvuAQ+c7CiVOiURmb78P2GtEz/4fWwy/g6RLBcMcubjs
fk9LUXk2UEpwgUFwrKOaaEReFPHicBMW+2ZakdGCWKVWsVuR/fWGklfhEEjfmLTwjlZhdsbHHAcE
sJwzfI9Yg4CFVersVL2ieaT9+Xv2fcWoveHX5y9YbFRYZYMJsYAPwzcx4JMaPOG2SNLKCbSLQHj2
OVHiBXB0yqPNbZpfbyOX3Ht5F9Qoq+r1zh6zB50YMA2elXPkdhEoJ+xTmB1QONADgbROHV4j81sf
XKlNwCthyoy7vulAHBo6m9ketTUyuoYqG5Z06LaQdysB6u/Vho2uCC/7+ix5S0QP9gjDZx88oK0F
YGuyalL2xRym0anEQlGDDiGbl6LXHUNx7CUTMmbDgFWi93fb3WaoZ5LoKUIeeEvkcMW9HTCyzOcQ
SN8hyLyvM5sHu+2c1rfCkzkTJxbIROKwxu6Pk6AIanXuyTOx0isV0KFWxtFLUKVYpy+CWmD6Viie
fbrr0RmFfVwD4TPHrQExMqWnadcoELNdTCQwB3+6tdQVA8jwHC3ChnmEV9TWMk5DSZ0YqC8MLFIo
S3tvnLwYzL7EkcOQlLez83WD1X7P3Ryybqza7E5KShna23B0aocm0EIdidcK9fEoSsDl5H9iPUYh
/Vf0MFt1wcHTHvGQblDml+fckB8mJKkxlMqoDL5hiXY3mgJJ2c6nt/+D0XA4E3ZCGJoy55zrV6O5
sbPV1w2iZwZAZeGd5bPPSoRcdxhCicl1GT9y5AKMiAzSf2fn/PEOBgS1Vafs7zQT/QGcoWiTLxMb
97yWRGR1eFqLNIVfcaV7a6C8ZeoD8Gn3EvAjkZVHbinbSa/H6GgZGOYIFkFOhV5ef1jvTsuhmQT4
nyillzRaKEjm6k/lRksfn0Cehp3oGZ6s+suvJgy8etk2Lf+9ytQdohofnB8j3xrapQsXWhplYILk
yJuUIgwPPAykWKNM9R+mlzqYxvp8vEdGTo3/d+UoBq2fKl38MeeueI3ffRlyt0UpU95cuD9dy6pu
AZnc68lxQMVWlMG3c1WdtyYN9K9IL4EWvGklvNgatbuSXhvBXMG7NpUd6MNNDCx1UGd8wg//wQPm
fepRv4WnL4CqyOt3/LsFzYIQ9BkyXW9G0/wJ9i7CQA1Lx46uNSDKwivdKixR+aj9eYZEzIOt4DjY
TpPa0qRLh/BfvSjP/GIxy6NWgb4gd9kW48bGkJZhyqcGjwRbPMw3mfIl/rX5n9gAZyVRJTXgOuQo
bWiJWVuxHj3PEJlJkcHXM/2zKbMPFm4c3LuI3iwhziatWUatIilKXbhEj5bVTlHLEs1ossjHPGN4
et5zqq/Qdv93Xr5K1x9zyn2mHYO9rG+CClQxk5UxpOuMjdFR8OCX1qg0vDRyJuRHCd0S+Q7EGeAN
tIMwKysGb58VVsrjl3zZ3dOnaQkUZZaazpB6p2viiqtQsFXEmm0e7uaxeg12rGeHjfnQJlzF9hGo
sfNhxpZRYdv28aUZ0IWnWYmTvqRfxgjO1ZT6D9ehljrw+JesR69bCECtWr1RZz5zYcIuFL2hezgV
EFHYvN/ZTdozAe78UY85NT/VaI05aG3Uf9UCvkxsNxQsIMjlvaZwozLIXULiH1BMzvrILKBTNHYQ
JhiGUZJJ61Q7/9Jt70lFCKxAMyxiHNW3JZXGfXLleHw0Y6DOucB7+L7oqNWi7kHyvuGDHqbN7lew
DNCfiJF55tgcstCVnk/q/4H5s8oBeKGTq5Cae6MsVDB8Hz8AIMBnf0YDq3dR39roYBX6ueVdd8K4
zr9C+d/cdJgcGle/M46ZDuuuOWP1oAA8QyGkL8aaP4KW/cNP4voxxG0nObgzmd1TMAtV/i8Xus0+
G1MJyrlpmnWBHFA5E8oJuIDkNAioAenCvLeTwv9B8F5io30XRPTATt2Uakn+uBvvOnoOL0PY2v5b
9FNbzJoQpXMW9Uf2DyMi+2lJxd7fI3tRIkb+ndXcqsGi9IslisbFjG512aG3h3fYrHKmQDt1fhY9
apkxAX5Y/k/a9kmojL1JLeTHOWhOBe6kQa1pcaQQi3mNadGfVxZou1pBFraEgyn2eTR39X7PQ2Lb
QYi/IZulx70wvGzh0WItVgDX1HYdel6uE0z8MInL6NasUy1fI7qZb/qAy/36EftczK7hccEZC3mq
cxLhV3coLTe9k9sGsYXAS48E6OZK/kro0Ju9M7twi1KFa4XpQY+0f3Ogcfgjb94jkqdPMi+7nB47
ykCkfq/7GI0HCDZClArMvICQ6nWnOo1S2JQFtpehoe+8T3wziHxveWGrTsRwkgL2DuqKn1NQKT/7
zXz8nMrrWbkLmvXLyUy+iwkWPOvn2GcBhH6TACH5eJJIXffFJwn2Jx5j69Wrs7Wc7jcwrcbILT7H
m65efgmGlqyHMeMqEx9ffBFYyv/FSZYRqMhJ9rJ8OpDy2bB79Ey9M8JZA3eRqsvOamON7ffJapns
joNrGksyIeBVZOBU8R+KYn+qACgzy5cl6MI4mIdT8EZXPzIyxbdGez0BZzJzASKHEitu7CqX+OZ9
Df7HLo2O/dxDBQCBNLmpHiZ6McanJBRI8VFy69Rf4wA/cgLPH2A92fgfUCXpcBwMm5C7Bn1MHvRZ
q7o284V13JRMINk+BjlYgsy7W0Srixqslw7cEBBGLfZBykZFx+EhjcA5XRgf0lCBPP+cES7FOlsD
1YiffcKs94iolf96a6gnh72lza/t44jc+r1eSXKq34gTE/takWSn4aoll1pEoSq7GndzLzy2K6cP
0MbTgG3e47jWAU7W30s0dZUYf1QhFiOSdu1GKyx6vxMnn1xVUzoB3R9JNQy8cqbwTD/h3yLh79Aw
qscmfEO3+abmKIF2kjl5C6Tz0R8e/1acYrhNTpuDHeZFpd6vjqtMGd5TweZYeXNYQLqHo39k2kH3
9ccL7drzi0K8OTfDt6pxamchu5vwNMKnwyiakCC4l5kQFAfyRfQVD21ZrSnJBcda730KhLFT7ceU
vTvHv++FgIYVlapIttwqz02BEsksPMcjQrX0jLpHDH5oiF6ImcfQoPi1aEpXXvsXkO8oZ8s/4HGA
wLQJU1JqskPyx1/Buq/I9AipJBk9zNJxgo7+SxfhEiFKtWob2ZyloX9H0eCHx4no68lSkAqmA7kK
sItdeUoLTVt03vbDWZrLDQYn45hpCSCN+XcCGd9uyD5SZ5jZVSf2yQ7LyB4nfFYLquJU1Z0N9u9F
gX/Xj7gekUtn+PfST2u6Sj3kc5t/18mm4dBr9HO6k7dCn8+6+WE6Ae2rjIHXiKS8HThLHnq8Xodl
0M0eUcjlAeP5S/TGluG45obIebneojsL/3QLdyAhbjTP7rj1W66DSBIOwlT9XnTl624zajdtbzrQ
QIW8bbUHrr4758AFplHi9nISHdm8IdSV693sPQ1SLP3kasUd4ybTNONDuf+xBfVv7RgRvN94Fc3H
QwmbykdX8nug1AWkSiFIlWC0aSE03ISHbj06vjOYvCMBJ2Rffq5RxMWBiKF3vidwkhX0pIBeSuLT
w/43TEitI2JcXhMq8OYd65FnBlqQeEdS1rSltf5U3dPnUR0kLRoXkQEna9+rtKfhLfg9tPoxl382
r7mMOE6q+CIBWD06a733Wu7tYsgwXzWqDcnwR1Fxn6cvRlFULtrLPdnFAf0B0vWAQIj+iZLHzE8U
xyQtrSs9eH9/HX1el7l0pH5ds85vxvrrNFhgpQi33D9o4fTo1WgxtLl+w5E9fi7eEjAgz4Y5WvDh
Cxx2j20KQvpSsvt5phbCELUXW1sXlu/f1glQHDbGRdgR6i4weHaa8jazb74mDEBe45wyS0z0cnmP
js+bOQMJA51GDdUwW8i78prbht+B4jcRfYWVExRjtpiaVqpYF9zTUkL6yJfowreg4H7pLGB4eHPE
ElRvOFgHDLT10wcvcQkP5WD+VU7nNf5ZL97vzm1GwuDIHk1kHXsy93SFsS4N6VkTOTNL/qSP3v3C
OHd1L3GV/KJdPxPHu1/VeVt6S8rVOaCCqZ9Y64GclcDte3g2ArU93Fj2nPJw8D4RsxDl369Yqo0r
N++WmWIhNVYoYYXkINdTcJOzoGJI8C/kH+REc2XoErT+idNfmbhJ7Za34MKpN5Vpu+yqkKcNqkAk
ZcUlGxSEmWejcvlZeV8AEc+8+XJdX29Kkrf8krh2sOFdWJgl6kP1WkJZAvNCU3MtMbB5WWLlOiAL
/pQgGiRvGrEQZI+Hj/IYZVW02qjhqu2+7f0S+Bl0z16ouXizwQ4XMAunRUQKgEZSm+g306RAnrrN
l10WlTxZUIi9pILTiGlfoL5ncsMNN6k+cF/NmjK8zEMjCGVXmMiAJ3/hJAbwFyWzQo5kkKh08cRr
W/VlCRY6vYd5ikpo6wbsQtAt3/2BRtZQDMlwPtudMOsHR/3k4eB+hAiOB8gu+8Ic4Sfte/TuIr+I
evPgNSog5lP0ZFNlgxP+j9PwhaUuvQ9Lik8U5brzIm1InjW/1UGPh3TJy9VXobFzOTqqnfBelFta
gX2oOyQwuPjjlLhaoTZQPKeGALbodBeROp/5q89a80lN3YXgFjJWFoluvJKVbh76gGWkSq8Sx6G+
q83fHIeTKXiVQM7/F7oNlm3fee3Xfau6Llvc6gg+5jR8TCSL8Ll8NH4IGw3jM4zHxm8SLS2oiaz8
ERMhYetiz9n68embxmDOnhH4jAI1+ALqqa4v3rKD8CjVVpsS7qkhHG3qh+NnWlosZlUuELCcoz+8
1Zpol4a4IuDk8djyq50ZvM91OoyBY/m+wEsM6Rk3XB+tbRT21Z3U5CPo1kmt8JbS26wQA7U+CYv9
YN4gxyi5wV5MsEAaDiDlRcfCWh0esBkerUtFaU0rg0SiFeLdvyO84Hn4HQQV/n0Z4KroJcoB5c61
sbm5YVA5vVUHPRRSTRYr6zbn9aJZS/K+Nh8RLGQaZuN2rmSQUH6G48nGcVlotrwAmxe6+8KfXUX/
leBU5iVaa64LNqqa0hgE92oKP+4/BHumo1Fh9mL2eHbWK9H8oGj1O3kXNeu22SaLzJ9Pohxn0wAL
82/d08uR9hrtMRpBJppXc6uHd8tSshATbG2d6I3IyfWqFf/FtShRFYGzdGhVys5/nx0GnIi8DV39
fYtLfD7pfy9HkaGCjNHgZAUB0+mXVUQsKgvmYVitw8/F/+Yn8nL6lWYiXd1IiNEHxNxhY8mYrn93
CH4rw14g2fbXvqynQM1VOVH0cZFM3C78fBeNPqjDSFbWO1nq8gLP/iQpbBJypAlnPsNKuaNH28uo
qRoHNcpNcJsGTeXfyPaT9jV6OGfoXC1Q2dL6zvD4jUc+/ULY/RZ0sD6tLP0e0WnVSlcZTo2noUWl
JyJfh3Tt8mFOahzzQMhxYXQhGgaF4BAkppashsvehSJO5eRu7sla7F3ji9Tad6a+L7LvcBplcYgY
LHHaLCqbnBFzPOvgiz3t722wd3IRYC8AvFw+7JgS6r30KgMD5ipNo1DmZPT5JPjF/cEQMUahQFxP
Fg88FqUUCr+bnK4RzcUjkk/ojiWagPvp0ZIwHKxMV6V572im/b03znYtq2rgdAdKbCSBPL77MZan
hCB3SIKJL9cILfgoeGttW56cRnWillu9bIOk0jEOs8u5mwZP0eRZnJW46WjS+mmqb8HM+1x25ZhE
fvv0ROih1U4dIMLto+2AK0XvjByJE3GMHCWgT7SKfVyQqDN1kPuDau3qsiDMGjFwvFuvl8yyByMq
3AFvm/l+M15CPUiwm7E6d0QMUH6QWOWMhsUo0sZu+5cCehsF2+K9W9LKOc0hzqMV/J8bx59VlJWF
h1awAuUVsag6YUfygmUVNC1KsVOs20gvdY8r+g8c8xJOK/JS3t6mCNmIRsocYMDeyi+S9h5Bp1bu
/m8rHIzCTfO5Z4/F/YuvbkkyYGaFuxFvvBSB48a5HU4S0O0CVktQOQb7y016Os8fFGSpmt+siQ07
yFw4iPMX35Qqwd8otcgCaq4EPVZckKmaHfQOpzphDTWHO1kbPFzqle6FujJCYJpFr0tbdEQKtHfx
vhsC8CONj1VEnq4gPV0Hre7pXImH4rckbGn9lXD1sVY/vy9F1H06mB4B88kCD1yCbgIMQ3vTSZsL
rQ4m7h27gn1eIS1FxJwqs0Ff9gt9uCVC9RM8cjbkIPs3j1v0toz3r9dpImjYGekFq7wm038aOmjj
yBStiYmPITXpTQ8Y5TTC1k66Khc2YnFFQG+RXU3hoWv/OETCBm/kMSeOndt5yuexnQkAgGGjxA9Y
Lk+ug8NqxTDlBfTfbZSwP1E0SymPHi0vOOEuU/mGC8OkHU6097TM53cbjsjdaRjuMQ21nXShC+mx
52++c/CM2Ad/EGOokYTB496l4Z0iLwBeObVs1jK2ZWax1q5mj9w60bv/l1bHw+DUZu0M+VdWJ69c
Fz55X6bFj1prCPkKZ/EQWVKggsIWYaHvkq8d7VDGWL7Ei/J06U/A7ewbuG6y+R308Y5Y3bdiHU//
QS2RXn95nkXoYfnOu8ZNn1PCvaGd2tUVkHbEAqYBXapCeQ0OJpTsCZ7dh36eHjOngrKu+YVEPYDd
kAtsFIEjK/7pJtbt4AOu0bTtsLtJLgekYilbI8nNk7YUVoGBVhJV5A1F0OwWPQ+xP6nTU3KU3AGX
+1mmSWBald5rOHKbBzTnQQ4SNHVFaNVo7O2BtTJBczLmJkpNtVbm1/iQ7FwRfG7p59ep59NTQJSU
MqzpqFjEpLVpDX1O4LOSRQyMfBJKIX62vgMBq7Q1feohjABnHtp1o24FNeKMfjjkWsBW167Ehy9i
HoBsYnVtpunMZC2WOp2jvxgxRusFTtMTcHV7eh5OBHOckZrJY0hnRP/+J+zl2psZroym1g3LnYzY
VkTs4+/WM0mYS4sRIPYZuOZajw4Oa4z8+OUQzbG9OIfLf0+ANBSdS8wFVHeRn1v7zrgMJd1nLIq9
jlVR2aDDjO+jmVa2eL8g9nboVMGp83X18cBioU4xyWZdJebyKrNvWdhnGQhKQW2pBu590TA7ig1S
RedbsCgeg/EIykI8x9RhI5ROiN0QdXs1Na7yk/jpC51iEPv724ih3G9O3UsVOn1REdDTA81dQMnq
DD3dDJ6AZNgD9QB7z1KLq1yobVGxmGcVx2rmZoloOqNnhstl2SbiQKSkHvVQT0HTbI679JU3C0M8
BFrz2PZdNVjkOBi36QMKWSFNPNYNHjwQbEkNExRloxndFE7WeAa/85DGa15cYfy/aZW6EGKYSEdA
p3OFAoCuDuVWvwD5fjCmJ9whJi4+P4ZbKmVE4MfdOTOecrqdYQXns525xDpSwJfRDfg/Am2lbN7B
ZnpvU1a7WeK5bD+27O9UbEgpLkypBrFijYW2CJ39HXgTQ/9/1LncyHItiT3UCcolAJ1BD6FvTIOC
97mWrqshReLXQJYH1X9mEGjxhesokzsgsgA4JXgcKV8IUEjiWcJZDDPSbkFjPWqbTZgKDEAa/XxU
h4e0iqnpXsENdcJYy5LlNiR3fD9nPFnp+1k1C2KlJhvrHJdl7aVAoU+HzGzAlYwfEIYEBJm2XLnb
iDYtD/IOr2RkW/qNzCNnvIHXcQ5BOjTJ234h1ZjEpsmWAzwwe2B3vErnRk7TV2CwyDYt+NueIUmx
IdiHnm9FMTjyN8TSjO6bVCCFO967x+Kec3uiyoUqw2BQzh49h6ZM8I4gq7l8PuxpyFFcsoeDznjU
3XC6cc+OMSjuSTPAyz9zHM85eWcbXL0gpk+589R3DtXrHMWenr3uuiJ6/R4YkGX+V7VVQ+RG/R9h
W/WVoPkloZiCW/2lsh37axqRM4cwd+1UXFYO3oZyKNRcnWThyTu2W+pymFA5w5hxXl1gJRKGiunJ
SO57MmduoXZ867ZisxJIGLzLQGk1qGmF1n2WQySWJWjDGezO4890RT0qvAndfhk0/VRramBYhaYk
WP6XEQJgK7Hquvjpzz0VrEogc82RXlL8/+cIYAa66G6NA8uTnECRUViNRaPd6ecKtDDaH00LiJSB
tXWcEHYKkJJAeiXwycLPnPRWmHAFuEbbO9IZfPkuBQ00dzh6tZ9R6+Dbm+UIyBXXr4cURURfeyn9
UkxhrziPFKcofCeyNjaDVN+RYKBoovl7g+V4QkmhADxcbp5jA0xEoO9vX0EYaBp0qEKWTeF0WpLH
cVcO4fHH8OtF1fzNZzxzHjUSa12hDZVtHSFjA60OZA0SVQLxwHDQMaaNIC7scf8pRUmJei6jxmUi
Faovt6lG2/rm03FCL9gGSQaE7jWejGlpfPsb1PriQV/kqBP7rWcgh70a4naowqjYFSJ3s5n3sxcA
8AEPvTxFXBKaXYYvWWRJKw0AWtWP+yyp/3IsGBpq+61uD5p0iTxLNP8rlKl45DljEN+cdEgfBJNO
pfus2Km9ykyVmAIggi+HHd/obWFiFhm4OoYXfO3VSMq9x7e70dAuQLn6vAcoQ6/Ydyu51R3apnAJ
pyxqfIlUzA/SmA8CryuVZGEpGI3ZssbnMo64H8vjOvGMw0iWYzNBStl75NOXr5toi9nnBKdiw92o
qMUmzy0kzeK1GXnw3t72SYEmXlWAj6/uc4Npa7DbBfhyY2eVlduKXliq7A5OjW3q7s6tuZYA4ym/
qD3uITZa33LtB0ktQUBM1XmeJu/5e8UTzP63UKguhWJNssxqJhYZai9f5i4YV9OSTKTDE6ZcUdrC
UvbyPxGFMFVxJwXEL6yt0ngjPukRpCAf79ucjeMIiHvPmBNR1Jpdr+7nxMpJGYpqceEhTLMXv1Pq
ItJ8RIVavRI5Ayu83Hdxj3s/m3ZXsPEcv3iQF0csDxaidxxAy4o8kK3C/I/BE7aEqfzCL/nbEYQl
Puo7iUE292W71ydJcPP76ge0X4jr+rEskjyo75pDC/kPA1Tb2bi6YdXZNFQ96e3Lh4Z77FsyIbWj
FR6FnWr2wSJklATiqbwzlWuvcHgn1ZwflkSL4xVT1HovTGTH3dOZthoHHS2CZZ8daOot4Zh/bzoS
Zia+d4KAZx78RIfFnNHps6uo8Mpq1tofxS68w0BeSg00KzCfLPYFilvgaebQ1V8GMWfUCu0EIqls
sEALFi2uDjzV8H3G5ynekxGD/d9t0Wbz1PJd/rN5QaZ6J4QbbFcBftuWjXb+CDr+NWcjrBe2EfYZ
nVf4pCVBPJ17h1HBMFb8K0fvGjKX9fqJm4TmlllI3WiAMbU5wOL9mFGEgBuw9nO7eRuJZBBkdp88
t9cLbIWsgDTcqBI30s5usxjDoAOoaLkW8aVsoz5CxwcZsDFjdzjLiG7ek15QpEyCysSFzpz7VSgF
nQwYGVAB1hXet5ZdrevPutvSxLJA6oVJojhkm1Pj31r/2CwSWAIuAADchWIxtgNf1SLqnke94jtx
IsexyaQBQjg2+gkuZ0bmidZmqJ3GkBPHQPtxfWYXSQzzTeAGMXTL71nPywFZaY2xqVyvPQVBf8ZH
Me2SfZbBkH5FdRHfBlk9Qr/b6JLQ5D+BCE/nMRNBPnAFtDZiLZjxJwunsNAuJQDefkPvh4cGMU2H
U++SM3KQCt2/jKGojVYxZ+TNfvrpFmChPrDYPU72pTHhC8KN+XCfGYRNX2Mr0BceJxBmn3ZurVNr
ALZDkU0BwEVRC//KcPjbATkn8wGjLTqgBHMPA/hg9T/7mhTWbnI7kTjbzXfaNu6wko+Kmr3A6gSG
91dg0TyWcDVVVn4pmX8o0fBJ51OnYyCFMZzc84t3ZNmYcY2TUxit5V+eVEr/Rs2edCxS1k/q6O5n
WS8ayVnl7cW6K+EFEzCcezrestpYzTgoJYF/FcHzkQTBE6mZTsqgsKntys1BB2Dv3fld23SGeUm5
OkycYi16En1TMWJ1ujlOsnOdldX2LpdYc01vdgzrNtbyAwy8dwCs0h1qHYPsoqsGkcHLs496CuKp
axkIVgqRQOzpv1hWSlLHJiB1EOTY95RZJasdsXxHxQleVqMyiikfpHcZqyvsisSlQ454uenr5zHl
0WRg6cJKJuww3Nwsz+qK9u/EKZpoOgveOPinYJsFy+0qas3NHkSFJ+o1cEtszSt7n2vqWehRFgdp
qH+/gsTxQXLE0hDCh8Bb9WI/YDLLGHywUINhe6Va5s+8oUgnj9TkHvwuAqBxk94REaR84MbxDUDe
3m1bIzbpV6DvESI7zHRrH7u4rjKlRVb1oIawEUYvMnJSIlWjA+JFjijIu51VO4+levaXO6OK3yzJ
uBncKFVjXGUECy91hCk+dEvf32utEZPfRmxVKD8nneDmY6JvlmsWxd+VcMfByfWaj0AgUveq5IIS
OgXKAabrJWk8YfoyElUG83QVTXHWRspzDto1YA2P1MU1iPJFPZdWMCjEtckDq8ScfCpMsaqB4J3K
U8ado33TqIikIZf4RQZ6EhffIjkqdvqGZFHnaPX6Wq4oab3FOF2Pw0xkzjl/F2trMfpBR8RzYipa
DMGfFFoD8zj3QodQWA0nC2y14239xiLL0wd1ThPGpY7BiKeCyD52Ow5fKXpaZKOTbJRZIb1gjci9
/QEv0AhL68DA5oDf/t3yOQQvLQ8OphoAWtig45COYtiCn3i/XbGUtxBpf6G2dtqTDWsJS69Gc0Wk
zl9pY+b70/dOeyFgaQanjh19JiXxsZ5/yhZV9rv6sdVtlO8m67jxGXan59x/+1yySDYWC3LvT1NV
jiZ1T2lRRSQ9+epj/kBeA3VPisfwlT1WY0+/nEbfFKXu+7oQoFO6D/TcPI9lp6I6o2JsaegHafj0
8L9aEOShC32kCZqzKyZw4L3G1C9ddT8sJFYMi+rwlNbVQOSs2G1GiM4HIISsV/LShiHqlBywTe+Q
G3yTjzq9x8vG3jw+MeccIckLJOTtbnrT9MgHb0qtdwF3hKv9DbilEtK7sFUM5coHA9E9IyJAeJxO
FfKMJvAkKWJEQiiD74B2rl4CercuVDTXLWyAj4negne5JKyOXFWxbC6SXQiKstXR21esFDEuOagD
FIw/ghwLAfiATs5mG6GP5M42H/SfQUE4XYM3PyUuHYNFgWmIWt+VzJoX5EgaPTLHhmqgTsGtx8MF
xzcyEBtgJ8ygLeGCeRYPl4IXTHUmbjQoevUUPZtGlymaOjKguEz4FtaezpwGRWeWlo5xIFJ24PSM
EWI/RUfG7xKgjfRbGbApZuDb6ond85xgIyCvbtgFDjXq5hz49HSvyG3LoCXtfb7LMGoSPNUQnD94
qDDAr/b+WxQXWqXi+2ybfvWFutr5u5pte9QiD2k8cBMx9W6/fsChdVEkznpwG0ONdnJRxMPYf909
A+7E7OPZ2F0r6hbzBblH40Wet9mRIchky1gXHaGHzOUXH/zgb6UrLxOQwOOJ+bg94necetHDx8gj
37Gx81ngClWBsbfiQgOzmESN+TZbPCoqR+/o/lnh5h3jia0xh8ZFLIdNfPc9ADVj7qt9m+vAHQtH
psw/VWkBRnZlxyKf1DrWasCFcBKNwSQlxT/Lv6QO68cRHyd1u/+/CWPKCMhz9urdbl9FtMGjjyCL
HBS936i8KkW1TkgmxmdC7fbRrfIGem3l3HPk3/sLLcN8279+VJKPwB8xi2Cumyu3nMHM4s7q4vvt
0rgDrDv6ZyPtwXFdBvsxDoirGpBoiCNN+1YSH8iCgNItwlGxC8w9kLezFRRFaM3vsdqHRygi1cNr
vrF/RIQrlvOUOOXvbNubSGrQZx9bUfNO74iByMooJvsU6EefumVkVYUhNMwgYmWln2F0uHPCJ3Mo
iYoqqHtfXwoGJsj/lKvUbAY2QKpraZzORuF3PyUVD7D5MfvHSOwS7vIWnFjnrGpIG0BERIa0B1u3
V0VNYiiGrVyaJKilXPvHx9DC54WO0hQ5UEJwnrW+MaSwCZniswJyLd2Xzn2aEXUaky+hveEIXvuR
LL0pxM5pLxJCcalKh0TmyzSbei9FX/So+MjfbrVrOPsh/HRL6AXtx0i17M6stBsBbQQSZAqPgI6S
qtYlH4LoTAp/v9pDkEV/WUjiiE0QJFd/IZZLd6YCWHStqSqjbbgbucLmIe1BMbL2lFfyR7OODsvF
RLfP0tVVF4a1KXVZUI7lNeMHLsg6xVXAbSySyCi5KPEue79GHf7COYbavB5RAocjFrKe+gw4m2mF
EMpiqz4+8m7DqZlC21PN73GDj2+qYxggqiDrJLFPdXDX+IcpTP9odUWysvtO8EvhQB8hKqriODCU
0Ctkc6r/FZDDqavLdl3YnlRPEhEV6PF8JhJE/cwAPC5fJ6ae9SpVfYutWcCYg/yXLQf0tNJwN4aC
sTu1a4MXVdkTyg0FUWxwljO1mTd0NwErPyqvvA5a+S7sDMC6UrwCtxMl7q7bYzqNXUiEcPbmKJM6
vnG/5DUgdaEqNnylBFi8G36XEQilpmx+Tmyxe65NlsstNKSmr5aNJGepY8WIWEwDGBF9jefYk5S/
FIx68y1EJg4xiAvtV7F2KarQ3ZIx/RapynoTAmTsXFFWxcWFLlLpbcMJRkVlHXR7P6IohNadESVn
iCUJmOwGTuW3Dx9S1A3da5XQ+fUUpFOjSyXIgB1yziG/BE3SeV5s7XnEWRB/skGvTPhWNE3NRLAH
Gn4wcwxMStR27Srg0/bOMWXWA4gocKcJ5mBe65hZXEzh0sZz/0AnhCMvPNLkVYNTDeRFeKq6muRi
Nyy0UMQ8X2vEEasgJaqikTAkukYWI09TCjGGLCjw39tvKLjHwcGXDQi1mKI1Bi2KqcsA6XmgR+uK
a1Rrgkb6CltclxjGc+K0LVVyLzlX20A5k7omX69xOT9huBg9dEiPHyTB/2LNc+WdfkN8VC4SdrhG
7D9yC/ATMwZHbY6b02Hw0xUZ9PcCQbjk3aGTahm9N8tdE65NcuRtCkRLPSnzYcc4vBAffesohvP1
SRoiUK8Q6x4E9MuH5q4rpO4CgmAScyZRMQJ8TbukUnovW1IE4lYomEzD/LoE+2LFK5A0SEFGPibL
A4g+y5TCIHD9HnPTP0vMHSV4owQrEf559S6PDOO6fvEuEFQryVnF4wWx/Pbms1ZNoRCM86094g+f
l05Pku/ULA5O5W+XLUan0b3Qp1WUggFTuJT+P678vQcKmpzkJEt0JHWy5MbpCeOrzWKrWV23GRCt
Tb+Eh5NSVmmmlUl2DGgmSiS2iVGoPSn4XH8RECg+CQ4lKz+6BGvJRTxcnmBIgQSkxp7uz0xOOhVM
qY+VQwXLsB+7GP+c0I2cRJelSxdktmrkXk0Xd9WPbbhMe8FW8jnM0kVzyOImX6y/sztWsrJmeFZh
AQuz/fCBSMmXM3RTh5q0zTJy/mmwCLKn0Bxshi7iQxoh8oeE/uC5MCCrE6BnaVPa+XbYOjSu6ubz
vZWJBvbwMRK+f2/d6wbnX9LxywFSUEYbJqMKQNIezeHR62nG3jkss0l7K+V+3i7jcKsibQGanycS
nIw6mVTdc8jLCBYEpIX0dZQP55yFbfSHj7Y3gPipCTUmIPiKmFAp4XRW8718iqjo5PyWi6uwBYVw
MFwc2s51hKVsLDPn8T0EEXpwQw0Fv7m4gJorCGAw+z63HanHR/UTrhHxBgMw89UyFuW5KS1gR31Y
l9R03r3Paqx53gB1P8fnWoj63Jxbv+bLb3qIodb8qZK+tqkvjDpJy8wQxbiSp+Y+WS8D0wTForrf
LJSVYrJwhP7nNPLVPMrMiJSKvUss9LKVMwgbBZ7LjYofoocwcoGAxu9LFfYAsnw0uXEALgzIiA0w
a7SzZvng+P6KwAhJKvIkXoMlNDCtzH+PA1bhMyZwERc2kIxNDgJuVudgyyZfaevZMMd91mz2UIlq
Bkg+lxmRPjRKFhYjG5Ee7naxBGUPlUSOUm2+AAOmMQMHRkHry7W4DKuHGviZB+a4QpuIv4+F3WAC
kWn0ZrDBHuxUf+unxro3EsMxu9mZNdCz9/wh7TNFeLi+1f9KRkDoRTE2ERhOmNlz1/QDlUCnXAtG
o4I5kIVLM/Z/IKUtQcBs5Sk1YR2yz8SkP/fO7EEvlJfTbqgDNORUUzQS2Ct/Sx+MmqXSTtbQUkxg
HaTShYDbKk9OMWcmcG0ZaNPgJu5nI7qP0H/6I9Z58vNjnJXnkdxW6sNqm08mnZQGddvkjuWlN2J0
nmy62iDH/X+93lXkeK+1OXYcksctoLT2L20WRq5dPrDUp/UxBv1yF4F4NEzs/n022fb4eXHMAgq+
eZUJhz9zjpi28vSgnWBX6van3qaWr9tkboXcLkEUP6XVsBGzFy4lRyj5d14vrSMf4TFejiu6aakS
Zyj45zRzWWzdNlS6q6tvCOGQRDejj8UbIDbn04FSwcNNgzr8Eiw4CUEOPTk/GxYZzDNVpF44J0Oj
6rb0JVCEUoSkBQPOK10Xz7sF2p17vKFyj9bVGe0metzMxGAHj1o99JoonKOYMGmR3B5Qg1+FkygA
BJemCnnaL7czVeIrUIzbO2yw4OWiBebpafblu/syJiMBspVcPSRifxukKSFvb55RVpMrXfZkXkON
OIoLv3tNWF4VQ0OmUDlWkOJNiJLjXXRVMgV9mueGKuJX6vx3DHg50PSRHshll5PsVlf2y+gr5YQH
FNrfQ8lsX2ve5+LbI7JJv0tdEQV5tgZUuQZ/uq/OVVK+rzsga64g4ElIPRI/NsKOyqVHPlo8cwri
gFxG4aqf7ZqS1/8DPuuTYF4VeFDz8cBZlVFckyqTDeONMydMJD7QPqELL2mWJa4xjFe/YAyGBtBv
uPr64Je//mt2ucdB2DDGhidZ4W7hSSY5JKaL0Fv+EJZh8mku6hYoJOz3MSW8bBeGJ+tzhyg/1ITF
u9CePk9BwqiQ+qgDnWXXai+8pEC/sXrO7d6hwbLamb59Z152NRWuHxKys0o+4TkQwcTjypBnkB+m
sKYuieBckYl2ioJOR6g3ThwviZpT8uVduMr6igefNCkNlMRiILGWiL5HukwLSAp8DCH8ouWARNa0
oRj/bHtuEzveKG1jwQSYd0rEg8NBCLvIXgHC+sfU/Mf/vJR5lCVPYslR11WzaQnQ9h+FmnkxQlsR
grIKP1lkRC8Kv6XrDESbRBcx5zSxHtGw5hmK2oKdcpdiHo+/w6A9b9YL3umqhOQ6xXCMIVehQFxd
ijq8rNiNF7c26ZkNU2nSyqs0HHBNbzRLastcCrtfKlbIzoNzVq064Pd/R8xUSchAixJOCn30/G3R
9YTmagWA0QhTww3t6+KkAShJXjx5EsNpfq654EEYseHGDGqn3ImjCLL1wosB/6ksjjdafXsv5t8v
+2TOVwQ4TJpYGp9fwA/RgmqG9SBiQuECutfXb0mYnuQqYt1Ro46A2V5mWlH7qJG3ywIDtGKeY2Hx
DRetV7X1t9zDwXTZQmIBuTDiCHd8npnrpiyVcRZnv5q/QIqilC1QDJ3GLEtdwsx6Pd45MJatCd9r
UKlJTnIJjRkRaExueldFEaD2vMj/Vx1wObC8K3FKGB8S0U9sT/8p8IT/jlFa6Z8bKEb+PQdIZQL9
nXvvRha/2Nv9QDV11rqPful39n2AEoRyf7Bn1ykmTGIRIfzwkZ9tyzfKPt7LfFXCpoBdw0KM1uqv
hldgadCm83KFVhrx4tFW7DyeMa13Wus8J6X2gzWCkYr1TswnK6ArKoOj9sXrBwu6V769wACzucNK
6Dvks9uEN/WBObdXRB0T/XnvQkBddukwV7LFRKmjWkgl6NM+Yp12Q1wi0t5uc1ORDCmbPMa3ySWY
pVfykcgwyQD9OQDDPxiH0O1qpT9tf0j2VwikAbfrCdDsN52hNhR47aWALkoT6Dwf6odIr48xqX4h
yz0QdaPVhGH+AHGwtvgRxIMK+5vj1/zZHFs6qeS3Ziu506lZQETbE+4I1bTdubV3UWfLJERglDdi
p249IRdISoWyfnkysfwDUY7xsL/BYTxaHR62sx1Ho/ER8fGbKvVGtsU8ob8kvUJvrpXq1VkT2WPC
IbgqHgiZwY3gmz1cZOQWxNnTQc3ogKk9y+S5kWAhxWTx10gTLCxAnwWa1tbPWuZjLqJkwadtg+J8
H6FJaJzDPPG0aJxHHxDp6a1gYqNGEhVuCm18RiDLx1P2DhzPGATu6VKtmcMrNExqEUa/A8RwqMjc
R21yajqMkp7IOAIXea5UeAQJ8Yrth5g/L8byEoDDMiwjNngO9yx+3JuGgc1rhTXa4Xp8YDHyi8D1
fBqxtgNv/jcee3PbtycxtgOyVdfMrBQ7O/jc1kTcxtBiwDsHTnY3MXGvkENgUZI7ADLpo6hXdL2o
EDf8kAmw9mpxoXGkurHBDih1YfLVC3oFTk5KzHeHztaCJ6Zoy2SjF74IUmtxV1nzVfKZkcrnkXqo
WD2nAjS5HcqGlOpL//k55p0t+vwSsvrhh67KQHKgYVjq0s/4zrkJkzhVNPl3ynVjzBlAujAqYy0h
O+21R59J5e691xHLy1C8n48Q7awWBWYzTt+6JiaqhuDcd+JeTrOmFstrE5eUtCS2qTC78bZG0Lv6
aEHgUL0xLlbC9bNBXGI07Idx8gJywfk6/Cyv3lybXTqtTTK+bfcncVSvbfnCBrP32XfvJWfJetn2
mjZx7bZl7XaWDemnI4UDDfBvRCu11oxiMQ/mc7ZRCxGwVFnA+w/JKgO/Mz5GnI1FIc19vSZaPYGV
0yzSM78nG3vVlZG1tNeO3cFkXgl/VEZ/KahhRPTddsi85updAJel96skXpCxY2is8tz+1R0Bdw3l
WOOCmoAkDQaXhBEkd3gRhiqQusC4eZ2EBex6wsT0xMNLnBRi+iGQOPh1qOs9psVx3UxQ7rM8PKXy
JIzzal4wgm6yx4MiyQYujF3G1QwOPPjFLOQx2IF5foLRfPAhljjSWoafFz6Db/o8krYnVmbTza2K
wfl99vzc0gVZc1FlOs+lzQkffrJMgYVBdYQ2Y3NKqjLXwOq8duTnjMWujsKtf43HAV6N8OST3a5U
psaBSunAL78t2nvJ0zR9ibUqmFUX+vPAQ+oZxulqNYK3PvVA9e4sKB30dAyM/Ik4Bm1WuNScHNRZ
JeiceGtKJgjCH+ooPjyULVdeqrKqXnk305dQE9fv5TtAXdBxI5LCaIevt4Q72ScrmrbAJOhX1/ly
Cc4PSOuLENia4E5CBuDPn8w28rZ+ffs9a0B2p4wUtIw5YmQ1sMmCNUcHKrNbpeJkOP+6EZ1qMvn/
gGQ3/O0xEIYBwjfvuj1vtr3UTTdEqWLol63TPzsxP7zcyOXi/5Z9MplbgVnykNk0z/pN4SgzAPRs
1FdP9pogOJfuRERLBp4V1FDnyLL3a+a4UvInWyrUNqDcuOPzvqXQkJZhuMgsPSZgqwyBnwJaE5hv
ipvoeEAvWFp4+tghiDfX1jL/T/8E47JW1yM3fjMZDKd5l+H/xmUJQK3KhbIF+4c7/GX70L7yaOaR
ixPl4CPQH+e0gvo4iJN7YFtX9+wKqfIgSronn4P7BoSqUINQkr+y+81dCugPnIrRCczVhQTNhbC5
b7QS0YLRB+CTl2O8dN1Ge4yHswiAaX4QdnoMs1N+8LsgO1z6oGfbLIKvIWr5GXxPJfowkG9c6Jlh
9MhPjDmm7JcPP/PTFg2/HW3iICQVyzl0ktsEp6T2rRLwlO+60uplYWVQkcZBvFPhDSyKxLf3QY02
beydqwvPiczK5k7Z/B7J4y+7rVDX2xjw6+BNUiVjrA2QP9f+PcC6HQ6qVVNVvGLY8V0M0vPHxb36
mKr9yjXo/SlZIDFSGv/eoU7jVTf0Dy97VeQdv7ciH2kmh1e+Whm/U8ME7VUSFLsS4FrKvKCuhBen
afg2InpJU9sRbTt4o91M0R8SGdbJlOisv/AkVoBrwquimW0Z32xberTFwW51quCSmbS5cKxy5eML
dHy3TjgI+5yIlv2W9DdQHQ2CPxkiQc2DnqRtJe+Bb2IgLWaG3U35QRG64Yi9yojMfIW6HqcwpiM/
M3FzEdMMfhVT0Ub73X8p6oEk7Whwi7dCLMR18mL1PRZP5ZhXCykMFEoTM7D2SbMXdPrikhlCjWAz
vwxwTcesdg5/q62nQzxi9OYBdaAuV4aBAk+UBnIE5KZ3K7Rxm/OPdK5SiQowW1KEpJIXO9Y+BHO4
y7bYPQm3tHV2KszLFg88aYbET+PXtsE67HzifSXWYXopbXRxXLWK/5ZhM34RpOYpmouw/ShmGf2x
nc8dgvf/WPxkbgxcRbCcwl/73kTssyIVAlfbux7R5TvGx07p+e+v7Fta1ryzwcdLpYIzcGt4lkEJ
LOd202Pm7WSUJNqKwrygfzSk8GpRtNymkbu8Z63T7j6HNgMwvhDl7L+wDR7MpIUm2ve24PZfhF0B
43LEkADWAqFs/czV6SBYtjPsO/O8b6KfvkwJu+VL8+85kPp7de7KbetMZxLl1j0wFOj5SqELw5fG
E8KJ7d68Qz4c5ZRgMcMaDVTRkKII/c4XqChiJ6V441+Nd/DdjvFXbYQgYyKGYcsQBnRhazpt0EOF
o0UpWDjcMslaNKycNchA0VYdIg2/XWrl9BAEpn/6VfkW5uZsTMpydI06ixTohJoaX55rNcNF6M6Y
nSiTZiyeHONo03cz1Yer6gyPeTZvnLfn1vRxPcXd1gM2ya+oqOqe/ZjBmoPwmPQwzmMZYDoqB9i5
2JYOyzn+Hf78EE2bjbFpudop2c6nqbU6bhvGjC55jwXPlEdl46wcq5Zw+UVEENUQ7inG5JRT+oso
TrL5yD93ttforgMPTbKfSzVFM3ns+p5jEgeclDN3eWCvbSYpxpKCWsRN6BjoDYBpIMbHxcAs9Q04
mggRsCnnMlfObnwCtnRJweXzz6EDBBJW0uT3MOsaGmOwDXoDRWgF37xYaENqkCA/sDC6BXFmG6aB
LnH9SRqM7DaSm1oStoYRL+FR3/j2zygyrV2IjBPLw3+tKx87kpfuDDdP8MGkdfh+qvIYymyCs9qD
g3qy6FLpTOJjJYGUi3rO0SMrty+8T257F+YcSiLevnxSvTOuul41HStEFbprTsASBG+ETjpuPGZm
MZHJgvKopIv2DeOQppsk8ccF0LN/ggpA02euxXdipcjzE5aL5R8jMb6WpQUk6fiQhoxk0X5z9qCa
R48vgKqvMJyU/3oOgZAc48YLDlY8VI7DtAiAAhWV2vwmnZPp/m1n58/JfRnWGC+McnaB9KCDhP0v
XZp/9UH2h4p7XWgIwJwH2GzYA8LrGy2wcJcaT/GSbVvgwiuvLy4bPX5zsHzmufQK8eHtxkh+1982
ZC5tAbbJf8ZZXqVo3OSsrtxekn2FU4PRjPIIT6/ia3L6ucftMS/k0p5D6Yg03nnKB7ld9pB4TRsb
hwlQ4Cmq8iSKo2b0DKDf2Itnm+1ieZ1CwVtgvPfpB1c49a18rEnntQ28XH9M5oFCQkEU9bzqRF36
gWDkTsqORs8i6gdq5DSA2Mfzln0XR4NeLc8GoAXsJ/xgd5IyhFBywPaA6a/uLyA9QKjGNxwAAQ4h
Rn4uCCXrnlaljegHaVoHQJmyYmWHDeAyB5u1Yu8uFRQQxFQiW8guoy84Y+9p8dg7MoUHo2uFtIe/
tvTkM9o5MKiPzfBzE2lirFVfF0KvfHAl6PqPb58S3xcFRw5X1mAFG8k6M4qU1MWvISGVSRZe1/Nl
ITMfUylhA27tqRIvHeXCqeMbRqurvXASiXvWkiK5uMXZvO+TOoCgJFw4dLcsHPDyq3vnIR8Vl1K0
l+tGWPcQsynM6dAp7mPYSjZTfaqabZW3O/466GkxxVcZRDuEoBiyTQX+upB2TGd6Iq5E+ME6n4C9
2vYWaZlosyS/QheSlhxLm62IMbJz+zudBRpOIedHqsP6MWCAqqBMw9r0qIljY148mMlKVw+EoNil
tb3NJqYHXHdz1Sv3CTUJBoLHpXoGxz3lJTaFwMcPlHbQJ7tGUN1fMGp8wMdu7CjgxkydjX6nfPVg
AYE6ygMqQLtHImFoYpjReVGEiqGbNxLGd4dddpgxzlb59g+azwOJGHzO03tVa1Ss0x7IeU1O/kla
UYrzYIEL8H+XZIr6z2mugYMQlJBDwSEsbY75RXzncA+33qGEk+oPlANKWxc8JQ5kL5OenEuVP8cd
98/L28eI8Trt9tGzXE5OjhHr3qgqtl6Uc+svJ++zbwRIOUv0rd5J3TAVZGfItTIcZC8l8DGvAh5U
+iUL5taTzbCkgbXxXcY9wgaT9gjS+nTIDcSDnUvCKY1nFZgQ3kQlLWNJQyv24Fo/Feb2f8V97xmW
p9N99wKbhp56TRU1OArv2HoyErVS1p0jZXWW+VyO2DeTJxfLPF1rQs6r3iqL3npVR/8SogALcVRp
ZiOGCR5WO+b6vzlYZb2MqBNEpYST5JrLQ9X4tgPdyfgVRe+wTVhz4dEAKP5c87ERQf44jw/6Fuk9
03taAuygppGbxoC60kAQ1FYo0U5oDWW/h5G7Qq5iKoT3hX4wR2FjaqMnldSKOTMIbU4IGcEqZ88e
yEPJQepr9vR1sOFkZoyMG5RiBLl8PSN6xD77H5Rkz+HtA+AUHL8A/M3iOT9cDGADIPemgqCVShwt
8YkK3LzUX87/fnnJJ5MADta/x0HtYI4fuoBIer0srVcADdsr7+ssrhxhnBuwCEigAqO9oU0VBQoO
PUcfMDs9zAkSEi2ToLFzotpsFyb6sgy3dIQ12el69SVFSdEF+MjU0S5dIVh+YjLZC8xWy9xKwP0c
wmfoWkZmFgeHJiHRn4oRdJAQ8/UTqeJhQE+hL0LswlqrJjF5E9k+QonztYb2aIWUDhobSinDLQBZ
5T3LOTRQ4aXHXm2LlxJR7yUBD1ufLDiNlPMbr3J1w/JfOdH/vO858DKtDZX9icBakYAmMsrTM61y
C7e8v8THVmgKPB1DF78Q4IXJ2dc8YID911bfwbGHBzOJVIdloaiIKgtNd6BUYraOfpUaXbdGp9hm
EaSTdcteJBzrCLCvbJySpJi4eo2QXeT7Zier9hlIafIP8jGkdRbCfwtZDogrqRjQt0mfb3hyF+Wr
N+gvL7ggwZx8EOjycAqzQfKEOU6+nXgSCNQsB9rqSuLhtvS4xCNahz9Ni2wEp0HKuMrsbpPhr9Gr
gmYgjSbJz1svq2BbCMpN8R2f7lB38epMp6IC3XN9f9V/GhevOY8nKkBXHD5Vrn+Gn3XlvhCVeiir
2CodjKgRqt2KVgJAZzw1ZArGl7IwYbN/KM4422+4/Jq9wCMSWlyaXc2ih2MXNokLZawstI0tuVEN
zg6E7pKl1tOsyNjtmPLU4Ya/8IpFlx+zoB7mG5Ox6fZeuENEaU/ttE/BWNPPif5RBCsG3Wz4uE4D
0Z1y5getFjIfwEAFZVU0dxV3aY1V7+DhER+bYt8s9jd9nxpx7Vnr3CYM/X6dTkb1v5wvlteUh/OS
xZf0sBP9SzWpvBsxjVOun6ur6lu0J5Y7rYIRDm6uhu+ETFsAgMymUGrl6U4doXUQrc+VnbJ3ocTf
bTttlgICOGmG2Nk1SLzhtE7xD4O5KlsYNaSohwztKgafjLgcvPvdRtbWpvWD4vfxVODB2hCR28/Y
rsbcchEA7IMjQC/CoR9cONWRB3so3u9P16zxpbfSxeUvOaER7qAce8XnWGV0c/TCZcZmStK+Z1ig
ZckzEjFnemPKM9sXb2t3jU+E2SF33L3g6LOljcJnJDcyxAwOq9fdwWx8P7iEthhOwkPNBlvRHTmV
6lSWOfIDWfcIkSZx4D5cIFy2IKquHK4tF7qJ4cs2RrIPLTI9pAIUPfFdLGxs8rHK4AE58NM6KxM5
DEQ9aoDEwSvlttVii5KS2bcFz41eQGPoYFPt50PIL//SJCV/rdXyESAriJZDLMxFO3v3tQhj5pq7
XO/a+FIqZ9lNi2HjnmgdyawVTl6H4ey2zH7puXw7xcq7XvM7HnbZv2IOXV+SIcE7XKHXqqrEcrQH
5iFZz3nIiL1cwCOpOR7bzp30B5Hv7NqNVGbSZ5qCUcOjBNLJA+sAjGwaiHr6aApZTheHO7tosGqe
X7s6ntF+MIwLYlk1twA4V6tYR8Re6wPVE2VZ2V+EFCUH2rKYgiEq8K7/yGGjhBOL1ctK96l4mY2K
a7VMYXN9TOCSvlEBSuXdd4QLGRwvrCFqtG15RH4bSDnMxaPcioDWISDoJ4n2/VbJghrwElP/eTcL
DkVgV9IIJ749HSX2vI7xk0qpIAsnJp2A+mtOp08aPZQhvkY/5aQ3htEfUzvzMg49EhMQ53mIlQGk
IF/IjzWL5lwpZRtHbmT4po4Hdtv7+VNOQDzHwwnEB4jQuhmNKB7U3bygYorOdQA/EzqhWOdW/TLT
GkrHvNNbLNFmWHC0hnZAQk1slgKVU/vjtfl9W+WLVMOn0+5NtfsnOeGk8Ls5L0Y68IqgsSDdPdqd
OVngz//dHlW6C2+6BXuBtM+kM5MCd2bKNnrF0LBFGZtSYg5W5JxxPyLbIQxY6gr48CIp6eFFXpmu
f0nC3QnE+Ft5FkMLKcIB3p2rE2M8Aw6kYQfNSsNtpT9xxexv0PMjF2vomFl6P5jqGzB5XY1O6TV3
tRIYikhKPTpmqqO6z+OjCUrS8JHa4wkxEyJChT9Wy662m/4FpN09uUyI8zqzKpqGmQ8fjK48pt59
5cAWQ+3xyctVuWSJj3fC9jzUL5UvRt3+97G6fQ09AqWcO59gQpgTPQM2j+JD+6p0/Vqb3+ERqlut
GoVTcT5jAbxbnWtwYKbJRIMt23yhxOmRpDL9AWZC8J3aWqHaGYRMvpIbcvF2vh4PRAGColDinVXq
AotfpSs/xhrZT1GlraNLQNkEbxgnX1s9YMq6FvqesFOZPPmoBt6M6HhpDLWyT/FBCZfWzk9ayYb9
pY37ruaQPW42nGqSI7U7kKk5lfRYWOLJ2+jBY82cPeP48UXUPbhqKqKJ80zYPqA0mJfWK8ZFJ0WF
6zjHdfapOnZ2duu328R6U2DUQ/pxYET0Re1D6YemcYj+fVDzhJvG4Xsajo8gjrSYsoOgRXC1/T/P
yWc3+XtVY5BWO6NNt9cebr8He2Q4o9FYZLxFGGImiLDqjf0KNP8agI/at5A6Lti634GxQPe+p1ot
VzRb00NGIPgjoMLnFcgbpHRu1GUG1DwYDrL3wZv3jcMHYFygXwYYp/kZ5MnUpGlE/vvOWeVHOKs5
iB0f3CR9nu3wsUtn3tFDUx+PAJIqc7PGSqqVtdiH/leYaCgPt8IcqxrQO7g/aVBR7xKnfPOS6Njx
vmBDGWNB2nIfIRLZhLNkuo3WRmBv4QV5vZ89IgYtCOD9Apx5PQqqPiDdGEqYs8BrEnPtkLu1V+31
wKygEOeUvnjsMLRxOPNiTgy46s51RdifPddM/Fw3m2H0LZ3eemM75WPJGpGFXCRLOw0qkJP2xHF0
MFmlE+51oU51UIcJ7JqV0MJPLZ1iXDv7qIRzZ3wUezmPpl+ayekMSsSq9pTgqtAhIZtgWyDIEDsC
tySq+6L5Vg0m0HJMmX3bwjp0AQfBkTdfY0IaQ39IiiatZDGujTsEH3dT0yZIKU9eElclvgL1bech
4MYoMjurbVMTH57tlfdHjFUKVIG+0YGnF8LIVUABawbn2v2gzVgO0w7HbcEdNNUSfIrzRwMo1IcY
80Z/9Rw2T67ikNnYnI06Lt21hGMtLS+viJ31HpPuLWDd0HTt7yY5/ghPwoVpC/QxXn2teZbEf724
rtN2QDq4sQzKahvMd0Z2HN/uhg8H+Ic5WtGVp56jMulfTrZ8MDtcut3TpAynKHEtHg9pHqx9PqeR
Ititk22KoMh9x/8kQncDYcHfwW3ixzCxWjUVyb9YdkUOMOKYWZPtWMzxW/qrG/NdcYfGKjaGtkd3
3Mkied81ZGidAnGYxMG0ezZbfFXOrY8iAnzhQhnEzFVv706EydPsjxwNSWVa2LPlVPBiV82SJUKc
lW0q3LaJjp8mKIhkgH8ViDFGX4QSWMHNPnthdeNBJvbKbdkSb5oPoZ02WLaOnlQ2AE1yiBqhOhqo
2gPhRLUqLMy6jOZfX/cexWSfQBLz3kn1WE8F0kAzz/mMoXY+TeJl9DoHHI+y1fOovZSHxzA65IQl
mFlqoHk3FWEOOSGqDlgVqeGYtKf+gf3+y8diEY8bp4x5IqaJ6AQP9J4Gc7xH9UFEjzyBauUirIXh
jskjqGxV85N+1BXKX1X1ysO+0F0gdvbafW8HNaXJNgGZQZRmXQTiyYSqP0XJru9Q0DRXz5LYuKIP
11wxG/LnTbEZs0QAlUt7/p6hvTobxEdEuE1fZTqlacZ7wm9bL32dItC4LIdIzESU6OujvCgn9W1e
4Pns0navCvXHp89DjjNPY+Qrme3WeHreVcr10edTBPqYdT5l8YTAnKx1ButlUJ3jIRKoxeCNp6Rm
tKKp2jDly4VvN34nr5yvSgzQqydhxGNVq41NuyNkqmluDIDKr5cB6feOCFX7ewfus8MCnmrTnsMG
SjjYuW1e/GA8kW5EVNNbUi47DDNdQ7GiH5Sule1T68Rfn+T/3uvASlY34CwHZg0VasLvu+hs5aI9
mMWBb9EG0y5JCYzB0fso8mkXiNOHVb3WYSBWnj9hcnEDc6odh4TnNS41/yVCzd3JmsCLRLSetfcM
5yB45HUX/Zqg/5+XEe8O26730H4ljg7Sd5gVU12GFgdJVB3b/BYgS+T7wfX4DAXEfTBCNwHMT2Id
Xw3qkcjkxMob9qUgmM+7OkMTQ5aAfwuCePycr6U9ndLSETl+hyB+i0T/yOeoUvD0oTHJfjTMrCdj
KsH+BfRlIGiSVGsg6qYXo+UnziT6luz2vr0tQhnGbMxhkeWrr5hJ8KhlwRMXfBFaVIKBrPPnAsJi
chXZUHkOI/NlV/yZ3becStQhf5hTDbXcM0zVgwXKoLiLdEO/u4wJ6lLRUyqTcytA5uIeevd9mfJK
anEhplKJwymOrC9fXQH0O80MGdLdNfNGMDJ1EPL8wAAY6ph48AsEhdl/QsUF/sOiX0WjKiS96usG
GxwAB4BqCZnvlLOYSol9rHahRuf2gyDVrA/AF0aJ0DlnjBpZ4QrYduFPHbKK5aOtL2LpttgbhnUJ
nsO9XDRkirRoEtEMQCi8nn3ELh2cqy+VIVcmUmE4oQQ1NIhS580+ajmyMhbfsoIQxNLWRzqOqR5c
AVV8kdGGo1xBX8XVlauX1xKk3Jc0kBhS8Ns6Ir45CCMATl6D39HJ8sj77XVnRFanZh7Mk2A7CIY3
dL0+1yRZgiHv2K58JFXkFxJ1VKVzKKzxlIjokJpbrcAFH9CDb1ZlFfZrzz5ErMq/kjTZoZsw5h1J
IMpMZvNE1991p5rT7+Rbx41hxxmWyViF8UiArhbPvw5MmhgMPB0XSZjuJxpnWoP61Z9mdiLVVbTy
8U5mHlaFDowq8QSSeNFK7rhZ7tkOMrcQ+SGIgU8d0Wqi2gVvuzJhnWTdhW1AXOE+kOx82DCt/6AK
TpSAP2qIuNQ/TfyAtsSIRF/x9iqW86aKkb8ouMjuSflWmAEETMnPMOOInk0lkD0QyZgPuWJ9Ng6l
yWXIRf8PVPMHObSx6hKOsg+pnM6hWOclJfhDj6Hi3bM37C+xrkuBagQ1+pOoBRgTTr5SxpThxfl+
huCHKEoh6mWzMSuNfaqQh8DGfakYfy2jw4vlMzXrK+2DS6Iq5t/epkh0UUw0gJt8TJbsmchyhgFJ
OVSt1+IZVfplPZJtPTB+yn02Ob2V/zDtD+ae70cYhj66XDHdEugF9asUXQucJ9+lNQx6QV9PMLVx
QYH+12JzyPGDJevue5ieaBqJPucUajOPKYANxyIUhC2+8+FwezMjEfeuJNOvT6rMF0Z+//WtRlCZ
fDvZS5szvVYZvf6oULV7DS+qUByz33ZhkljD1EPWy+YKsox7kfPPouluz/G79ASOMMa+omZUsX2I
Z/tFnTyYDanKhCdeqp6JC+0RbTVXbJjAvwpGl1F5kZFrO4R93M7lBagw/zGJqUtKJcFNkGlwkg+k
g0BPGv9O8PaqKlvIDh0/6C4JdpCNDmd4I9WCsYt0dlyViuujxU25oBoGCQpVVy5eWxWk3y8pxO2a
4jv/2pt673XdRNtNVTXD5aetHkaLu8X03LETC7JUaeh3LrKrA56AXeD89sXbMXuDD05HPVD4jPub
MWLug/luJpqcG/0bhQT4rjPUUS3iiQVVjmy2a3zXlmAa1vyEzurs9IgB2/K//Rl0sJJRcqcc2PSk
OwA88+egoVsPCpjKnqtsZQR85CD0mOwXXm0KAAGzOS9OtX2Z0kU516cgY9djlyNa2MEYCJxTmjSs
RkAI9euAw8wVo4cUuMFG648ReX9HXd2VGj26VhNy+X3S8pygzSg/I9jMnh0NdxkJZq9zbunSwvKE
EEH5GGf2IOXaIyalP8dLC4mCpALj3qF/4Nj+XOnfW5PdERwX0mPrDzBRBOpsI31f9WWUiD6F44JF
dfTD/0Ry+tT1L2v2fgfyGgIC6a37TZ4n1uuIwWKLM0XcPWVOfu1FTPgmkLyJovQNSEBPqTjLaDzw
QSHZPSb+4K0zCXSyig4X4Tcrg0Xdbfk6VlUR5dk4XnVRU6kZx04WJUMYhkXrAE1FrizydRFp/LUs
RNQ1MlURc4v78Cm1v/vIFda4DZEdV2S3e8s9HHMRJvLP/4RIJuN1iXJLohHZOYjXioYkpmXnL1iF
0q4Mgd59svWNE6X3FK3m7GrCNssejI8mDjX4L0nQy0y/oqMt5Agxo+FDD3+F8dVsK7gDM1f1edu+
/BMIhjSFn+uqhI01s+6q7grlUTYxLFaSq8GkLfDkb4wEr2hbk4csO7dqkNes0QyWCCNMKUiD31i7
cL7RITU64OzKdhX7Letd+dVWui/MccbTwlbqld/0h+inFayz08rfqERNzvSmYZYjjl+vxDeSlVGE
/FlZrmAmK7QD9CDdBmSyKmCmXlZUdRzi+QiUY0WQx8edhbAZ5EuGbvH6HAt18X6uPCtzDyrKuWbD
KtGEmfrBjPRg3vOxJkCIj/SBbCtFodHErHrsqOcgDmgYm0hSslH8uJBbfoXlDsJT+PfDX8+nK535
lSj5MJOVytlEIblhzfrX17FPpFEwxDVjeQRsZm2GgXe9V9rkDb46GX49HiGd5LdJmEwZ3yTrz02T
r8VuAHIfvowroXlmYDLYXviQtCWyFFFKk0a7eLCtW1zYY1BTQTMxdHMGA8ARztoTV1r7DRVuzHZm
y1ljzlKtcBUlkRy7wT9Lr7T8Tbq3P3BsCtvJlOS9M3Yg81T4PtrpFtoAoavusO4U8IIs/k+S2LTT
S0z49340CNawhqm0WruAv2JYUmlDOdF5hXMDLgo7tlZ9zLPI4NJKMa51IwLEdySLIvQB5BTQeGHi
8eYN3PCE10JujeuysYD0CB1DPoGrYNKh9G2R+KBqdBatFvIHznWmW4ednL73OjcJDgh4zIwiKPR9
HvH5uvna8vj9WFEJIgzVTBdTk1eTJaKCA7SDBC7sPOULTyGbb4oguH25CxSYrZhhjpkU1UKZDkLa
QuP4u+FV1rYAlNdddzpGZD2aBp6WSGYNulaRFqDFxHAE3TvZN3yweAjPYlFtdJ0BPCgKbKaFqrfQ
9J3fRr0zYp9jDRXvwe2x/U3MC4z3T/NBT/PNkLGAtbcqilNsGaDHCuhjbsY56gHcR9ZwQEf5WO9Y
/u3RGvngQzGvYzVtOBtgPZ+j7rFYoWMeY5M0p/zIJFkspUUDxFJ8M6usKx7wMdXKo6WAxa23Kju5
QVLC6JY5ssZSwYcWstImbrImnZL5afaziipKF8uXvPNxj1J8tYO5RXDHu1jRqjZxM1rYkUkYxLpW
KEiQ5wePvDauiSWnauGwIRstEvbcKd7hG5Xz9/fDR8yMYX1pP4hryusApS0yIsndZ8a7VHy3kAkr
6JWidqejdqJXBxJzyV7cSZL7np1FaV6TriErS0Nn9twJqNtAx4C0zt932Qr6Jr0vwt6HCW6CPCUG
HVBeIxoQ8iGWF5I1WQfaMjCEPfQWw81J8XgL/HyycCWs7ceCgsepOzUYC9BZ9zMPbDfdYKbku/kH
yP5ikG+YH+f2u6rY9OAnjsovNnN5keywnrSt4Fvgb9o1gz0zOlTbJk7eJQft4jMIlln5Ug0trP7j
eItLEt88NhF3v5h0IaZIRDOUOK96REfozr2oAOj6JQLvQwqSQXAfuyhkP97TMGzyTuD4MIxR7KCp
ehQfi3E2ntZhK3Yl4JcVk9gAwciShLrwSxv6LrjmrTOlLMHjlcgxvS3y0WrVvUinTPwMRha7ODBr
8SNRaEYPlSO5e+m+n3zg0Xq9dQIcKXXuHyX1jImAqnKCvAQzArLpOZmXbzLla4nbMevjg0Fm+ZBL
Y2lHtdYcyuBn/GbNrNEvUMrkc8DveDftbMJ2ZL0J0IWW4dLKpiFVwa0cbzNj/sCc72x1j3bTGUc5
idLFS8LUZtUN46ayxW9RjJbwNEk2ENDjcq4Gc/KUZ9k5ukENt4Ozd1H1ROwdgHNK5Dd1B3s+Psvq
H0n/suUvwLQO1ySNepMzD2e2enZBQa39jv7Vf16V3PTbzh1PO1d0vNSNrSsgYtXsbfc24VoEEito
xxmK0HNetd5d9gvqrAWUj1e+849H0vdf+pZFuH7GWB+h44JmMrj/biDs7JKni0E6ypgpK1OcXqzj
0X/bRpV+RTB2Tv2ppJbikwZnlWAfyMZ+FjGU5jfbYCr0yI8IJuzS0LP7/16F2ALgBZRq15MEtzWA
2w6SWUlK15Zka+/VvVLr6I8a/ofr3iQlZmrVW+8cPq8wgCFBJ8L8PpeC9i4kNKuqiRsDXmWCMBWS
ii3pr41+TwE7nsbSBF72ob+Lg7urizQQvzV1vAJNPJZkVkUvyMwQ/003FX3Whk4oWmCT0NTtD+SG
JGIdelMlmiV+i1AXEja5wS16zOPLbWmw48JVZItqM6USrQtOWtvJTksyQxU223NGtbChiy8HLDHF
7E+TfvlUNRwAVk/uZ23UbTQ2eHXy+GhGUiBzTlq6NvhQvVlo9RwPNmQrvgDWqxBI4QpC2gEJe3C8
+L0H5kbX2V60quDtkwDmHxs4zztQZc7+E00VTSf0N1PRNt6UsDPYjnoo0pw6gBUJ4v12svPagcnp
HaCU86/j3qqrd9vwTFVAoQ6Bp3r5WbDVoO7kvDPEpI/d683RFbu2e7yQ7EztNTdHIBmRqc5QpS3o
6e4SSouehQl7tvpxBErzpw8nmrKYM9lM5gbHMR1LO0zTBuY5E9Yg9cQgXSeXZVD9pteaU7KhLKrt
2IV00iNSlt+dm1pb+3SPCyXUuUntBzq8/SLkbytvufD4kw8bUS3tDV/wLYnJAqA49vOV0anFUg3V
JwAgBBDibWIYWdRkePRpULe1hedaFoxfw0nyU+X9IDLt5Gg9hhmP1tGt30D0gDp3LOZFXmrinOJe
DA4WFXdgDIYEldkpJmEZ2ry6EdFvfL9sd+N4fOnL6L5U5cD6Ke7Q+E4Z1dJ94YhS+2tXlx/l9J36
FLNbPMOeFlpRuHtAkcAL8c4B93XOsz5+cgTS58wyKCcTAG4lsysUtibCkDcnCkwEV6zVO8izQnuD
/xR0buJmvX4uyWpfuwyPQHEjYSsozui9icZ2g8JBqp8XJ6kCiMGGjSA8CoeGfXhutBMiVapbzZUu
6w4JXZ9W+tAm4XCeiTbf1p5s3ypRtkqlrAv4skkqKpIyT2ycDrFdZEgTz5uWwU88fW6DnjlKdgFo
awSdiHK7rUEwCl/PL1a0X+9BXUagr74wwB/EE6hKwjNAR8s0qTnIeIUsp1NBoHGBFoTF1spTwxwu
HkqJPI+mV7zZrAtkKRKW8k0qrJIr5PZoUkvZwp1hDTjuUJGT6Qc3gwBFTTUrMXR8QQKI/NW8oB5U
1l72SJDMVKYBXxusqsG9pLhGjlTgV2fV+FBJ6vIDaM8xOSY6TODCnFO2QJpcS9C+okXafyaHDc5t
ECRykwmEuA9CD5nlyAiDuQcE4ZOuUOV0lzxsp75KxX9gTV+exFFQvbMyIcUEJ8L/yEmP8YJSbF90
N/Bmj2snRenRc3nZ+DHjbZJPYQBrKBmZwOiFACHDLefdUjRMo1tYFyM7ZEsFUJLM38V1FE6Qs5gF
X9w5T3rgeW5dSlqCCfjQhvK/uFB2Tx9JwN/6chjAYAU40LdOgXisGiecqhydDCzzkXyhfeLZuNHv
dyqUajjwdSMeslPkX8FUifRgGpyaA8rNf7sPpTo6Q65mjv7ApEehLTaKI7SFIqhIs/514XfJrISx
CUcJIPCENK++KZUCc6eR29uO7XzDWdE5FvO1Zoa0WS4KKV0KNLnKvXPAT8oTfcKtJofPkvT7WHk7
MH7JIaZLQzM87ZOdiYP0Atix+Lo5qT90WKNlFpurgM8UcSborXci62AAQTHTZx3/TSOOXPosx3jt
+bhhitFqI3WqmEmZ4iWSp72SulZcWt7CQn6r3qP27oMvDf6IlIQgfQBdm17peb1/BKqUHKkLIP1S
sIGfKB0oqAiqStkvwZQty1TJ0DWVUvilgGu7skAYFu+VpdpQGspJwX3AwA+f5ccD/xmPmAxZI0gr
BwA8wC2AMn/5GK/QOBoiDqXMfl+Q7t7iz59UEoRfxhVbhSEUEZy7IgFpIuSeW0l+bf+A64qY5G0S
KXksVB7kl02wQgc16Ss23j8vkfNx1tjcl13+zA5Zk6W+siDHrV4BVy9NwYj2J1+mZcMmGpRgZU1L
AQUbuvB7Mm/wsY5VMNlxb9pBvLPIaCslrnaaGqZ0quXpPmaTY98M/XnfCa9tJL0PTe86oAEAWt+A
awdi613MKFKuo9Ys+ptxPwtND7UoO6K1sILf4PZTPzwgNNWGFOlD3XbYf+yxkESg+mkIO3gXg/Wa
tVNPDXcmpEfY43+NSf98S+NflB71M+C46YcfRb7idEHU161F1AMm1h1Ugsf94RAMda4hz7xY4D8c
mfPRBbKHSOrbt3Izk3L8fgbIDhre0MfSNExF+O9yBsCN0uGzz8WjRCKBu/aLlrkuNHbb6U+l4vPZ
sV9Zau954YJANxCwPkEzibWRXbSexiXdlaL8e2wxI8hSnFr1S7KvLnsIi5nduf0sX1yWGwm3xv9j
dlPgaI8sm0g7wXCqi+RO1buKDySHj+kQ9LP+iWe1C/+9N6ZLJHFGfz4FT48cIPN5bMFvuVR53PKm
lJAMmoNnbK0dgPv8aLdubgguCZL58kXiNSVxIfpcwiA5ovw5oupx59xiQf3ET7IFn47zl38c7LvU
JbiINj31Mo8Veed3AQGDl72Rf1DiiWM9Mwlimew+YEotb5WEJab1EbrZgG7Wzzgz/ufTPzY2njU6
7IAdpd9G/IgjYFivRY6KsmXN23YL5apGE5h6QJ13VUUbAxkhI75+DrUOJ2OE9/gKkPeIRQvdaTsh
Wv2NsuXB6ah3QUKUHi4OWZ1BxdEoOhx1AQVxwXIwktjCmfIC4QfDksycaECqfx/QLrnESklmbZAN
fMWRe0dg6r8yBPIKJ5mRf1Swq7qKEEQwCk/d1xTEvKAYMGvV0xvzzasuRYMN8haLlNoijNBfEIMg
BXaxJ4nLF8kQz4v2cYcM14sFu/k2TYDJn082vub8Dk/lCEiGI41Hl9fPj6kOH1/bWDpYtCmSxmio
3sKpZpv14m4f1D7LWfg5k0mDEjI/77DwLro1J6Jut7odWNLKZBpixDjAFX/8m27D+idmDHGnNqrl
aAWTUV+0RQ27URooGLeVI6gCLqr0pBsC2gD8RkjjtJStR3hhTo97YIV1zEv+20PxvtNBhBRJ9JDJ
K4bAfnY/cncvo7k3+TkXOp4GDdQT6EybFvzxqto/smbwKx5XKr7vlm+OPDM8k1IGTvUoCLTwLPjh
1zebEb5IyMdmQOwC2rERCINBNu70tSaiiDtEibGxkjpgwIgyQt5EZuHZZ0mAPST2DYtfv/D1FYO8
ezA+TTPKK47GTii0B8Qi1NoEQnfs7qDD9n+7IWSES0d2+Plunc1so01Ij7wL1nuPIRQT/7jQ1shp
V2K4Xe5G3fs4Bhb2FUSTyhBqLXF7HCzs3lN8JYvtR0+xxOznPN9yY/q9zUbaqcaLUnPGQYmrsC3R
drWPsVqZan41L8MPTyJES/35MXjYKflWbEc8au9ysVgLG8e9PfDeBaQ/Tbxn2EyFmndS8zZuPORq
440tpK4ixVOSu1iNZelOHBZtxSHUdrYf74XSNvq54cErwOTMYyCsLhslu0gnD+ah3tjqpK7xpmjS
Bveu4/08sSu0hHzKdiwT3frkqhSpF5tRtj5vVMX4PYlp7iyopD0uauiMC6muL0hYsCyeOuLTX5sm
a8pGp+dagMMAuV/uUD3gdnnXaLQ2BHUjgrk3yQkIN0ui7WQaxE9svuWbTk2oeaV/KRTXGbgdZe4C
SRXEkM+5Yu12+q+us0bTNjkXRtr7zzjeHjy+g+bCGMAZsh05cl+aBmK8nU0+2pCy9MP4+ysoSLEu
djq7gbMCZwRk4bFkwA33mA2h/3PCbpEJMa8kmpQillRXQtbgtG1tA7ccrS07Jl1bVqtFKOXHru5y
2Pl/E0iLxdMT/mQ31EZyimKsFfpdMvy4hrDXu9HmMoDuvGWB1yNJgOeH8oA0tNChR0S1BpzrpWnT
T2Kgg7FJvOI8mY6KXvtNLkogTTubEF22InLwLq+2oCb8Axy6TBw1/notigUTQr2+QC2tTmPqLm9F
yTOGOK461NL9wcC3kfSaMUgxRJLulrrjPZyLEMPerm7ax1SBIrOJ2OTy7KypLUBgfbzA0eoWJ3rZ
QsZUBXy98o1y3aK1Hj6deZSsnhihedR4jufo4g5Hnu9wq+y6amoc358CKrZtf58VgeY+9wh2zb8q
6ZiIDD3acylC6+0/h+WafE7lYMwiuwL9Wa+FFYxtrr6qT1wQaggqWg61cDI7rdFXs4NF07/wc6U0
Kw2xqhGB1TE+Eb1XnsXynaLPfkMjW5mUgQj7IB36zfYYtZcpdkzRK13M227XDyQ+fUNskzCN8+wr
JM3fgUwi58Nf4WBUgXY/iJuQlfiwMqoiiWNzhlUuwkgYcvBiYVh7QNFNh/ZUKfiSYYXZFoh0SaqC
R088P+wrQ9Au4B7YGY6QnVVUCpss7zZSJfY2wvzTs4U5trQuJmf9SPxHxRU5Bs2hM0xlgw0hZy74
DMuTLirXFqj0yQkty5re78XCBHAtox6IKM96hDi0w2/E5g981zlSjVpMClLFFT9CyH9JQZ5kmBzu
0U7xwGUU3LB5M4lqddq38LTwmgtumWCMzmzBDzHThz3+25PqwRS5b6FXHbmoPrvTkT+ebmZX4zTI
VHAiFW6PRiSEEVF40Ezg9oVpg/H2zul+04iN558mvKM6poT23ov/fT+L44vtvVserK3dwUpvV8+l
2rjMWnyQ37d1y+EB6R19xlIgg1fCnAqFVneuCon6sLr00CLXCYMVjDZoUFz70VHnuNjuSnNhcuZf
rZ/ft6q1FCt60I9R8wqti51+lP+n8M7cYyD2EhjSyR+D+2IajspVSXdYnTclFt5EA9WGsO6vIYf7
lCe5ABaloMxlP3HTYzS40O9rQAFFrEzlDyHcc9H9/q51CeN47lJrPBKNDBb2Mxn2UZEgY3//V+e3
UedVlVxRSrUpSbFjSGa+h+pfiptrzo1KIXxDae6rsjForLZHQwrCT6WQPOZ+XEJhScSuT2XDFkkI
tK8Eo2lun1E4Pu5XIRRE51cvTFXecjCOvxNEJOJIrYWveF5fQQvgFB45wo8O3EuMCO5WHwT8jVcv
79qnwsi0gh+TXID/We2i7xd16sHcExANX33K7T5TgDp5aF354JG2IEgKTrc+6EjSJn0vHRubM4M/
p4+qd8Ufp+eHJkgtrRlra5gz3+RHuGnGEX49Ko4/hrxAVq8xDV6ugZIEgyGtdyF++4gZ/wZpyygU
5OR8+mWQu/eqxGL3Hha5a240THzxBQIz2j9XzSGlu1govX7kEukKE+JdfcNLF6gRmOXj9FUyR7dT
odkYWkieoKryXKh7U0XpHBWx7j0o4cCVcUjVFGcsat16nLL5NGzW5jQuhaN1XNK7xxEW+YvnI7L2
Gyr10yKidyBTVwGWjlcFbDY6C+ui1siTzmSLssWTTTCsf0F2r3D6z2ftFw1jze4kVwHN23GvYCdx
H7dI08qnxiFAptykcVwV38KfwTJpeCiIIuCwcBVfi6ENKOMGGCnXpVyFxnkVAGqmk9wmIQel6SEB
5HwIVLEGdXU+oc0IBrNAh6XZiu1YmhoEyGoXAEvAam8oCZR3EVq4/LRNkoY7/AAwzXQyzdQuT+av
j5LrpRC7XWTO/QArO4k0phJuLpARBAi3YmRzyaxG2iEvdmtWYN90myG/+qQUXit1ac/EbP4MGPN5
mZv03z3xERzN714ZKq/4wVXCmkHIP2oz0NJ+6o5RJc1LYygTQJzyx4ErgLCYZdlezxUNdCA0o761
zDAB9ZBp4sdOkoES1uOYVyI9HjIhxPoBRcTeTJBNZaKkkjqwcQ8nUFQBI9RbCXbyNOx2A+TzocIx
PulHjtdEAE9xX6RHcYxrP0CVyXi9iNfxfWp8cIrkIXZceD0DXWsZSANKzFrPLS5tRK4X8ZNe398E
UgAnVDmpc+zrYRpK6PTca43MA+/WQ2ZcLQBvo4FZOVDfo/TE02MVNo7XXE+DbHZXnh/sfIRo8q40
ZAOcdPIrBHJRZ0HxQBhVsUk/4yakt9PqL2Ms9KV2bCBD8xbtNIC07z8aktScnd88czmfgdcZmMoa
3+TmImLcyiOw6p82v/RrLMtKStTfooSSqdVkg6foBod+wS+C7zoFLkQzPTzecpuumQfo3obPfhk+
4V9JUyEm1YRVUXVcFmc5ammrVC8OhAHaaaWQ/AXxgYpbtPYewPBuRGQvM+RwT7i6zq8bmovAPsl5
bekpaohHh5q7wLwsPzK7HkdGexkQ0CKxz9PujnyvIREWsW1FaygQHwU3itw3ocZuQVQ2aRyn0p4Q
SrxI/Khl0aIspMeJ0GCmQMmUzq/1bSaW7b/9GNzU9tq5keWt2mk9v01V74atZ3UcWp8XFMnYIj0z
fi1/44mO5ufZEhXmRT0WRrgD/hJKtlqYFfFJ+B+AiHSnTPY9I5uh8sze8l2ykLCqmtV1paGtCs5E
8ny8hzTw1jy96uR1YXeWbpu0wykjH0I4SiAf0Yx9803AcOtJH/qfmpmbZjR4NcNwmSQSROS3kWbb
DU5RGuCjlZpFpszlVG3X1AECCts+ZrPi4togKRtzwGxZ0HgjHa6rjzHYvXYX0DWF9v4c0GAsS/LZ
wfAR60QYI013CmINjUcX5vtgSHzK2m8EOL9zCtH1V3uFNfoN9jy6v3srEwU6wojrUnnk6me3rTGQ
OCM6di7Hs9OAf4adfgKNzAeHymtzAHQLvS+FRn9KOxepeamllVpAgaEXPn3lekywwUo90NrAbcYO
HUo8HVJ9qY2HmXLJKkM2lV9xXngrSSeMf6KUr5u5e7xveRcB/58rBdZv/XgULKUp3EsEFiw8o21H
XAYC5WK+aF6JnYOEtMizAgiuQNGSeV3tlIQZpM0Zuqsr/I1d5/wIpAat6tpB9JKw+wGxjLVSCb/+
PMBoliF4U1tcynLNJjzOKsN2LsmaWZmZOAYtx/9K6P6Ltq8uymZbUjmsgJNwrjzcou5gz0knQgd5
Nma0JcgHbZLmWst6HWAWEMkjRDasAWotcVDvqr4G9g7CyWuzcQSLpXaAhOGUK9Ymu26lGRcRzswl
20E2S7HwOpgLHLTUNhp8q34u+h4Pnb4//NmygXpzRqSXz/jZLmht2RToIcccDGVUp/1wBIueQ3qD
p1wTm1KDmtOVkQn3HDm5ZaYnTUGSVu/30gUtbESH0D4ZpSGut2aDfI4Hzi1KIxEAB0sXmy2Fv0eD
ZCSD7ao3XqeNTa1xmgBl0kxB+G9SptN3cE6wr8NW3aHeaKm9Qo+McUdLVS/mswFp8CQTyIC+VUDB
ZqGX6nCgXiAKIlShxRVbIFr/aZLjrwr9LVlfZED4aGgHvAv2SvYA47d0MsFAtePRLJfd+U3Fe+Si
GoIVzmTgolTew9avfYee53q1+ouEQPAcyHXF0M6gpsvGNRE5C466RXrouR7yom3ejaCSjJAQCYmu
hmP+8RiEd6lPM5vRUKrF5BiQMkh4PeeapsIG7Gx4tKQnc2l/l/aICoYW7Bt//LT9CFg7+CxJKIqy
zPA1V0KiaW9rnI8Nh8zYSLWt4bpYuO4FRMKgYoVgqkOrL30mKanNjqDvsfFwc9ue1fNa3DT7Zgxa
jYt8S0TduTmp78IOGl/G0GzwJ5Dq/rDRUVIeHTZa3pSdlJ9voMdpGDI/aOc462K/zhylpDleH1n4
0Okp9PFLnMu8mCoEvpLE3BaYCLIaSWqEviG5klLojoqWwxu/AiSgy/nwge1UnxRzK4GdMc+1yQaI
2beI7ZVLBO+lDet+Op1nCHs+/RWpIbbz+Pu86GtrcAOR30d55lWruchEhj8zyJGugVGpEmkfEqaE
+sxqzNE3sRBiuQpaeppRdE/sUfR+JQGAaoNNNih2cI4gnd50jtIHXQIv0RMBC8eLtLsNTEN3gKfR
V4CP5jspU5B16+7hctxRSEtQE3upU+qKE0GFWgnI8jO42k3Ls/lCwVHwabXn0pD5HTvPfYyTAsO0
7SbssozmPfkuWlGMAnW93+UAHrkdAKRD1rDrA8ALxZ98CtGZDu3aLNla+OBFn02ih1F+LJMFQYko
dfbw/W00uLzRsHb5dNIkAdunppXilAcBRe+Zrh0uX4sGT6R+NAdyqvM26wixh0jNehDg1gcb7eWX
hkfUhusVZngnap/m7pc/B3p8gE2SeY1WMzVtfsCq3hZS3tXd09ESd4WkfK7MvdJyA+lfN8/q09ZE
kuJIkZ8mRVA/iWp77/lle6B4QR9X5yC1WBxuKCXEUUJj3xXA8n50Cbl5yk2PnZJr+KUx3K3Qm7w6
uIBafR0ZjV+LnKaENcyIMAOoUeVzeIYR7z+tB/7L4FHQ3wY2cQW08GA5ChCKeXR1YaEg+ORVsfqf
/Gk4Dqo9GOFzhuwKL9Y1YrbrgH0tiNRvPUqBereKYh4VkfbkC5RmgYB+vipgmkcA/se0J5hbLGVo
iQBlg1nCynJZuGkJ3kKMAKcfZ8ZbUipkq0TR9IxLyQf9oAkNtpkDBBtZDDplKF9Y+tdsFk0eBnGr
kXL8+ercFUMDzaSlexRbeOLckY72ZChPg6GdOcdNH/j9wbjLoFkyFBEUnRdqM58zrK427xV+dWL8
nFiTGUjQfpllhzWg2aKNePO/kcluFoZmO9qUs445WJzcVQaq72sasxaWfhkNqekEWYiqJfa1EmzX
fl7Rr5VSSdewrbSmxfE3deSA5OpyTDZY0yxPpjRyqNJl5y9raZRumrbeapnBWM6EeSoE+41AQmpo
BOVo0MdVxIAqCaOl9xgG6zXi1jxC0Wg3ciaoOBfKjPBxkI73DWyaJAXxIEnxls6Fu/Ir4DPKLeaW
NHoZZhFEWnZPJTq/59YGxjBX61YND4PQDnHO7HGoESDXl7nR3X7FUYx1/93Csym099K3i2biUFJe
kdB/wKpp+LMKpCPxRWTXvWDhcj78eQc35az4rslIyw5DdP3XnSBhFfNKULUHtEnGZDa5LrMr84kT
EqUmQuA6zq1Ym9mUEw5pn2O6CDT/Q4kGZlT2qbpBO45P0ONJPK4TOwgV4HtcFiqJKoeVNVucKECs
2EvMuGCNLfGOvX7hHk0zYQTMK4dL2mkvppmczio+aBqcIMXizKTKQA87PAqwNgCfP1p/3uJ28FB+
8Y53YpAtBkHv/iPQCMukK44ruqOD1IzLUhFM3soLRN3fgLHNsbnT6eLsrcl6N1r3leXkNpDYtERp
JSrmQsHOcN6mXQxjI6F6K4Q9fHPjtBNY+v1uOOsCM4Ww/7yQNrxmZF37Eo6ZtZHDEj2Kf2O/d/WP
PnTO1b4HX37N2Q7eCqSe3TZGSflh8GkeGqyYnLh4jaKoZ6jOk5BVhANDU5Z3aNfIq0ScnoVGU3ZX
YlnFRy795NHfZ2GRYKBrCrgujCpxO7dEGsuy0j/U0c87ZtBMW50LwbcPGFq1uL1bvuKjCHdXvbYp
JbqAirneXzwI+YDdMsmFMpdgybhCCU675nUNVyWLDVG8ghyqHoz4oIGwtMMpv5HZYeS0Kqi+lSBS
oQ5FYZqFOiT4wCtzuwDELS3NqH+ihwmrgknyDRjlQLNtjIAtpiKJhAhEapvUkqu9h6mptytjcZUR
Y7o5ZCP1LeQhojaP6ijSJP4iCL4bifRceTO08Apb1wdBRKl97E2w7AJU7QEX1nizPItM65DNXeeZ
edfUxiZzFbQtnMS/kOGgEgo3VWu1R/4OIrQ5JIceDbbqO1RoRT/OLtBpv1TeAcC6GK9fkE7VMM8c
5uoI574+kzvDUy4jczEaNkSX5kSq3645L/NJ61T/jpj7aeVIbT8gwg9HwW16s1CSlT81lbiVzvkK
nLAJ1aAnvh4VdGiJS9QFaewi+OJ27N3ZoxCR1SkyZ8F1Squ1ZV85Igza4+9IAvKHReKd56GGOdIO
cHKOV8RXC8hGPGVwAJk362TPmZ/49rsX91+dlfbdPpCbqn2/E1yF/Lm30wfgfYvkinLMLSbB1CLl
JFtj8l9wYqF2VNXNwbcePH0/gbiAk03+K8cWtO8M0HXy2WGSaJrI9yAV8wJocK5wj1EGi9z15Cyh
+awEeiaNnp9MPP7tVx1FSl/jFR1D1vqosjYdit+K8ngyd11tDdeZ3hL+oGDCmHYV0PXc1PWTziK6
fjS1YJNTJTc8mPzFkLkZq+zHXTSHOF9gVtFNg43gpOlzzymmEso2o0AEswTQouQ0pojCKC8mfHs1
C2ZTGJ7aHSqTJWPB/0azIsmy+pgv3oPhlva6sE2oO73bfvBazURS3ghE1Jt1s67Xfk7maHUvC8Ra
1JsJladSsyA5zvHhOuuQqMUH4mec6Hwp6To254Qrtl/C/NxW5eOygC8ruhyue51Wjdd5HKBRC0R7
6xuYkS3GXZ+kq1QH7PLTL0A6L/v3iPqVhmzqnL843uZbQpwvkTrH4aCMd8hddUi+uLvhlelpPsuZ
UVTmrk0oM2JVaQ6LgZLUIPW5r5MEMsfewzkjw2DnmGKcU2gYfUR/2Kf9jAzAVVm1CZ+ok+NA+GS3
2+1pZa0zAE8fD47SeMB0o2jsnWBQVj65n/yA0wjkRXlEnOgeACj7Cd0SqAlJGlIqn3ZZ3p61UEF3
7OANHmsfTT0sb+5kSYmb4h1V7pQHozvUQy9BxHqMqQgh4NOC2cnR2mYNR/WrNkiiWTdWbCgBow00
SgGkISDBFgvmfUA+OoFX5qP+yeBe3GjdorwOI2t76TtXVmtFOErUnHYpk2JWTmAA9bUf6s27dUYk
4LJgraL+P9DNpTU2Se+D6ATxb0YwMVaDhgwQ75h+MfrBZwYe8GQEbQ7yUdpjr2vIrANak8OzkbuR
VZmqvqAOGuW/pda63MMdHjK8ONj5vWzURP84jzoqnpJ/h+6KSWwWHKdJLaq5OIOfmF0DEftaJrbx
+2klVWcI9tMTW30SJVBxm0RteSvInBCaejfUBBjjvrmelkmBFeKhUuFKlkoJZr8jM/3HWUtSGvhN
XXBZuNBzcoHvO3ia3tqc039z9reGu9eFOcQWWZjnyIw8py8RYSvw+yxIKfYS3JTvrrBzz16ghi3Y
wYJRO2coUO1VXmITxrkQMEgHLfQ9qRnWRS4yoXAgEbSTfSYwlWmSwFfROCKZDQlO4GCYwSGaqX0v
O7hrGluLEhCvezeXzKqYJstRhMoMcCJAEeyQ8P0hAw0+ovEbFlXj1n2pY/eC91AII6w5+ZOvqj0w
9O9uM4SlQ0qtylm+CsPULMNK3qsIbDdjoxCMTcECoppK9pfNu9DdrVPk2ifu8X1apAV3YsMq/bds
ChWaPgTehAdCIQYtiAUJ+n2ApCNzD86xq4o6sEDEIdUCJjK5eiRPBJpHiiz5Nq3kAxzSLzcl7IxT
pu3iOmwMUnMPQbh2HnSvp0TJqWf20FOC+mlRdHYzDEamNN+FbdXyqlVJEVREz8t3PaJQG5pILWgu
tsdOJ7JCEKkfli2stnZjTUunh2ZnuExFG/yRFPhIEIAT3zBBQCeFwvCsaFeDAZNoW+fRw2QBWQcs
jAVGX2g0D7roLVLeW4j7x1+jQ+R31dVBUviEmCz4dZd8a9vjIdtXcZXj0kSKlPwN1edeHKf8Bz41
WKAnsAAnIWFPxjZajDWGUoDrhq6Hs8mp4dtYdciuMvnBYx6q4eTBloicLJ56+g52bxQ93d/+UkKy
RyXQaxXNBRC+Ocm5O1ep7XEqg/TjqvEvONgB310SjpPaBiLmDyjuOUS0iVXTAXMc9A+0kYwTGbZL
p34XtWyLU6ylhAkomdWKX5oaQys98Ux6ksGV4EGhPW+TwxfR5F0+huubGNaLlrfupDiVnyE6WUK8
r+Ud8kM7akJXvZF4x5wljvgAmnoY/qicE+i6nIEa6qrpxPE0T+9g4+xlFGzqVYRxKEnO75QwMguN
590RVDgjCmTJc4RXgpeVRcqo28bUzVW9K7KrLBA0ZXNMvH0Ftu20Qi9AQSl1Wvfp1UBguWsyWG2X
5PsS07nYg6s5A+M6vmmJZ97xuYOhwuxbKX+zB+oRwVa0S7fGmzwgDdRIArgTMsi/ZywaZuITbeMD
75LdamTjoamIrdL8jcnhptaqj0PQwZ4kQM2rdMI8XSTa4nCX/8JXTZ5JCsmd0wVHoUOh1CDcApep
9Q0tRF/NEjrGxdEtR+4Vfbyb/RxjqB9msPWE+T9/XH+HaOJIAEEa0S/e4t1IJkxLzGeI0IJub/4N
k6AO5PKPQVcBxg5mcoygwzc5bGvfS0Op8h+zdRHn4is4FNu9uYmoieQJYGEeHhB5Lewuzk2oHv86
HhrnRQfB0LvRDFppk2mUkgQ256/p64p0f0SiCmXcfS1vpY8RZ1o293sPjFK36VSwHi0PX9bjW93d
ugpALRDP9fZb92KQYoCO9vFaRoKZvsQnzVlbtE4CJbXw4t9uArA/yP0FKYTMMEtvCeirGWuzDGfd
X1vj5tT8YWZ4lslTAEby/XRFpL4PIn9mGfIcs2AV6T3HDy/h9F0Up1+tCSG5DPbA9O4kmy+M7vK+
bpX5HksvJ2YmQmDmesShbSKQLaxpw3m9JxCEcWMlQ5xn5vHWrDhAilEE47KK3iOMl51BQG+WAeJo
30b8NtLZi8+vBAdRrGh17vR9awYKZJEVgyGT/z/445zY+2l2zFUjq4JSOzSIP+SPJkJ3XP2Ekb/b
cE6TQTXv90AbFaEHbiVYTRpuB2Wrr8Un06kEfi0FPGDGZM8KKaQbRSskzfD/iwsogdQ8igVjSfQg
h6p8L+FDTLGjllzj3bG4VoNYCW8svxcjgzxH6Ndot12C2Xyx/FgjNvCEXzDIoClHuitNhdnCIq7U
tAutMMrBk5ZAizzvJ0Ry405bmLuz74srOpPi8fw6cwIwe6MHx9/2ZrBxWj5ZQskNLx6dVIGZnnu/
kc8UOy0uavdC+s9X8gmwrsRf2rpYniR6s0spa0Jqxc2/Q/JY3j5+ptRSImIKH81/AO1dvLKT2MNu
RIdNMZBYYS6dIPi8kyxdhDXuPedfA/Mq34bhfK8rfDaS/KAriqONtrUWRWUFKFrgoGkMtcRsvK0C
IWlpE0kx2Sb0esFtuWd5NYtBxtXDJfGXrQZ+KdgQo2g+0phHzkpyeZiW4tyLErj5SoA3SwnzgTmB
PSvonQZ28KSDTBeRFp4HleDhm72vLYEwe37KyG7q4soOyjfPlW031bMSZNQSch3cS+nN8tbZ5J/y
4cssRkzmOAk4gKQtUCXtb66F02n2Sw5paIMHOBmmPnAgzR6xQxRz8YvqhLM8IPTyroIYoIC0Vjk9
7N2nefo6oFqIEKAM+kJYZvk1kma74mLfJun0PQNhMMk4uNTdyRVl7RXyvd6AFghZk52vkI2INT9B
bWDVhxz8SmQLh00avgQs1/oEXKliZrLdpSCLIg5KC9sPYCHOswiYS+f2fS7CdZYddYZRfF3xAL9f
5CWiKtQRux1H1qROF2jvV3QI5KAGwGi84QEX7r34x43jSDVdoJESFxGerObGAX2xPU6ud78UCjtu
Yc5/ZZsO2V+mCxxBsc3EgbUr3rSWzplqEhI9pl8ArI743jpfgP0AjCC+fd2dfbOcyh+9kGYmRp96
yFt6zBjW5X09I52UQM51nF2Dj++WlSRJw3rdQNoEGv/pgafhKM3IZhJskfN9ShIk9FrDc5fnbexE
eiHpdlE/vxh6nmFPuyAIj/pcig5yKuKjrvUoxKy938zw4/lDDs0BnT1B4vH32oa2Jf7LAHe262Vd
iBWltUf3P8KwV66LeoobLMYQw7L3UMh4rTIgGcJKCPBCqWJbP3vSTsw8A/VgZ7KaDwlcCEMQ2Nvf
YrBnyxLpsn2eApiYGyPU+Af4Abq4yYZ2nXbfrjjwzI8J9mkOv7DLKJBkPspfBKKPfkONGq9Xtgrf
hHwq5DSV374pSspcGTAjalDCTDdHdEmqyV65c9rTpO7qDNvniCT2DRCbOhiFerCQsgs/MCSBATEX
/syL//+bylDFhqjLZONUchUGe4fJCub0+GmBKiAydgKMHmu3Na09oK90eXoVvwHWSPJA0DH+1s4L
erDV5FiohcWhp0JTjzvTrKkMUpDaoBVK/niHgK0FxZZVn+Jer0nvgVoIwi8LfD2LhM9ajbUqLltw
H2fmgbi8UBE3md5/O0OUCwxrlxelqYS//WvkdPALw6W/KQ0+W8SQZuDgkyRNYbSmOuD3UR3/63tg
Hj3BgXaik94jeNx5OM8EMISr1PMD5iz7C+WIHUc7KipOXVs6LojwN9LMJS6RED2OEWIJmorxwjhf
DMOs8Ff1RFWHdpTMrrs6Q7w9gGdnsF6xHyaDrtEh775gAlFR66sZe5PMBhk7yJb7UtsiV7wzCwhT
z0xXJUGaU22lY3RDeN5fPGmEscbVhbLXc1za2pOhHVElkdsSu/E7lTps7j8F/7VSQ21MUqJJQjE4
JlFbAIVFOkNQTxe1BUb+svEh6ZXeGeW4/oxmLyV/RUC5UUiMAwVMkEKsBanwA7SeyAPNXkONGBVj
EpO6lvGEBVQCheo85LQ/p69rIKmhfyWt7WfvUg/BvULa8DWqE25Z7g4JJjX8xw7PDE7Znrz7IooB
0G/5jEBTyH49IZeW9x9Pw9iVJ8sH+vTrC9q/+dd+dYwC0whaawTYyesQD1S94K/MJpLCp11crIge
y0k6dMgibNxorI10XHxWLGKkkXSqcWE7SjdNUbFDD2+J3ewJHFV/VA4n5EYuOv6jX6ou5wAHzs1s
Rq92+LsLt1kq3ZZ3eoogtbULf9h7bCmAMR+U3RZcz2Vd4+9iRUDfzNqoKEtxdKYc5jZRzgJsE3pu
qMEPuB5tVdxOEFnAVZPvFDxarymaa5+TjGo1rdxTYD1RL4HmGYasJDzco+i2W5ncXEvRpDbujuym
QsKBQwcpaQfDS94Q2lvCGvho/tJFKFplfcV4KXNyf3GOTK02HVfWOypTnJPEawXJrEMdqyWZE83f
9DbuJrAMmlHnmA+j3U6IOyh+MYpTHF23ntzHzfZJBDYjBcWirw1Ew2EE3aIQLxXwhsC7P6WKGRNc
uL2HQ+HgtdQ9RGOfBZHCEeHaKHLZ32JQnFys4As859fmjUGEjdACDygf7Ux2UJWj2n9mxd3so+/V
dePifUIVr6HZ711lHTunhv/Yzl7Uw9wjqIQ9i4hSOLi0XD8kSdGIzEbnmbu8lTXf9iCUCIk6+cM9
hSSXbeTSmolFsqUGblKd0FvZkdUuTjodejK3sLB5JPShqm/sNO9onYHoi6I+K7JAc5PCHO3rqcfx
yU+qQjCmaO7NHIsDAok/QIJ5czsxsNJmR3NFbY1kPFwITyo/SLUcq/jHqgF9N3j1GL74WYoCvT2L
qeCVLHY6so/oFuWp99PUIKSXe3NanGGQvNO5/eQ+fYqZi/8gDQK/iz1WePm45TYA+3JutGulIZ94
rYvfj1nms5ECP0d0MucYetBtfRV4bDunF5eUbwtzEPZkWm4RJvyf9tzXwytwVVVLjwp0maCnTe8u
IoHE8It3CqqXhXn+uqQhEc9UvcBtGCbfjsWv5mXY/80ezAXDRXza3Z2yMlJqI9M+E+wVwO0kvQ51
c+nSl9z2YHnVXucrP1s2ey11w9v3PqU92d6SnRMFuyS+r6mWzhOthmBZOdb8j0BaNplPiI2JL82x
UE2VoHn43w7hYglQJsIE2bsALlDm7DZID4abHXVOyvh7+gC66qAFq/3s+4U8ZcumBUFCtPMI0aCO
SUrqvf0EjecGM8ftLsTKjwk83KqOy0qaO4nmRCJgmvOAskyV1Aad+Wb/ZEA/88xcrjnPSnmQDCqf
1kDndJULSEYZaMxMLlS+ZY9OflVOnjJsnhVyTYOkU5ssrxW778y5bjQkBWvyFeMaDwVBRUNJnWmn
rJKlLClwV2qYjQ0lCPvacP0POGgZaU89rZFDgqlmvg74hXhjVHEqXmIhpO9WjbQXvpaXhU6LYqSU
RM34T7aY+VwFotk9hAbvan50AYtyradXPeSQIKtoIHFG6HMaQqPlNTAxvEggxeNc+1aDFxKDn8ZP
qA4WhkFtlRaosZMcPN12GH8TBiVeqSq/H4g8M6mXWjrCCLGLKQCk8Bb5s9pGVfdiLM2u/gTloKhS
fvdkR5PKz8GE3vhuOBeomHt9aap//b0RgXcd5nQPF8C4HCaD0RPL7qB0lPofnJ+TRSR53mTzivJu
gK4SqXt3206Mv2lsrIvB7QQuwQxbus/W+gZkggOrwjbJg/ptbIpAYz3eqvl/3fJNCo+FYxBrAcgz
66kLGBWdFBI+FbvMZCGpYpLP9FmEyflHYWhTnvba+oxXMYUe6VKQ+7qY57x8HPEusYxF4K7h7rXG
5jrW4i/XEEGQb1y7UzEBLAjDCe1GzzKtlyqxi/SzVmE7DkZR/Tb/Jh0g48JXlD0qrawTA4d5WN62
S9Hd5SY12KO/Y+mQqT7nmOVLfkJ/waEtg7kGlS323oO9XySIKr0yPDSwXyoDe1kqYrBdP30Ro4GT
u0GOW3iHuZ90BffbsMwbS6QdTrLXp4R3ZU0e5zQURqzSyWtyVTyY4GC71ucOKksIeokTbsBHOb77
Eh8BWMgPIZ83qCkhn0I5xU5jVqjpWDCtm2XEFto47Ed1qlOIuDTGVs9zXy9cp204r0S5poaiar6o
F7kBoY1BX1K6ECmZm9CJmfGJmAOm56EVp610qkJB377DjAsxaEEpBFAorKF7nZ1YbbomaYcSJniV
lyYlhcaBsoWZHDtRvU7BOcTijCqvKTDaMgJhQl7Zeg8C2Kb4qnxe2/NjRezAQCeiLYvFHUwBs0Ib
sQlgyGUJUqQ+Lq1zOMz5fKqDD+k/1mbzZvKjeMELfUVArqnCtPRZVJO5+u3JuG/wq/DfIlWdJgSl
FKGfhRvNXyEwZKA2JSgrd4PUteO3BJ4rSO1smd1DXzMzglFjFRjVlXiYj9kHAUokcL4mFUDD1DJO
LV1KvqnrovamC2fUsvk0NnA7E8zV4BZ7R3xJlLKO4AUOX3LMyPIYU57+DXOq5P57AYsyy6IjzN1O
wOcycnx+ZEBz25iq/h+ql3dJEBtxjUp8e24TkYxBpv1ZTMtx+SyOcb+SkZVwa7752pOK0/6vt5CJ
onNdS5444UatBsedurEC9eLZhfLZUAUVyUicR8YU65Obb+J4E2UlVtIOT9yhZVR0y2Ue8XeDurOr
uLoB1LrQDrOmUuGNyjw0OWm9Vh16SHizjxojxJX4QjzCsT/NP4MTGX7G2zNntMi92f7EUWBK4sVT
A1xWK9fwnpdAzD4km0Wix+SU66ZhfCb2dZtLCVC2Kksh7xdTPBn3z0FpWiuD0uq6r8Y9ECIIEKNA
dXOxvAoKte3k9q9eNC6lGTojLvlyCiaE14xVpGcCAo/N+HT8PffI+8M1PuIgmj4K7kw+6AZ1eukC
K+DKnw828uubGa8kUYpaM6/EM3SRB0jD4LF0Ce5oGDJbMfGzO89hyfVQPi39DePEHyuWyUa8ZpUj
wYdt1SRpOzVdrwn/Ihjz0Bb603O5wpClwIGESKNr3VpZRV89/h47jR6fmmpLeu7feh6nT0GwbDp8
QvDgU0MVSEYuhTQkLYHssxTvGO3Rq7AwGBcJu/d1uOZT+2qNrZV/EBLdpSORCA3GAPMuOWKnJfH5
X20RJACiCVcL6DCtjZ8p/CIsz28cofAtZ0iRZQxQ7wVabm69HPwnvgthxl6KdkEc+SrA+psYAEMo
4Emk1brXc9MkKrVujXpkZl1z7tEKhWHFpEyKqKZ9zwMSvFtdFsT4cWhG1FV62uBrBo68oPQ8pho+
tZUWjbxQbddaq5/5yavtTBIRO1h0B+9frf6e2eQGedrAbhTI7ew2v9h+0piOzwT+KIoO1aNZO7in
RUrmgcFG3Pm95TLfLmStRZmgDWSLxgAaxTLlTO4W38AH6s7OsHS2S7ylJr7fgVrbOGSTK2ih0e69
6MBMmhZp/OMoVAULWzkHeUnDoMntBirIvFSSmBNesN6VmU4wn/cm/A94gfc/Wc4YpO5NZubw5jrh
5eTNziU9+YJzXo+kyq6WuD0sQDMs04AsWzp6xRHeCpEJcfpSusBS62nG1O1GXciWHrP7Vab7A1te
mtsfeHwMzPJZ4ADm9zxc3u/K+0lAZAr6w7lyGrzgK4RLG0pP5jXngdyxudL3/PtJjiCuainn75fa
czSmdWKqccqvy30qLkLHI6riO11hYey+68anKGfeqc3sA1hoSuKYwrUHPHeCifdqaE62PB+nxmE4
mNhynfiL3BoC7O6WclyT4Bazs9NM0fAzqZj0Ny0te4q4aazPPJUozxsSorpc5shIGuThP8Cjk/bg
+N3mkvovun2LNVtFlrNDFHaTAykoBaiTE8BN4iMNdjHSxlILMo6CRb/6KQi7kv9LbaLnc5jfqjf0
7BjkbWqjn0/1x7thPwNU4ApePD7G413gT3brU8I/ZgVALjK5UsGOBojbAJWmDar1zl2rCMKolQDq
9CcPxpYlhenaRPpAPLh1jT7J159LgL4L3cHHRniqJaFxiTvZFYdSPurmlGmKkp6DsveWTsRuXU9W
sDf1BF1nPnDf9rj/E3Rb7dY7GmXlIUoFD9lkk8uhwilWugezTkQcAAfy/4mG1KgrolEovnCCvRjJ
fmqYhSaLkDDyD5FHqV4Me5dg3GgTIBpqYmXNIwIwUdU01NxY4fPn6NqWjYtK+Xaej9k+sd/kEjWh
kFMKaQlEhBIS8cimbOY9Q3c2dMZbdKbaekzeCMWACNlSVJnA8SvSJq3b1DZzKJbLWndcprYqoyl9
AqEBeLKJY2bXWet4Mp9pXGOs9L4YNBqt/gAtV4juV90WxPiG7+CBeDuQXgy2RVSUK2GUdFVQe2LB
QDhP6ofzeORFh1x8BQRqmdk8VMWZ/c4+u5yNVW74MRPWcK6oF/qi/bvbWCQ1MPDqWijfM0UC0Ky2
B/my7lxbJHFowyWwjxcz4OKVN4FaPsqaOb68bSq/VJ2z+Z/GXLXTKwY5TkJ2nB1rCTsbUiTixVl7
YBKWO1qTUJ83JPAu3tnIDzLULfV/+OQKpXHH8oqvAS4sCngyOOysWkkBhHXOxD8Hq/TOrqWB4Sbe
0rg39Q8X2rQ2Kmq5NRG0PC2vN56Ao6v51KPK/lI+NnGdqKtR9F2XVY6yMR8qCABjTbDwas76lZMB
qscHH+IXaHn1V1eW2/L2wquEohBIxZUIckwRG/dLRVWGU/MulscXKjnixt/LEmaIbMx3UXmrxPfT
agf6UvlKptO30PcqiOfoDrtNnA6cCgTMpivqBXxg85CPVCYshaAWLD3Hqzg/VdYrWpdOTb/uRJlA
iaIzrmAgqF1+ggs1YRPgzY4BYgrRfevd2oeoildONyO8RE6HAYK+A2RH5QKYrt91qr2D9qifkw6n
CUhTtXZq/hcHUUmywkMat4kJyPVFEVgsYiOgkbN6AwIvB1smvu08kMGCjGKKeTyBnj9AmpYXIfcn
YqSNrT7D6u7KzvjIuVU0fFOpEpushUttsymtnIl/ncCWA2k+6TNA6JLlIo6CsGKhDvoki3xYJQiv
mgvqE/9F1aQhx41QP21nm24FzxJZA7YStrJwai2oppmsk9OOnNhGT/XJISjfuXbR85IlzhQz2PoF
4sqB/il2zYmsGaPTjaAnN/Rg5M157uOGCV43yEDxlWi8WNGiErE63vtG8S8RijbfjBpp40XCTbPJ
dUfvPfKOa4bheeo9HJsgG4eie65xBCeYeTuNf9qS5e12IvpPjaf7uq0EKNSjpRUbt/puPMNUGPRr
VtY9CLKol30S7zK9iF16f2gr0iZwTml+fKLWOghLRYusBsVb9e1g6A9dKQXTQZc+/1sCxixGWyn5
XEsFRzArXD5WcV/ho96jNyy9Z/MeuUn10Au9vwBY7NMl3gd8c7WwAQMEJOQMeFFJSlLPYd5cJGsA
oA2R7XcA2bhM7VIOQSi+YyT9YNvMNX95t/6vzewFIyV8+XXLcY/OZeKpWAtZUxtU1IspiCWYvlA/
j8HMQtaPP86vrobO6yfSXws3AbexWwy776cr20s15pXXvxw+Wqo2RevtaEFFTWKMWrS/irsKc63m
bozAieIOchy6IebUGgbiqnI1I8miZj5+MRdaD2DunSgxrqf+XzANDvmeFF82F1ioJToZKfTQIEh3
oB/TcobUBsxv7V8xnYBJRvtZLaMN3H5jWCNayaEBNGoO98Ta4QAVLkaW1zYw0lPw1dYFe0js7s87
i8Trs4itwVsDQ4QtrWlFTVW9Gvd4zMNbrbZIX2XQE+u4USu4gE1k71+Kz20GMm5dZikw+Bv7LyPH
9PW7E/MSebofTUxWVK+MiWA7xVRX6/5+Y4htJLr3L8DPmu/02DdNjJoe5rki7EopBBSxadumiEVG
Xc+laJCazl/Cf8lbrj9nB/p05YCblczl+PwfvwxwJ6korQGQvlRaHzLKyhAZm7PUrKPiW7W99+Zv
vV6NiPIacbPv4HWjxzG3szzXdUUUo4X3QMk1LlR9WWd/fMwetWtP8hcLLGzNC5bFPWr6ak2d2lu1
DlsS4mcwPJRu6e5Cx5OgHpx48dAmeSwPvq5iq7Jamn/92gxONYSZmsBJiYWe/zfJIkZBY5TPtTHe
tC3KDFWwP0Zx5TebeRG7raXlt1uzfI2TjhW8tlTiNOYEhFNDXDveHc+N0+rk6kwD+J3ArflYW2l5
+QqpjzHAV0nvOPl42y0QAwe9na9GW8ZkWK80AJq83I4X6uAqWgsGchItrUkgK74H2sYauq6bHsRy
yDrfsg5Eh8NdZdObE8gA1+CwhN38cZGnYh/xN+3pXJ5yK84Ra4yQ2HFrETVusMi+lqcl5RK6AfuJ
G4TeB1ng3lJKFRoYsjPmDa0LyLE5BVwoNzXfKabBx9bd8+37TIdIcEyMHtK05+mr7c0zuiEzUzzi
JHPZsCcrlk1Z1CQ6la4VQVZteKXuiiUgwPld/E9IloRT9BqU0UqxI4Beyna8jhxLeqO6tKg9fUNC
u3BIAYM6ZNdvJ3xZfkBD4mS8kQT0BazBtglzJSWEfPJGSlhZTcUikIrcTlRGm4j5uIMXMK4FvFRl
Dq+RXqpQVO9XLjicRxcBAgARswxfXCXG4/XpvCXHyGBaxJb+lRwM3lggKwwkp1lMPKijEOQCxPLc
KkAA2mr+pJs5aoKvvWMF604P3zjn3YJJYnvcTWopXeq1+MvCy2TKnLsxQiL33tP67WqNcWheRxe8
GXDP7yfPU1oaa1gf+wtjlchKCZ6G6Bbi9RGqsTSVaHwCIZOmW8VFDOdjevzIRBoHSPWFPZFyZ6HQ
7qwJ+Q36BAX00qUvGJHSK8W0X4wUpL4oMH+M+jKv+IrWQB2UQfMMLGa6z59jHoVPSXuf47ITjkJq
N7eB25+y1QAwPKX99Z9W3829L68l6wy/+BBvJI2sme4sJMXWxRlonMXxbuKE0jfRg3N7ltMyTqhC
2G4R8DS+bZQNQ3wBB/OUYXy47yRfP1t5ejULRaOX/Y+O9lcPhCnGWgwefUbDTyGMe877GLIFISQ4
NUE94Q3uw3CxShWmIdR5kGQ/r9SPffD3RpAqpK9Czqky6hbVWMJV4ybLp9h7LdfUO+QmEZswPxSK
CIA3LE9RvyoRhlRDVHENFlW0lUTkmF7tnk2zFWiCfqUJkagWwXJhDcAiEOX2psOHNT57iIov94kY
VaC9AylX4ZQNXYUxcZDW0meD06UI7qjHdT7Y4hAUcSmxyxQlgjzgA1X232K/J6ceXuq/kAh2woIm
JUZge1UhfR1UAtwyuiMNs0hJYoPCwmSPLB6iVjAKKWkalzmrtLVZvK5OermNu36A7pfz/WMup0Aj
cIHcXjSogDjloPdC+AAU7MCP6VWK+CYgomdu8FAgkYh4txhxJCcxmPAdoAfPLCofbARGRoBYJsJD
1l4FNpnFYyLR1NL4oYOsfaXZjNHb3HVeg40zvyOXWjdt6lIALY+DOU5qGqbEOGYUhSQGlqugugH1
Fx/DiB6nHz4ve1FUmil4S+Y2Uke5hkxpJGo75sfN+fd25IyCE4sFLUnUYbU6c+2nfogT4boHiCAg
OLo8V+2TnVzawUExa+rHNrTWXOhv4ceDda9eMd9rgqvBAUnPWaTzdjt3j3cJoy9UzTJ8cvRyQ2Qf
q0BLNpvyTeSnay8UMjecEqSXHrg3qFJlm2fNZy1k3ggfoqrdDNAZZJ5oOFPNX/qPdJK2iRcClX6Q
O01muTL8TcGECtviEUsHqH/RM9Nx8q54PSjZzTynQXB1eOrIahuKgbo52bRjL91noPZwMt9E0RCz
ZdAIxGbF/BMGfLxeu2R0sQqZ7HGHU8+LPr7S/iSNeHhdOGBN0v/nOIaF26oB6Ve5CgsO5m6QUWdO
+impfF9jId3xRPnSHO9fetRebnojJiupiAjGJ0eYPqPyHpO59sRod4Z7RqOmypb3iZ8x8WfRY4/e
91+hhF6/+cGnAZm2aqh/UoPnLZH2uWIRW3jISPx4cLiesZTdGPRQmNLjp6343kcpu+qUafz6X/6n
CXkB+Eq3cIwYK9ZJhCIPKg01eu48miR4UWkp71yFm/IdzGyJ/3R8hhI1wJs+us/DbPowAgB9eCVZ
oqZXNBih0yCuCnI5zf8Z5VN4BW4xRe4X5I1KnFYyd5AkyMGjkd5axHYvZAyeJm1Rj8IKq++GUMuj
BX3G5HN87H+OYx8LjgL+KJDPr+MGjlr9Gen9277BNtNzdsFtGy+yqQ8Gm96Fj5FlVMurXpKApRhD
itgVcB8bJa4E+XzSkZbJ76Th0cj2Mld7/xIdtDpDPAzIIHVNU1SfgF9cJTAHJpTHh8q/D0zvt42U
+BtM0NQjfmyMvI18XERPuwTv89VSnEXH1eWbqdbzJcez+a/XefGGpLq3nouOoIcPIEkpu3oEogOi
O4q8VdFKmesM4NJvHbdrOdbP61eqFHawNnvucVexpQc0uZp4qbH8aikSZXsqUnV/APwiNSjB5exy
aDhyI/bmUjfvJgKp/X4sJYjwZ3DCMgKKtPVAJnuPjayRg4dU32uE/eNfdP+TqwAGlB/JVhv1ZIVn
+rnWT2QvcN0hRGQAEtQR8D/Epum3IKaX7h6mpvAb8a1xSs5gwN/k/clNgNsXeAS/sYX1cB//BLAU
qgwvs0Bz8xVPIhmtJ2HVCKJguPRJMxbRaNSctqtw7ryvaNM9+r90or4LY2Tle4ynt498qJpYgAAq
ALjMVZeWr6SQ0DCYU28ynbZzZat2fxZHjHMf0CuZjTqUF6I2j/RTyW5UClAdqpgC/w7EAFGaZvSL
uxSaGkwWkShEGqWUX5H1numYM3aL1HnC3WCFIsopqHQ3pX2xPp/HrF4A9zM7UMOx+uZ9WRaX6lfL
5iMhpxMM3GbvIwANrN4QaZmv2hpwk7UcwckqRoZLwPzONukx7ZEP+kNNRQJbMUdVqOUuoZEdoUeL
j72OqDumI5csdjgGFm5hhtqvhzOrI8mn6C7YW91bVP3nz+am3/AIsFMPtBo9Gm8MPPpVGb+pm6Y+
5I2NZpV/n1fY062f9lGL4EfDJ1jTu4w2OmjVJ/3t3DcRGrt8qhtZH4gl+crvILQTHhPB3rxFAFjq
t120vwzQjVHxk+Emlll5yIUWoCi2GKb5qDKmkCs4jjXOLTkniq+DvXAfFl9hAMNvzGJERkGoM3ZJ
2DpuJxGQ9hDaVHZrGz05gYl/botV+5TtCw6DNceHYpejZoMVGrqjKatHMhbrojhJ8RNPoTqm+E8X
xiwj2cLMm3FNSIBSC7syKMWUlO1Vu8smdVdmb+hag1iNv2T+d5uU7M2v/zbechfZ0+HgQVcMxEjI
TXLWtMxlvY/1/4gbeIeFZbxUZz+G/ktVIcWDmsp8lLNjN//z6wZNs324Aw4xU7ZRZK2o0DZmNoEC
IOYo6mKk11IM6FJZEa8wfCpqB7TDz2wlfEClc/Bi+8Zdm7nEvfa2XuxBWZUo3J0fEggBgyfi4kry
Y+W98k1PQ+UgAYtEgM7fOMKuieUdfOy5G1PfcurKU0gvT64SFXzRDxP9DmP1pgQasyp7xELSqe80
Rdd1C4JSpDDvrvwm9ja/OrDQIPk8A22BSkhb7nzdQgyhbsXKmrM7Q0PTMmOmiwVAD32E7LJUD2Te
bikAxC4CGyw8s0Mtg/00on/+jPjKI+DjkWN2A5MdHzo6J/hU9kirR8upxIGJRBZJwoOH1ut++cGq
g8VOugtrubX1bLne6jeZx23qFahL3nmOr9ot4zv7jwDBuHOXB5jk439kcJeSuLpDwjj6PfgK2MZP
u2p1S/E8SZ/MYricahSSlej80Zscllra8D9pNY8vOeFbsT08vwwKE7Xd4+uem40UE3kRga1zpq1b
q8vvF0MxJcjOrlvxGruLWhXFwPv1TWgXq6fQmJFC49uwIwJo89CTlqNSBb9yyncbxW6B2TBaflfx
kx0URSWKiUIMzm/qc/Ru3s7cJz4VCiG5fE57mXiQrSwyOfWo+LD/lM8S+qTQBCui2DeD+eGeAriO
KIx5FzkBYgCIfB1VXTuBpqCCAxs76IZf8YI+lwkHJs5UKMesR7rb5JvlsEDczSmKcL4BNcbyAUR9
uODLbQQKXh6BtbVyjQ034RcTHlrI6iTP9SVWvLQE4KrJiFOoWShlJ0WAp+hC/BTaN+wtFlM16v2+
fqzuEXNLoABJaobJkF6RJgeLuu4Z1ZYD3NY3yJBtgtdVMynOqVIzQjIY4YScMfddybwXbjN/opCq
TAkgU0MyAC5sy2bsgwtuIHnduPLyPvE7ajgsGLbmYrImOibQs/CtIoib1iqJT+hD3jNj2QC74UGr
9ApsgJ2N6WdazotlXEIV0k7zRqWFcakNeu4Ac0m1mwSjQ+SJg56og3d93FZ3e7+XLvgOscp47Rvv
uf8zpGFRPrFDoyLuCAdb6nlKcD1XBpEiAZ3WnGbKx9Dej/KsXEDan7PDRnKecjdVSBtPd+gFwFiB
MVlc/pxNz/YBaKK2j7kf1ZXvHSTl1qO/JOLVhF4kfRxonJBs1IYQ+5U8MWPr4inFh2WfqbfRcL53
T1hR3NBMLqK1cFORNUbAzUh+itVu2OWrXmPzgsvBNflpwbdQtMnbHfncC/lU7psqzMYbiyLJbG1t
8MmD00I7sQOec2hiXQ38gZP4VzxkIkSsgFikrfcd6+/EDxiuHVpxdk7KlhCn+VP96CHuPmW/y26r
UHHFI/jrWa2+JO9BrXL3BohXgrxwsziYTWPix9Vh91lbZpRRwcdhNPtxvEsXo9+bvH5qM0FQY75f
767LVCp10rRaG7AAQRyhzpsAFuEPhPMEYVah6zErM3vrOfjVahZ0Z/23Q4dQzHb3muJEsA+wpPAE
f82O4XiANR37SFjmuX15kEzRxfX/WRHkvUeDyWUAEMmYv05NS1paz9QggrYd0+KntU0ZTuTOT56L
OHU9vvh2nXG57v61y5i/Cl6L0wxlu2YvMFMrz/d2IU5N6rBm9s4hUBBC1P8CpbWsc50EyeUSWJDE
tnsSN272lBiGYtrxl/LLMOHqZWLJVtZZMfrBbPWB/YsMS/LUURK2BwY51+6NCkMWdqsjoFGNdVQ+
ML7HkrTe+UVCJoIM4d+dUfyiUlMUY2BmUGetCqr5VjlrhxcyRWqUQFNxMRDL49aT/KUpIzE7pwjV
dYhSNCGcwBz3C6eGe0ASD8kTsdVwIcOdLfMXls4S6itD72wbO8YyXHZftdCALk7TiMO0vS3eeNxE
SwJaBRSlu4VUpMhp0LRhwp/vdUp3HpqDHO31prRD+AE0Bm50ZIW4tpT2959KADN2rsu0ywY4Pd5m
0RxYJlSf88DlAniXVDfr+K0VCkMJlAhasSdUI0WzJU9unP0UuxcrPkzQH2//0viEGH6oFdDZsYkt
sNkNmekp/Qc2hY4CykdAI+ct0pyY2GmsRxCvAoS0n1y4Vm8/052k15fEJyjudmZQhq0Gma9rRhlv
ALeJPJLAyjpoJ+t4nLJyPwVyaAngwZ2/5YSnBw7NLccbRH9iT1uvODbYYW6RrTEsPEeoK2T4niWL
RkS6EAZ5q0ZyAOQ6af1k8W4Z5D8XSyy2ivqnFX1zuC4FjU6uoKsLHL9UGOCuvsW9//9Qt+h+ncnd
XLGI+w9LDb4PVqHm/nDIU7MKUYDi2LKTjDo+8WbX8KMy/iZp3MvucGst03lHGYZj90ys557iS1FD
OS69VsU0uh9klRHXip7Ro++OTcpnqdCq6ICYoZuQrTTjGBOfaI1c4Bf5aqV/m9dFlw/kKjWp7XqY
MuYD0g8zWDkC0IIyHvtrZ30tZDq30ayIwkITvi9PLTa3dKccY5YH9nTUPpxWnohCWsh1KKx10oNS
ykZ1B9r66YxFAVhApUg2r7IfrevqEmNYTD3HFFhAf6sy6NR3NpX8YjTRtlVkCMZ/e3837lRRJPut
g15xdulwo2rWajDABkNh+k9Fw11DVpIoEDaJxj9Ho5I0u4zsDj7HZ5kHVlrW/zBLK0Eo4y83gbfi
PDdVrFjTHNKfQR44uinlmjLXU/KYM3gx6h+H0A/NtSXRyy5+jseqwb9fBgp4j97gWBvBpmz5lOaO
tJ7z35bRXAPHCc++XZclM1f2mlBl5SYN0oZGQQAMldfCa49U3OI+N+CjMxJCW6Dx/I0eNBOlSdWT
kjEgbm9Om/wl8iK1OPz2WXIQFCwTfJMEJd4HHVy+iZrg3wn2T7s8xEoeyDcsGuyA2PbXVEYszU3z
BJSbRliutFIiTt6YVxr/hhoAD9FQm41yJ3t08L1HMZ7Iv6KSFz+mrn3NiY5EAafDN9KP/4ZLdfYl
yzNxnxVfGfAMUn+zdRUj2Sv2hVk9KPE4/Yaf0vZNufCnlzlLgaidGJTgoORIa1f5H2rkJ0M5usOd
v3WntxuU9xs31TOAYuqv5149Uxf+cCjA9Qvy/lyaTzSWsyvyQizbwM82IIZXh55SkSz4j6BwS6uC
Q9KdRkiMOuADrcEEBkK6DgwBLH5lhvq3k5MleZklYV0hVcgWDm7as+oOSX3H7a8QGp1B9hXHeIIo
U4xLR4A92I/oZhxZ1nPqxm3xApMsZGuZ4Ai3glWqGOuRYvJ3Xmq3lyM2TQBhoacNbCOVnw2vjPpk
Ai7XpXQMaH9S/S248jR5V0+2Q6poFAdoQGFJhcRHI5mWTjEjMAoNc5sFLQrOjQ8TyjytgUQ9r/lT
ayjI8ZBg8v8WZcQlLw0v7J+WlyVU+rtcHcji0s9sKGawjV+LM3Z1TLm9oHZcg//erpR5AbIGq/3x
mTy/NPpnENbAKHV4lFD60GTwM57rPM1fpi/EF9zS3L/aW38/KaNKaV5Hl9Zgdiz1clpLz/HaW8GZ
3q9fqJbjdq+9zEuzUP09uStC6wU0Zht1oBRcDnNcx29bcBabx2hQxh0aUcfyqymdcWIIsRfh6YJT
t+FObYO+kxZMgHiUIFbcOA+m3xknrJwfyohxEa2EKuUTvSbiKqfLP2d/5DaLKh1vWSBWFEozl4v1
TEYKN6S5rifEGDilMaCiqKSd4PRe7TLZS/aSjGoK2EOFcqTHp/qbCDyFpx3r1qOaPlzO5mcqbJOQ
WC7w7/JX93kifR91Yzjr4b+6m04+VNJBdEjywVXNmFR9l3at67GteaVsUgRe/ZT4NgAowujcWxQY
diAh2agYIrxPLFSU4SgiGGiKao73M/BxVn22NXw2FDKTOnpOR8yjzo/nn0kqmTC8tioMB1TzPNVa
vLLMAT6nCEpP0Z/GLsb6S1+SldfjQzizC78/Pqiz3aGi8ORIqEpidc/vLNGy7BhTwrvhWovZyFX9
0eHDlJ+UqL/TRnhX9Wm06EBdpWons9iXiztLL+ya1W/NcO1SMiFKKAqxExY7GHzgJTBOOipFolAT
spA/uNrJWfgkSmHKernb+bMPOG2RrBemgyqL3vcbn9c7zksq21mtVCZfUH1gpnkhF/bhNS8AF4d3
QM2uJkaRh1LrxB7T4mWiWKFPDJbshURqMeC03cIsn5ClIPUprRTLqB4LWW4+IN57pEd+fG9tJzMS
AJ2HmQaNcBoU8oERf0A1pAeJC4jyiEoMP/CwCUc73SBOZLLG2vmd6T3eejV+brabEqaz08DOYkDi
ms/QdpQuRcPV7d0cAXRb3z6WIxZy5gTjCqsKqXMeZ34xmH3TYlapOhZE2JRlZBww1utPl1MXDFEV
mnGUUa+9e+OSfNIoLNwUcgWnPLzjnbcgQixSH0Nz1619TYKJg9QVJPdNiV7xdg2F1W4AdMRt3Q7i
4VPzcYzq3WHZjaiM4viVBtN7wE27RxAklNtO0GPpTS778Jm50IueYcuziPpLtyuiV/ZYeBXPetFo
dOOVQGh0muFjTVd1s0O1HVvqE7KNTYuh11C+DUYycb/gyMRIcf8yA8smSJLha9KA46JbV/zn4OEt
BIN49wrOiwnhV0DZInRaVIFpYe5BV0m5aAeCeUcQt6LPmvDDyPdgd0zkea7Ha0RM0yabW9pwtqS6
X5paaupiXa1YcsnU38nUNjYluuG/Wvc5kicdNNy8TU5d3NFQXGPefOWXk7K35clDLRyJHV7NONn6
fDVk4M/Q06LI6ywwJZaw9Aeg056++1wcQPSyFJkDLy0WVgAIDAi/+qlz9y9RivXM+rCqdGGK4yqt
RgX7Df0UKmhSkCp9SH8W28RbnwOaTY8zavCE6Aw050AKM6ITb+Xxtt14JDBzkdgUvagVnoOMPpM7
bfL1M72qG2vZ0QO+nWmZO2MS8Y9tDBwqf12eEcJgHy/Ulu9g2/+/afEI0HXjbi3yLq/jzXRp2EWA
pGtClEhX3E3zOy+686ueL8MnyOQJ/sIyg6URJQQ5KpfWmb6Yz+FtyQavDe7yNptPiRjk7Cfmu+cV
tnbHEYge0ql0Xddu6J/QNMj18MDd92CqccT7ZdVeaQyR0rbu7hFOzRT1nkWosymdkYRRVypeDW6G
Juyt8VkjqJTCT/pjw1+aoHs42xzN/JOLp5p6ag0iIN4HK55ewHTOXdlZyxLAUe2Ld/HphKB/FanC
GGJ9j0ixs3KfxX6Cy7f4FVpXzN6grJkrDB/4PibsDSIiQteZjw3MjL1rW4bhGG//oENbyE+EGfPI
J1+CRcy6RJWodPr39kAi4u9h7PVbA6myAxA+MUgBpSFZ3RBSSNzZvkx2y8tSpH3XMzuSDSCDiUo7
w77v9EOCwjZNhmo7eYvsuLzeGIPKfFXm2HIN4IuT+1YELwpYgyrlBIHsmr7PP1siasmEoN7OLfil
dGJiorxscQjdy8UJZIIz3nrRK7kK5nTiQbpvkjAyeIKDQjF+ZFHaq8psiqK+W/DZS0QZp+HxSuAJ
gmWRlGnjMbsh9TgiKWg1mm0G5+g4nHtkI/ygcxYttEguQMaqfD8kYFcNqW71fTf0MWcsX1nw7A6q
+CUgSRcFFw6smEihnYHuhJ0F9VlWRZv+VmY3mWcXQODttLDVDjSpoxc6vRE7h683NAC1byZBM9UC
mT83huotH1MV41IkW3FCWxAFC8sVBCQgfrmzdZRCEcY3VcGS2d83CcYARm7OtegH06ac+vRjKhqJ
rolkNbRKQwZ62+O1lUfc0NGi5AbUGWFJtIL+YTs27Wl4L29O5gOQX+lQxYrkG+9+5ElWIQxJ+wE+
dmi1NAlXa09+odC7rqKZG4ZQ7fNdWUodCrLQYVHGjwNKh8IojjDqn9cRRNtTj+MQL5LH7SmQvM1C
pOioDrlUhWR0hIYrSoZOyessEauzRx0DxIdpSIL+Hybv+g20v3Nspg6tWDpuL5NEaCRq5uQ8MxX3
ffg3bIaJ0Jr0jUkrlkXyzulQx1IIfzr8jooAdB8SFdJwydoCjDMwcohnqLPOetTRobkDNT8eoixw
IQfwTmY2T56Zlss7/4HX5kNPU4dzQtnXB+KJFZRDtF2PtPUWJyPOW72YgIBBzUYR3icwP/R08Fcf
lFkavOtewBMi3b5y1DSBU/8KdbCjWFLzO6KoQ5T2lPPtjYwFRVI+0l5bgG/1h/pbB+G8FB7DftUT
3IxA9nOe/74sgcZEBNvOeE2/NZclLL92EXeQTOgFL80vfv3SH/YTEMxTh5P6J8Y6DOJK0bm/QnvP
SbOE2gwQ4MvhysPly+B64IBz9HD6jOUuO0jY7RSvoBDurvaON/LI+8jUNGs1qSFKESE9Xp8BOpSO
WHgd+UR3oVM4NtEY6dc7Z2vwVU3i2Y6HeMiWemL+sT23/8pxlPb3+4MTAgNWYM67aCxidrJSOxNg
kBqUV4gIvBrlDyuqWSpGDPz3NM+v4qLxYoCzSaAePLLJyYdri6z6BPc7JqJuU51/D/Y/xAUFzM9W
27m1EryQTEZRyt9S+6c4iiuY9OCoF7bip5hbASnJ1i8bT/sp+YIr5vPFhgSf5hC5NOW5dTrlrIHo
tdrgbsG4P72gAW6yPBaR33qTZNqNv3Z0f2z3M7X7rax2HgWUbB49DZRr4b1mk6fLP3uc65XpB1/o
rAWdtzNc+nTAnn8e9DU50VQnTg0HRq3MzgyfS/HmIQaau7cxDgEuhpMh2xs2iPjmWUxrncJHOMEa
4l+wv5yb8UUVmp+Uzk1/VLl6H31GQz6QQPGvMy/IDLVhQ25DbZw8+UjocnaIuf6H62bmnhXlX+/p
I6hPx7Z1acjgh8jZyPYbShyKZ66gYzWxEoY7+87rmnkX92YsPBRU62W9S148G4g1ekdfOCDxWd5N
G7r1CFAyS/cI+8RP4TqZw3jYMwLjFs7Y0kQpZPtb+AEy66CGCAamnKKmVl7g42arlzGUgPqFh86Y
YFdAgaWlL22J+Z2JA0B5AB2u6hXRx2/CnWL8FuiC7BYBtVkLpwBDRkr0nxF2eETwykuaEEgpPj4g
EZNwqq5s3v6PdgSjoIXtFfyiwPY+nnj61wA3TrK6skuwDgVUa7EepOucWYCdx2l8DodjhPCw3TWa
+6DuUMbJtgPaRIHw3IKSj9cJU462crgPEGn9bWxO1mSI5UmUaumrcGNAW9Nn2i8fSJghT8SDxKwL
kBYFkC+RlFt6mlazDu5cWyJt1lOFJ4cEuZIdouK1R6XeAVBgB5/XZxyDe7aW8hyM/BUB8tLU1Ltn
ztAn39Jr2arKbBRgyo24SHU6cSX3jIFE9SFYs2uVB96gIO9G5BPVOiSrq9GFdNn30VUOEi9urnxI
u5jB8fYZoqfT9ZojlAVdeIYyB+zY63HiusMaeZTpqf0pbHnybzmRO9lGBFa6cIj4x7U27zerGCcg
/5SvBd5ar+TD6aJECQOaFL14p9xklYpKEdPOHSzCEyCH1w4QwkCZhULIUGp5Q/z4nytvOxa9w+LF
T8mVlTYhAQ8uuQW7+DTojwubI2mJ8qdHo3+fBWkaVAmqGAyhut0TgBovAeFHF9t1raZdIKTw9aPF
dGy2o/xc7eya4R6H4Xy9Y/XmgBWcfmqtElTVlvL2ccqVYNaDkGAy9SM04HRsWL2kNYD83UVg+CBe
sFMOLcE3so3r6TLF1XcUUNygcJRFL14EQfRjWu+ditojsKz2Et51QCsdOdwHpIWkWl8bdJ0Qpr+R
K54ahjDUJiB8UeE4rV4ARvNrZhbiY9m26AgnxTJurDOuxs1uCP9zwISH3/gIKKG4CTyo4up2x/rE
wBeN6Z6NyijFoXgXQTG1qa0c5KWykQSKFgJHzhXH6JUFYc2tn61qqDC75q5E1NXYFdh3h9Jm91Xc
DMzrgWTLkDiKSW8H1OLCRCUGQZPbFWUGc97Y6p6Sp+OaEDXx1VDWdYPzFuqseOloCsdt7cPMbDOY
WGqlAzERwrZDKVky34I1ftUZ583h0OALg7wwb9jFRLNNTNobIy8WpADoNRSk7SY1ATgInv9C1GRM
BPWxsVP99415oPu4mAyLnyENwYskqEAjaNK2bk5djGtvYdxWsfISzcIIVdSpvQa/dSYAa5JQydkL
nyhcrnakOy9zmZDOYaIvkNEV6DAmJLnKaLAKNjJ62+9dYeaNdfF7skqUHzepgV7WKwFP2ZeBww0I
DQZosCgdG6N2IS2kZwch04ioMKYhH80U41oEiwRRCVVvZnPmqQ5YsnbB1l68urh+uYxFenJB8Jrt
K9oqthSQ5ICaBubUNkJHMBcfgOn3t4PnEkZGvlaii2SJf5qNzgxSVXos3kKRkmoNJydJ8YBw7cCq
/No4KfeAdn+lp/ewoeL9+pQ05QcTdAX/aVFNqBC6jq4zOUtyV02PxheXkivfpmmB8z0AWDLvhtFS
jdDRdsWhihju29r5qX2YXf+zwLNfiWabbxIPFFgGVpWGBT75LCkSS9ARQZ9+b4pxI9UJpW337qUH
scQfE3PWNNo1abPAnmT5LWXQVuij9GMLqFKGIdxVtKL9w2M5P+miVwWBQEj25kDUjzR7P5/oMw1o
3r0Wfi4IJZ0v+mDHc4S5wCdr32K+wVl1MaRyjM9618oYTjTgaVlPznAa6cSKaNTxqEl1B+JGEWt5
DCKWO7yRzSpJp9VSD8KOPfNjEHCkSyOGCWxpRDk8wNf9TvJP6mVF4/XKD9V05CuamZGqEV5tRfsL
x0T/6XHy/EII8HWF3uq/xGQAJEpJV+K+Va4tUCr84EjSf+DNS2ajl8h4Sj4MPSdHxShu2iy7x9NY
XCE9vDRVktj2IXl9xbPrsIEs0LFXLSgdtSsPKrYO1wYASorC5+4bKSE+gxLSQDOPQKxY2SZ422C1
zHEf17WATUYvm4EUZfbzA4r7iBYet6fsaI6r1lSzaFohyXQ4FTQwoUUUzf59bwYSUNXK5UdQmHfc
S9945iA/nQ8llqGuHRR2JRcPHfIQsdFWsISEsAPwdDgSCkXDThf3eDQ5sLOnP5owOOQEvkDYwvcj
Bxr9FQ2jMiqKq/NYZAzoXBgA1IhXIpVXvY7nQ95ahUTFqIz2SPmg+PB/CakcZKBUpvXZe0OOkw0a
kujIHRz3zjVibmVVtbHPyOBizR2MJEXovCBXuTaSQl5PhGCCell2RHuhVDtes0uq4BUE1VWeRoCt
75AzY+cEt6UKlaITRKgnJLI4Win/f7qh2Z0Xg9kPMOsAYPk9cRfCMrygvuhWfmJ2U3J35OX4REtD
rocSqmmeoyDqxVLOJBbL/WEbhlJh/HEN7KXl2iW001ftQa2QqAwTJOTFd2zoe34sMhvY8yVFsDuy
vy7TyMHVhYpotYgb1/ojDEt6mdcjgFU4iKmYZ8lwz3ulYRs4L2VfONt2QKY/EuPqIZEJVw1rrugA
j/11N9Ww1UmUGhBpmqvC93VooyH7tdAIO3X9B9xjsa4M7HjEz8MjksR9tYw3YBtJ2pYIBCHt9dU1
VUPd7ecoYhGlPh4bkiZKKPlDCeYxVNulMOiarkKw3DzKIUyxPioVOsfNupUBfXq2SL6SY2g8vdZZ
jvR6YXPhhjr9yBbsohZSNEsmIEsRXD7vROyn/nhtDK0yQ4N4fG4b3DoJ1TTFC++SSUaYPvV9u7/B
rLZZseaEQTSGrWr9UaARSWBhUTx8ssuSXiSKY7J85HemefqTrnNejjnypqv1MctNndisYRBfK/q4
cxYmjzx5z2pnfwgiQ1FEEK4AxrU/0LHL9SDIR4GTQeEAZHZD7xImtZ2wHhmScgll2qNFsB89eFCQ
8UFsMYYndZTo5I3U8miX5nn7QsJIZUrnOoCMgb1Pe8KcuX+FWVmJJSN/2mD8j7nSfP0ZKYRQlnbf
lPpGqshnR2uEzwvNNBLCwKIXprdoUkQGjss5JGoeeTMLaabjE+mvy/bl51089q7TLGer1bQRoDiH
8XxiaaqiRbJ11vNA0lKlnK/FX33OiHhky6JFRt5yNj5BQ/svF07DZYJNH+MnW7NphlgLHs1QxQSa
YctvHN7rSiBSRzgpyUOADFTlU0EqTPba5K9mnOLCaVpdIV5foxP2Bt4xxl30tlqEg5kIPZC4u9pM
hnGDHcRdy7NweOVucucQ5zLphwRbJFA4fzpKnXJRtzsB/39o2++CqErOMso8/lGbUrY8R1oihHKD
Q7LLp8eJ024Jn7jjyeAjdLD+Ro+maDixMF3wDYB+0U7jB0x7zGZLgxzE/y8ZLnoPR5QcNcidc5zU
FHnYAMvoJ9RDqi7EU2MZFR6YPjOWfzMB4H+cwqgRPIX87Co0SHydbRuqn5Fx+wvNsMz3RaLotKxV
w0anhF/IRRwBBkSP14fs8f2st5ztfHaDu54ajmi4Ff6+aBPkt4RUepD27hvsNPKxkIoTD9MUHDQB
nilJ+STUhRn8+P8MfaQZf/ED/qBfG6QEX4anBMTHkb1fNQDQ2Mp3mLjBkNWlR8t0Ro0LCZsZz2/j
3JwzxepIMpLlJyTU+yQ3rJLzn4wJTGW5c4XikTH1WKFoxmN7Mm8/M/YlbmzFpVCTWxfYS/If52Kp
9uh6Wt6180TFez+BhUeUjl9FeEur0KCXhve6QDAEmtrbyQljpwOepi0RdODv7bXbMW7t3eSixnqE
EGJgrxxSi5LfOpQE5eAHMUv59XYaNLhiV/m7vNvJp3zQrD/IjhiwuEEgckXAupLzJm9Md3j6H2Ng
VZW4WlS+X8wEP/S7xnhYq2I4nomWOwQhoctL8XdCyfkdpPqKP0SIueJVsSdyjT+usCI0QUEaE20u
UsYBT4URZCr6h6YYezRumfP1a/tLyj2OPUzz06um6Pdro1uNv6jowWMhcerDIV37uy436FePmZzH
VsWNjvExQ5+Idt1KzF/IMdZbZONbwkMgFGcnXLDE7TcGZARvAqz5bTbbDcVJikFdNz98KB/YqMAD
LtZOfvOhxyYml5VQ2CnnUwRZK0bmJABwV/+B5SvkJMPgZmVP4FtQK7NsmvOTq7DCy1O5HNxJ5SKa
GtQyKzjZzUoTrcOeKnZp8kACAUnP58rXa0slqMLlPpZfOkYlzIq30lk/2GhTqKnhl8n71VPmU614
89DpI9f28YhQSGjtzjXrndGlx/nJS8zxN9RIe2ZiToSlkHcZpAlzIvQmV0GOqi+SiZRwuFZVAxq8
BLyZ0tbAoUvkI26jP4Nkk9iCCmJKh14VZI1xWFuVaJJGNPDudYSr2lajnldfA5NdsyisNZmxr2aD
90FrQIHQ+upypDuZmQqpJHi7In3l1Wv1IEFtCJbbH5sUBjxNrUUtPyWcp8BLyhDBsfkqegLnEudn
p+bKEjBNl4PkfqqqZQtqCZpx3uh9m747KdZVtkdhPz5nNC1leM9pplnaSKbZEuWyuy0WmvwECRw7
Z5G+3CMIdxTS5/bhEpUkOfpq6e/WIX8EzVsQ3WZnTJxYaaSjd/kQ/8E6YUcGNPwipFvZwTgvyxnr
ZZtCuxwGCxKgPcQH+qwalRmOSD8hoG5QEObStzT7Acvg+TRe8MvAS2rc59Zj6LTFOlQ9/Sy+v0ug
WJDCGQJRVL3IxDPH0TMqs04X7bDIgeJavXaL27xHXuU3hhELiUiliilQa7ld7jPIyptQ15OrdYVb
qvJt/pIQW2B2h8vYETUQRSRYIUdy5I8z1hND7isVlcXCb9I2XvZszcmdjWSTNjcQppF9LIQtwOl4
2mmCR+e6+TmO69vykPhTuGjRdVLYZE4Vtlc0L163LzfMfX3OOb6YdIsXgHJiU9224bP+P4UMsGB0
HFtH8MuO5KOAq7M+E/wr1wi9k0g2XENSEfLkLnf8h1lx3ceO/Dm9aSxfosWtmeGRLbjJXCjRU1wJ
05tcHDnrOSMEm7UIT/ey1VPF0CRifE2d+d5+MJ/6fU97Og8/oUCHOZNDpti9wqv0y61nqreBPc9m
hCgRZkwzMCa8bGNtIBf6ow8JbQ4JO6gMcVmA9tdd6i90AKP6e7vyz8sYvA4r/rHYVQ0zF7Isq8WY
einfGhJQV4KqZ0w0jQjI4okY39cMAVSV6TAIyvRqAIIkGHbrgJ9lqwgEb/yiEMsHoytnvhmgkwmZ
x7a7YBY2chXtH6dfNa0OUDUV74XAEdfeP1lGcPpyk92pTEJoIguseSCLzyF4bP1fdIZt26yP32R3
00mpRWmjzX5htADARuZUgBBGBtPHHIOGyceHeDGVinJRVZoZAiwcis/xHpypRpI3tpeRymHNdA4p
r0ghJo+MUV36Zb7BijQhT/dxjDhhJ+AUmXzLeJQfXciphgla8pgcUUFXbC/5nOrEtookqISdjv1I
GpvRAgQGT/ao0Lid/h6yLyeJzIDivXII81wa5Zcyu/hG4fsc1qZFL1IVN5G+1SSb1syueS1ZVJ7R
NhkiO6mQG1PZOU8GDiHR5PRT07NRWHIvygbFnsDb5tg3WWdmL8rt30qlKlyyz0zBCEudLEcHQfSK
BQfqZ0EDngZCEEWgSek1pMqEj0dB0Hlx9bRDtomxfutN/5orFvq21HaG3YaGQocdgBvW9NHsP3AX
C9HYWTMMcEq2kkb0/8GRcHwScf70XE+Kds0/qVhEPO8GzkhCJi8Lfr9uvnWR17TiV4pTCbLR37fK
xqPRTimX+kOIdUltDNoPrwjEC0+xBEdPkTh+93hiIA5cSZPmiEcJNIzY+SblqDWR+SPqa3oG7GHC
3sxBj2MISaGPpmDcWMHCLqqs5XKRDlZdQnRV4XjKp03qYaRzPL+q7syQmqvHOGl/PrA7GRG9zm8c
b1F/io1vDzB/aTF288qi8gOOPorTIVddooHqT3rOQm1lKvUR+kBbaBVg18eV9ws2FhhlmE3Dc+LW
LBu/1k9jvIIb1ntrImp149jbmtoHsQy/qbmmedXEaXp47PizIh3PNmhW5RUH8lNxSLvFc+56W8xs
eGlpxywYz9k4lZ6OFwdPAC3OjH2jeR18yyIePL4u4gGGjuG1moZfxZU7CzFGcEydhAYoV10b8kC8
WSCDzE7tETwExpKobouIXsk0mUx4IoT3DasRkqXnf6bDC30YiwlaAnFnHamVt/YOnyP9KYZbg8Yp
LlWzy48U0kSp7V7veT4RrtZ4lPKO7Yi9lTjftaKJnXCWVqfifCGRtb3saqqhrok5RFo58uAbieKh
jstSh+cDW628nRLLO7UOxEteSFFerR2cAW9EO+WMP5a5KD9XA1pGnNFTmjRc3Q+BPcUWO9nj/M8d
ABEJ9mWRReacVA/bD43gByMiebz82drzkKRJuC7QpV8u1pYZT5yDKmdZVheQ/Svn/mRaBIz1iqJL
4ualOoXSIVHGsr8CqzoyCOVawK+VIHAeVICiDhKA2EOXV1EIYQIP9LtnNneIaaiRFXSiT9nIAD89
oIpfVg9M5WWQs2KRTlGjaeyupN3E+w1BY2l5QzrDIDbgJVaiik+apSzsmLZXWzPc2bPKMITF+jfF
L2c9PLTgxv/PqYJPJRgFiz5fs599YpYuA61MqXiUCBYrcyXdPyezIZs/CFpijrfk5Fhi+5y6WsBw
3AR3v5LRdSmIXKgVik6+asJskh5F0JDWcrcAyp+yt+LCN73ogzPsBer3SiqkvVRm+NBQ+VWhE/ba
SyHy6FD2Kj6W+2igjwYho0Y1i1ixlP+hiTbPD328tQEL9au73BhodX1DuPyRZB5qvU0ovwQ+bQoB
ZJrq2rw1VvgQhIkCMpIhXGIiNRY3k+3o5pVjJ5ITWCWy4SUdHrRG49j+4Cfm21MJwV3O3o8s2IFh
EJ1e6MtxX60Sj5Wkl4uN47bPxSUdV3gUTCxmD3sezPcINedQAI0+vjSQebAn5Sumfvwa3V3y2lT5
WARTAsWd50g3a41AdMjKmiVLZabcJq1WqgFwoHtqe8ePhSyTK/kgO4uCuXWALYEG1AKVlYMhgf4/
XTB+jZeafaZqbaGX5IbMyT2IjI8k2RtRsDfJsAdnXCSRKi1XEAIBzh8DIcdNxg2Iq+1L4ROynAQR
bz2iZP6jwuInevKlaeftnGAmrThXgjonYRyHnLnpIb+/P4eWh2xMiHvsqPh9kiS2sBdoYJwO8O1u
CiD22PmFd2xb1B0qvLENedGF6xz7YmpasBdF0OClQQZ+hm3ZUveE4lT6RWFD6smn2ugJ9/QulenC
H8wmjk3HZD5mXssPfQxb58IpyUKTb8MZkF47psdw3VAwGrRFURMThpKpsckbMuIxaDfqmqwl7A7t
iJdxX79eOs6oWNE8WwJB4a0T0LSqNzOMtnYhX8ouxp5Amj7Goojsk20c6JkEbFUFKqT2hEJXh3pK
IjJT7BcJvCrnypffnH4v2Sr9rKIJrFwP0ajF6SqBKlkquwdupT8g85aVVFYO9IxB2s7z7/Sy4ZzR
5JlFL4Xec8tq1D5s79u/aTqsZneCVYpPfFMJ6NI6sB3ONtSUKeK5s8OYQ25vGo8FCAdt0I8JsI0B
Vsv/9avnamOP/HqKfpLqCi21RWYHTG4WzDva1V6b5hpGv41SqOJPaEb8/+uRGeSLQNG4MNPH0EyG
hAYusj9sm1fR7GhQ2WxnihJPja/PoPWbEmq0/YmQ7ovzcBlU8/3M7QHchgaFwdllGt1/WwvQWllM
nfGUeT9oy6aF6A2hfm+yuuN9YVO9FjSZgHoIwL3dv7P3zRk6c3bgaJk0YiRmsa0wCG3QGoX4Gdny
6t+G3qSAjSCUIRCW47CgS8vUjaB/M1zEnXT+hSD56GtcLe1VDzoMsGW1VKDTox/kY86y/P2cz9Kl
SvpFYwSE9Xcfgl33qUc4pwoXIwiNXQcVX1x88TYPWomr7x5syKZqOQTlMjtLOgy28m+VoeINKe2f
Z5x5XvWPKFAexJ0puKXsGUY8kCts+3uOpfWErY772bTqZNJVs6lUTw787BMPSzoLgXr8B0fh6kUL
fGIhm5UOV9EYEYEb6qnTTSdIkOJYK8be/adg+4LxGBvGewKKHCMGCXdyWnInJbWCb/ZWcy0BKFif
w9v7oB8g3gO7oBpyaIdXedaksuQT36GxLmzVCb4UEVELII0SR34vR2SVJ0ZGVLeaQUQlr2yrq0eS
q+hnskSzTXbNL7AcVn+vMLM64mN8gY16E9I3VyEe14lHB/mCY8jrvpjggRKd+3vVI7ivqPsdSqf7
oP48Mdb69TUfoOzsdBI4hRY4fO4E2Ii06KbOS8Gz0P6ORg0p7ty903yvwQ0AHPdadWecDGxZuFpY
AFIaYQlnstoVOMN7YRlfjwBd0jCzthf+4qf4T08VK8IpCKvxHG860e9v6SFj9ESH3AMHu5LVqwEd
9tAjtBBmefnm/9RXBThXuslX5TiN44UGp2izLfLBWxrnfhpkjXvOb+HlpuLzTkwuZ66+ggJnKhz7
Bh/Jx9xzFfKz6kjUWKIUTxojELlfmAqHM+lY4GDy3ciVThYYDa/NUaV0QC0PLjYcAssrpuevSENI
RvyK5pMSne5kVM4Sw/uBXea3xTdDzv17Tm31P11WTGFOtskle/How/hCriaezn9oR0Ga5+kPxM/+
kv+lhz8mONyN7mN6N1+rEQmaL97KQu2OFrzQlMd1Ta8/YgD8+7EgOpQ/eiWqH7Vqr5sv6IWIZth3
w5p4z14FEitBmi64rW/TQeP9t/ljKJ1xClttcCg0LftQ39D0cRyRk8xRWDX4k8e1tJzU7lvYe/wD
TMoVRXJwvvWApJI2/gK9SsOug1XldPrKgTK3BAC9qY8QjU9F0sGh0GvL1wwIMby+zEg/gSQUmEad
3QSEEPNGp4I/ExgsJV4WcqoJuHsgBL7X+Dptp/lGf3Bs4UoFFO1AMSJwtAbpluGrb1LwNSbpP0Y+
NgeqTS558S2tLgHVkrVn2UgRBEPhKoXNiuluteJV3ITPrPONNJXomYpYqgp3QD9teSbSge1lvjNO
dyJQ29uHksLD5+r66cXI/6Vf88DVTYgTOCmtRO9mp2r6bX5tkjRfZ9qOvAmLSXx3XSB7t8EhYD1x
y3X6OkWrNctam8ZGvZmxWt4v0s64WF8FI2dL4d3zGaFP1s9TFFIvr4dyjt7cyWlv09eCk+XDY82B
fwMQI2K0lpGWBl1aAhOL4QkK9HpTmEkLCz5Y/Nzuvj43gYlM9CEtY9DXy4jRDa9oiO24fJXCwqK8
lec1LGNPJdkdZaAgLGloi8T3eYqmXybkT/Nytn0BqxOD2jY6txpKkanmzKAPna+qD5RkEbXB65uL
i4IFjKWSH74XL21fwZrj1cjcLOBzO4TYAaZiBSoYtpLJ88CQ1kUBggnMsXsJ7gnaddxrPN+bgHKb
daRCRSl7W2Zue9wP8WSc6nhbu5XjTczunfVJKCU5oENbwRhvbXgMDl6ooqTcSc6Rq3XRYbcDCbKG
E+CEdknyxNx+zLsK1Us/fflwi0TcjAF+zAQAxZq9QdT4LyoKh9f9vbG6I/VZU8IIhPosBWrjGfXq
3gaUilDHMpWpR9Gc5PWNSsxSwoB1xU52dWeIc/NYOxBE9XeBq2w54vDQolXEOx3mOokMSZ+Cdgnw
wS5vuhFHMndyVCflA74ZkFQVrSYNzPMx23vkMmh1EFyGqMXBtn0S7XIHG5no9xJtFBCN+6c1x9J7
yjUVB/3MVG8PilFCbeNGlA/wyI5izCr3kKLUeXtpe7VWlrAX8v/gIP6Bc4Yp7DFQChjSlbC2x0nd
gKTNvD0ydVZe7EqhxjgH9bR0PKh2RGe/4yo85/aapQIK2MempnILkES2kmBhIprXI7oJPRa7Wws+
Uan8Mx8gy1FvSrqM3ye+r2Kyz/4gY9LSEmyO3bii00q2aKx8plXixL+ENMDXFhqNP/jmCWQ09rk4
nE/8KxWNH5S7kU3VeRwAGx4ECqIXOUFZVA75V1jmdBU8o1jrj7BvogKN0duKRCgmXSAtVMNHUNIe
Nsj49JqmsyTHh7rzTDwvnqiqHR+L82MpqhdBbnbHXmol6jHG3YJs92xOykDPKP7S7IGGQ5uBxDrn
u0kzWMZwKMlzPSfPYZNRBdNykO3APLn+fNJw7S6vXTjm6QWJm+MGAGBz5IQmAAWsBM4rl6ua2iQU
TQRxn92g7ued/JfHc3issvs8KBWtkfyv4aIrzrD9DOAJt6ugqPw4pGQ9rspxvX0oFbrmsBt9AcTf
AK6IKqLvQG/RWaYPtTJjxG++6pfsWJ5lSoneywNJCD8J+hSyhqGklEraIGkoasEmZd/QL6r6WOTj
++K4E7nrryp249J1AuBmw/bQ6ojuB5OkGU9IT+xiYgyW3K+gPujndNybVX5Q1XgTnvW5JcLw7Z02
k+wgwd66jXdXWJnIV0+D9D4S+Gei/WLaiiw7c0B1pr1ClMxzgm/sc/T8OBGLXBZj9Xjyae0/T+ze
K84xbphCNTO5OqxHZiMgXdB5+qX6411V3dbAKa0ogIdXBd8VbM3DUytVAOi0X20gYlI7EzH/Npu6
2IJ45E5zPJY0Mr5VvX6lx3dphp9bNtALI3ba6CHYSdlaNJCC0kBNb1b22X9MbkOxl5MXcEurKlQS
30CZiaqGpgws2Hg0btAFp9Yv7gtVveSZU/Rp8qmzkK1axfxppIKnEWnJA9yqhBPQecO/wsp1Ellw
smy/BR++s/RcrxkSHTKIWlnI35eJzmR6gh9QdP9VR4BYAaXi75aXk19B68SIo0mU/ipAMFFWeo5s
DVhEMhIn8uoJWwV0328k4DPlQqnc1KLyaOYCSdFYGc/i+VnJDuO74RJmIdaNAKfnjYP81NLNj31q
54njqRUmXJ1fdob23aJExd5+a7a73SwWJKRrI4SifyFdpEMDwdjGilUnj63GQTnAKwIHgqT8JCX+
Zg2Xzm1lzWHVltJkkJCY0mY1wKPUtfz9bsiTPLIRaJOkDDEATEbOSKh/g2l25etzwpeXaHpX4CCC
cxB9WpNhoKigaXxtxyFkw5GPm4KoeuKGLEIoUXF2OCS6TWXc/qni3OABKXHHlWm2aOqBKBlGR4Tm
pQULXam7C62Ee7i7rw3AwpOB3TKNSmSIaYzz6b8qTCHC4rpn/rsQbIrkYCEj0HRrR6P94Z3+RO1U
8J9sl9OYbKUBh8N36EvhQfBuWk5bVK075D41huJQGtb/Ti5SX5DNK3NQPgKKeOdSSBXOUcLJAvQO
XIWi3axpDg6UOy7JtPKxdMLsFPDCYm2+pI9UaSY6KOUGn5htt+ageT2H1a+OLZcQgJ57Fyy5K9dv
b/45Xu12naZ4xhvcu9Hmrwj2Ud2kfuNlh9xG0fqaVZFgoLLbEMp/Sq9HK0PRVYZuAteze2/KpvU2
t0+0rQOBMZfexzVSzmBdFz/ImBcMc0F3d5JN8YIpu9GLDUnOUY/M708OZNtUGuMk64acP4wxjDpP
GahrAbLpJg5FceSXKDaCnSqUN9WWYvcKNFSZay0y/GfYcpnSNV8Pyzy9kslLsmiGwqbX9BlTWonf
VBYU9XGQBMe48ioEiPgi/qhNkTT3nmWOyiJy/QxNdWBOUsHl0YofLzz01NfVxTKjIWJnsfzo3W1n
G28ujxCU7AdNWXFEiMammR9jdedZEoUwyuVtLzmOeDwpYGKfSsu5BnHUxiOUXl3vzO4ZzlAXFuSg
jjBDobcNuofrFcYsb8dK7Y/sbgy2K3k2cPA149QHRXSOBxcW0Yw19orwXoDPEh8cutTv+zwB5o0A
yB7eoOUVYX2uXAtZt25SFr5pXNc5qiN9GySVulPE8cwJU79af8zGkt2j9nsVEp1TexZsl97Pl197
/6N1DRUOMkyBh7zMzv0LLnwTtzJ74CeS/WA3uoxhIGb3eFM0XS8/V7SziE3O+VeI24vaMS9L80gD
hDNkIHKDFOrFlcvuno3ugC4NyL9aDHvO4lrae1nHWyaUhv14cjWpdY71TXO+dDyHYYdEOrJTcfCY
LVOttdVK6Imxn2j1ubEODedV+Qp8LoorSRk1y6+x3KZVIOs3VkYzqBHDdhy8TF6H0cyrLPIw3Ci2
1s19eXZbDEUQEOWtKDgg0DZYQ+PLyPwcu44Gtmq8rRzq/9u/1Onbwy7c+uoqN+XB6TmvsT9JeMFJ
uHMidgc8r54DMgBKF208ilKJmtKs5+F5C47T43J2uz+9gWHBAjeXK47Q0vuGDLG1GN3u7Qi6pFGW
FCKHRePan4KelsNCjou6xd1ZS/1VvcYvaVDWNVUdXNInXskGVeeS26RRFj1whp4RFE4aghnpN9pk
tCUjcSGwb8gW5Af76LzPUWRleDs91y8fIBLPLEnY8Wxpqtim/fbCJYE0+lB1CBsTPKSWy/+ePIlN
LkBTaSzwR+nz0irsjkMV6VlZKonR99H/E8DtFR/3Evz9js54CK2qaWqzktvmeX7OiMHFNcPUcfBl
TghOBx2XwAjnvcEK3uWsB0PRiJZtUJUbaCS1OGsV8P0V6dM6NUKWn2w5xAIDx8VKZS5eOIjD18Dt
jJEFJGR8HS+8wlt4iCm02QGrzJvpOVhxTVUf67LyQc8WHUExQwM9teC+2azANeK8cMUEcxfgrjuf
voPT1EgSQothkVDPib6KmUhEcW8OXjo1eBM0aZXdvnEPCkVVBm4GLPUhhlhoZjn0kyqb//n1P8JR
7faMb7b68e8zCfblZ5pO6+SndYYw1JYSgSLngFZjBXd/Fk0WLvFyiXjCLlf/6kPoJuTeclzgECT6
Uei9eKQkF6A2IGTagonk6L3EULvzJokNwKrfvdKB7SP/sCP/cin7OPOjX3YIAESNIeBcTtC1AugZ
gu0tgFYFZ1PRzeGzxvWQT1TILULxfpanAgY05fFXQ5UqbBdI3qRGD6DZhRjhZlmpMmChI33P0E/y
mZ6LOtGxfXGnRZ7vkoKsNFPbmBITOtATd8CGcIbH6yecFWSs1y01dsv3JmV4JFBQZ2HJGr0Udj4E
poNPLR0bUcMnzLdM+NIlaHa/Eef5wbzXJgSYaPJ07Hs3fgtNO3pNMAFDu1+MpHszu1O0hbdoveV8
CRafuhjKTC2MXW2zA1SlswEAIqsktelYvkuoYqzOhz7ktONGpEMSkMaOkbJOOtRRu0jS8wxzJc8W
NI036n0+OzDBzWWeSOfj/oQHhK9zKAdiavpwrcRGMY0/q/Bh13r/nhFZ8s3OU1n2VpjvybZ45zgz
Z85+NH309SI/PAwQTNsdxf0JQHytWSGkEIkXYLg+wK/9ygIYkSXYIFK9bn3j/gdtWT3H2UqFL0fY
c7kTwsnMDMfU3EbwfHTDp9GWi5vmgoVO/lxY26f/NZe/8Gsu2IZOjnlsGWO/LjgAvjqKFrBohPID
gQG0GGpOud2vLHOxybmiyaJiDBRocl9PYrgrNxDvZSbqVBIxfTJ497GCRaS+8BXO496ugh1wJ0aB
GmKlF/LYQrlM0KNtlGSBhgQS6A3d7jYOC3r8dm20MOTqxAe4+lm7MG5NQwQQ2WJPmp//nT782RuG
qJFhZ4vi8NhbULSbqsYFVtTGDVP9U0eq3yyCo8Ja0n4drLp6UxZMyknrmkwcVKSu9aN90Szl5rD8
+E1qvp0KvjR0jGZrb3Zx3ZBlfMVrG5qvvLSD6IruqAv6O8R4WNREbTcqj06dceA5orD5tWBEotXr
1CfPQIrP7/ZbFpK2BOloOCLtLaTSF40ATJ6BViCKENBLYRLkYL8V3GzUJPrdf4Ua3tWdOtk1gYtM
RKgQosmLdOekkgG1L0CMh0zVCaq+agSbF51SRzigjeuMevPNSbCdtcHNW/vxuWN0Pey5N7cQNdxD
8Ven4oSAlkV+PIwONLqsIwRJhxraguTgCFyeLTJcp5eXX7qWLO/7GuGBuWjuHzOk6Zwu+8NGR6Qe
/qI1F75gvtg0E396qorC252ghuQRMFI/6YmDKQ8vFGBERDtpkdYBTIHrlGTaaH/8MYWmObMz/ce5
ALOMWzH9jDj/VlXeEBL47rDoNOeJQLW7v3JaM1rARBe1oep+Z8LFMjJDCyv+jo7YSaAdsXUJu9QJ
YHvTp6LwjUVfHdByQ/ldhJszPOaYQzO3BMFXLxcdqj5+YZPXv5XXoNCU78oHxFHlIqMfDGlxx40N
+rL1fmVkFR+uY4aglOx22FTSVfQsU4J2sGAvObf+jv9klXajiitSvm1cTKMc4z6RtF0mb8xNu76B
fzUXC/bcqKY7JNmccII9NAaI9bDjDW9x8Vb5baeKC/om6SEo2gEPAFyWbX6H0La8wuV2gKtdMhb5
3Vbbtg5/ktUl6JApcT6b8oyAekwsgF5zYZn2c7uBhoKsS9zjMhAjUY0wrI5QiY6wM9AExVMF7tyL
mBd20HFmygWCmAgyqYWZbaRW44EpRTZeMA4FWL61O38pm5Mqm4wSTgpd2gG8KQl8lV5oW+jUtfs4
a6ieC1KVeBvCP0Vu6vrkTXflpaucj6UZz4lTdQ2mGcd8RYnPDv+sBxqHrCUmTxPeTJLODO9jgOwK
I4QYXxsOCPgY8okV+IsSJElCusTt6gsjMzXB/4ZMoQZ+zbCYwc7RfVP16F0EqfQUoam78xX6s0eQ
a2tC3BCVvhasU+p/mCSe9xhUYOFH5wcb071xg3JocMQZ/AqDgefOclUm/T5fCJAgKjgECjBmf6Qm
Sb9Xl1bkt09+Jz4xpRL+uYEiOSAMhHzqHT8flUOy/x/uVUhaQSMP8QtmrN1UGGF9BLfHV/9y0vYv
npU1bpx8duWJzXiDL/huzh4hNV4DfY5jWI9tsw8ojXSKaqnT11nQY8ggYb3lFXbrbrZJ6A3EUtuc
90iZVEREH9J7Xh+964YvsP7jQ2JsqDxlIFVOdb0ye2Wz87mmJFiHMEgAQsdSgf/4QJCNFgFLOS2l
UA0lWrdYpatxtzDKQDPIIXtKgo7c+tdhfQuR4g1TXMxxiFxlOjZyMOLbzjQpvxY3EG7Pixl8Cd6h
NWCprMInW8jX2gi10EbnaF7MxIb/QrWqmmz5BOUcFPouxEbXtTEA1/GMsoaqumq7gPe5GRaDqAYt
0wwJ5jsvFWIsp8+MMwREA3cdp49MkFgkvGxe05BBYCFJMW87ci7sg29+NPHS8wdwl3CFnPdeVeCu
kharlVdduj7oCApmim0CZNTrkN/5rVZp9Ld+1DY9D1XDl6K5MSH1f7ntwfvccNhEMDhdmG3tNi0w
HwlEJlcmkifNumfSxJ4nMZcqIbHIhFQa27RF4mbZl9HPse1EoZEAoWXrLBD9oIjUD6JTRFwpmo37
2ef1cPdY/Brcb/qhh4ZX8X82a3glEVRzBIRg17DWLiKFFfCFigNz4gizqtzGF043kAqPp8UqqQCf
lUlyrvuDT3NW/zkHmLA5J9biRmz3Ygiv4WrWbE5U5St6WH5Zm7SKRbBe5mw6LFgEB3H9E7hC/HWR
MugNfb7oQ3CbTMhJKruKECw27uhDsnVL51Cx9UHsMhCD/onS8lfkaeeQomb4aIFNCpk7lz6DrCYy
Pn1pblmczJVjr8ISPik0NM4tIqGQh5zniLvE36MV1niBmZb+vftM2YqYwJZEIGoJwIJ5CtbZQ62o
cS7by6crWMfXkIHBJSeLjWHSnYcR79ibgKzGoWfAHDOFMF2ttVbZ57LTfmnIATN2hTJQPS31nCTj
RTtwyoaGncvK4esrj5xtF7lr4Uv75BNxqp1QBQ5I/uG7aT4GP2rWxomDX/WlFTj5ve8PKz+j9Yof
C5wOLILVG/i5BPGLpPPZ9azgRY/reuv0dgzFo89T9SAwnxtORQ0DunFxgdJv0DgSTduEMN9mROny
jYO1rT7Wsq7kCDv3EDi+ALiq5/L5iEyNpbkD29HtxlU7JbWq0c5leEii216j9+74l9Q9Q+oEhXEW
Qh+fzwRYScA2g3iUvc3WnL2bHKdJHGx+6Zw2Egy4Ii7AZ2DL+Tt5JQ6cq2fyzm251iOUYXR2so9/
3IdGJnRGNjE3uUvMzA902UJsQmaag2XiJXRHwzXxwFTjjhhlvsw/l32x/M805C7ksMPPw4DutoEX
DLRsI5edgOMhOg73qv5C7Tdkr5XN6GnMcFZBtsGFrmIlNhqj0nG9eoQt6r+YVWtSWR0FAfGLP6an
Bwwo5/5GElJvgtADbA5OhkxWtUvuxtnOiYNs27rsoa2NA8Ru9CuJhpGjiIOO0nVT5INW4lpJyX+l
96ECIk7AHwa5Z7V2MgoPzZIp6WRxbfXoMRD1WJx7wGLK5333tyW7v3QPIedx5i5NmoPAviOeclhi
dtghycOCBbEAtUrI+GldwU4zK2dlG45MIXuLJawZ/jeBgGr3vUAeDhj3dgk+xKliLU8+HQsVgbqc
VImud/ly7bPurltC7CONPNDLyg6VC+LwbBKdOgVcI4IE+LLAK7a4N31WV1q5JYVeseQP/TgjRuhV
0auLfWmCI7KUtk5IspeSii3WtxonAnD6vPAJ0kMDDjh2pMybs5BUc9on/kfi+O00KyuCmaKzHoHC
lfxeE1EI7ubmYtFbuUOFhhMuhGVv5dkVKbrxN9pXykjjrs3dDQmRDduGcgw42JK25Jw+yENCac/p
GPcCAS2JD0Ibl+eZlXgrG+Vemwh6hKdNS+Nht+udEu3fr59zbSfowoWyZeSww4bdjPJopmnFBuHU
7llocEUYib6ce3Q/aKU0JKVeUAMZe5i1sApV40icHL/OE6M9TLTEi0mNV/nbsidtAU+HJjnkOGca
zj+5IDDoyv5Bnqkl4DO87bd0kff+ER36+kV/KEXbqQcmgC4QbCv98HTa9dUwlDA8kTo0AuOS4Yfx
TIJ2SXOz8L/DWFXWoHpnC51DAX1uq1RMBc6EwQ/lshpG0xZuwIv5bLZGh6oEk7NS6lEFJP7XvwpV
2coWSWB49KArhRVntdqrWCIZWVePaUbaDPirKUKXgSQMYa+7FNVfSnb1iQ06NTn8qZZLStwwBZhB
6a/WzN0sGSrskDtuZjh4dHfUFhzwckQ7duUD9QlwMPaGrkbySHO0pEqHyvr1Id/7WApl9sUHARIo
1J0Eo5+KO85974p5KAwDvXEtW/mx7LFmxJCWdbKbabUH6iMaEST58jvadYABw4XzZtCDPocPRBgt
CTxCK4M0fQDPv0OZrZ7k5KriHRF9iglfD/a5AUdhluLope3SLePfb5FHabvhpQf4BaalEyRdVqHu
Jff1v/oxKHR7sebOEEUa452WweiS7cWUlZVTlxxfkxyTqLluyfS8cZ2Pmd/FwEgvl1PtrdRQRpjL
0bpcQWRC4H3aU/cFhFh+44flQh7tq6P2aHyWBzlpAJ5tL6+rJTNwDkuB47XO44ELmiB3mbfmPHPO
kgNsS7AwQiPki7+olRVzP3ml4PnMCcQgdUVoRg1/tfjWAYspIrc72zbSfGFAZfmDv8ND2fAFFLKN
uMeLy5n++v7v8bQQteM8jyvvXSM3ka5vyJE2gcnYZwko0DGcbovO5M63VUcfAeoJEy04dBCm2SBO
0OjyyoU2EdtWPCB+eS5EFxSWVRPWGQ3jVx0/UyTftkxTbiw9gg1GP4wbLrVlK7VjfY97CHrvCoiT
Be340bbXjTMwhQr+3u3FacKD5Wm/xFFFS5r9RDMKgN7tWPrIW8aW5QDV8dTvm21mGTlZT5CkJiRU
c2LSR35/S3XtfXOaZRi/46ft/UHR47V5lCOWPcwNPEx5rYF7H4Z6/KzR8OZfxZ+n3EjqfotOa5e5
PZ4xkwsZTMwfZ0wkF7Nsh/PfPjM4kAFVaiFyP6wsuwKUnmZKaZdpzODOAiGejCrzrbY4r4uzjyJb
74y7rMF6j4fXRsPkX2ZNA8Kf6HwJ7zZNGP9ZPiP2BClLc69YIbqDJT9on83iR9ltVVPJjIOW7wuh
J5RF4r/RJe5bppFEApmRnBSnU/DiL46Vh/NVLJbbDypIvllrZDMn8zAXMuUy1pTKbRCNztAnM9Pj
kSkn7VSzCJvdSztYs6A6Djz79GaQD4uVbzhT8iisrDiNb8g9Jka68IG9geW67TdotzWnqeID2jSN
8Ps7TGEYDfnptxlv+MfEK4MZdk4g0OKB8LrYI2OIGCMlzlbd3k0irOMQCua6CYUQJq0DgG/gHgen
ZxORCctQEl8hBUsy+FISX6VNUU8k2Zcpnpdl9DP/C3UU5iciARm76vWl1vg68in4jKCZTJyRPD8/
grPHy/isEY0ZoqD4alWbV1MZup7XE3LZb+VTr3jALwykxf8y/gnQKXpA38dQ0NFnjyhIqQxPfQNZ
ow2JeivMe0p0a/wtTTCF42qGRinAF9W9pzb0G/YTvdCCi0xz4zQ9fQHCJXRzQOOpLvT+ySAk8of/
1OmK6u7cWFD9Tgulrad16ovuvkyBypJNdYFPJSXTpxijFqXI/BNBpeIJsjxGgGG0xdTOLQxTlTZT
X0hEYP0dkXdiYyNkrv/9Fp36u4kgruhZa+4mhArRXuyKSvPie0LfF0RCvISYZ2M3DeB/alCSrR/T
G4Ki1QTXJBwq06YRQ4OR3Gk0S+rgn10SByKvq5TVTd5aQ6ndNwLJfUF+ay2PfNzF2rVQanAcouqE
WZnx50Um960wrV4n4Ktzpj5bxAyhSY6LgjePWjtK6id0MyIbw7O63jntX9kwIppZJ3fx62VNXOUl
3YLyIA4MkgcTDhicU1A4suB8lcl7m0Nig2e/bk7Z978OdUQ0XxLxydEFZBQU447m9h/25OgARIfg
FPtULSoK8bMTEi8Sn01hFXjX+mq1kM1Bg4q7Ah7r16c75n0RJjJs5pBA4SKtO0FdIcS3yh4bixMo
EYDOaKeI1JYvv/46MbaB0Q5QocN0CGLmfohsJ04rHjTXcGaCa4O7/jPr0KbyVBsvysfvOIC6JJMY
DvnQwDGftQbbQDUjJ7qypeEn7RecNYoE59H3KGtieIXNr9hrGNhmWp3jGwg5PevWo6WagpKErgHk
HOj1Yidl8JOJ+Rf7nNX8cVmUQWRFutBTvNVYLOkU6kmWBH/6v+0Zdh7vPguYdLgidw5A9/ZrM9si
WDkW/VheWPdkUp4+uld+RiN6u6HernqrRTl5WLrcoIn+fDaJn8j+63GnZOhYk5Lk4r5oBkBAZ6D3
HnZt8XOuHiowmNgXHtTR1OtuDZkpLrOorgWTEELlZzwgB/kFO9XvtxCDMrpGBZg6qZTqaRdYPkSk
/kJLmpQWtjwAUdZNpvUkCxs6CKKaUt+IMZwtOPzDBnbZqSow5S0VilP2ZovTPY2cby04KTqNk4Bp
soC+VF2kG4hGarHkkml8Kek7tOL+9MTim71oS24vItqDkvBG8/AlRuJI6DYDgif7cuG0qze3KvS5
hagAvRzkGeiQBttCP7hSr4IEY3Q9qm04qgPsoCPSc5CAHBBvf3E/nezXWwwEWLLGveOs1FA4LirY
6bdPkx155ePNzbDYSl1j5AY2kldm8azCGy37g2cs2U6cpUCM/UZlCFQoPi9hWc8FIg9ppTc1D0mK
hN4K+Ax9kwarpvI5M+T6taaTPaSlZpmTW7/tq0ePPMggVvhs+s8AstvL6QApbO1cFjynzOYiTBR4
UbuWCTc2xU7DioPADqHIrM/GlLzOSMdiGeTCf4zsQ8H6iVoXQMVoLt8NhI1gGRACd+TmN4byy9j1
rOgBb53tgaDb5Ik6d1yDIs1Z+IFXJ3eKQa/hwNosKnGhB4fakWBLff7g9uTF3id930NM1ps9+XXE
D/P01cgCf2ccrTlCYw5jIDRkInWzbncC7ifPqHgb403c8i1lEyP9XE8s4qwM89RAgFOE7mNZ199X
pH+Sfn3uC2ad33FoTfIPJTylBi91pjpuPu9NJRqE6UJEfpgY2GpY/ivXQGCW1IpaoSf1rtN2DlsN
NuyCQ7QZgCpN8e97KWcOXaw1pHGXrcIL9kt3BpI/Jb8Ku7guXVfIcJ5lOgYtgjRpPI3duS/PN38B
GTT32Ti/mApH1GxbeT6e4HyMYS2+T211cvPPcR5HiukcNqh+4x4UWOZ1JQfVk6XlAAy1DmzTAZp1
TZjd3hQUtKTDgRzUcsqbn25MLyEcd7dEiXEgVSYJyJ6Vt/YS5Xf8FUMkVBsw3k6Hvm91QdAIGwsC
Wt/iPAmINZIwWBBOjLNjJYIymz+kVOOrPl7CnsSJmw2itfIXpJSNRgNILB+akNASHRrbIYilRyGm
MLvC1mrh++pPChnxkRK77E6lrSpz34VhLEsjBbv+0EimLT3LyVpfWSs+AjXF3o8XMFpvZCp0Fhp0
CdPFvnTfbDH+McW8d4rYj+GEYCuKG4MERMDstcQ90I1VUjJhjGMavCl7NY6A4vaPIY6AN+Ts9gB9
lHkc6150eVXLtBKxowXeEukY1d9hR5QFjaBSMSvu5yhciEz6eDrip2k8NC/prMnnD8am14PYUKZb
qaq0to7TpB7/47DrFgidiH+hmwZunQzxadJVEsTE9SaX+KTfltzdac4z5BF7U0FuxrSGcCbaRJOG
LDmIt3z3d2pAXMXTGk2J177N68HCQWlkaekrOq85xz7oaT6IrBYEWHd0RTb+By+iUG0RyI3T+SoW
1HREeFnBsv5pe59dVgYqT8YGX2SITmKBfPfj5avvANkXdfcScJkuYJyfrHZdmo4tqFLCDfVOq42Q
4xdceqMbZlFMui2xvBOc3ZDbTvaZuzeNM0AozoImt52hEgDTSjiTNBNi6ujBgmdz86B3R/rMFH8P
wO8+Fz2T1+GaB4VEb2njm/2HkdU0PN84QPien45K1Y5ZO9xdFXqtf/U6+nka3tz1cF26/8gl3E3s
2Pvt5UZ6xk2t/xQG+S4Ok+BiapbQQGovqMvNRWUBRxi4qqOyetWMBhJdtZ3feHIo1fpa/0rm380D
PZ2AOP2qs80uJiU6GIj4DrCxmOeH72hnrBbe1GykW7ZdwqhN9bbAqlX0u+oApi+cPNJ4x/XdE22l
u/kLXAloSYio9LJEbwNtx6m+aJx14fSIEUAF2xz1v+5fBbWsHBFIxMLhfWZ3xoNNCdcI8PCk0saY
fbyCPYyDmeVZs365DaLd21V7sAh8WIafgoc2JJwWUCneTCF+B1ccS4ErRrogZGkO4zuzIkP9+H0U
A1dCmqp7tni6eXRicNWyROf4+ROLZFgGSZiuve3nO8eSrlKpMobZ5I7sRD+YXxc5w8nxBcLxSwjY
Yu5hjl1j4eUU0YAZH0AOPk7qP34oI0NSFJMZV3yRNhzGVNKn2qfcPoT7CjhoO9TjQ7alnLmd0G6U
BoNcq4n6DARBpvH8lqe5RdfshpR1tdCaEnk33y2UhDKyBSBCnYWbKSP9DMqE/XE1nhATGmXA0Qoa
xhs/SngzH0TwqaE+SUKylfFTvkLiquphmXOVXObolelB6YViykpIrKDqfqlYFwSxPl0UhAvnHlyi
XlDGGruqFRXjMdcnkDUf+yKc6sz7Kd0qb9Z8G+ZyqkqqibSnL7xK6A61kPI9ToIy8qQjrzv0OAbb
a3Mgce23cktx8x8oMFk4e6liyxD5dPl9EhK/EEHZMJ6mYccoy9PlYTy7/euonzgdDfB0SSNFHmxn
gFqTbq/BCU8DYlctcsosdl8DA6VTTgfYAw498t10ugPxUUbD3xOT6PIu746bHkiWlgWgwCu5/KYr
iQG8rL7L/YS5vMrqqULB+L6NEL96oESfCUSCd1It7/t2xgS8MFRfeDwmmSnjwwkyvv5KF32H20pC
0pVevHZW88EiDcnyIrPjCmdkuVmsiOsA8U/JBRp6jUhXvU5S9XKxKd6PEDMq1ffnk59gcvKt/j3N
fYnXUwEeXg92w4xuojyEmq6Zw36pTcGLTqEK0k8shjveKbAF3GJ8ok2qUzWFbOvq8RQAtWlyi6mZ
/0jFeEGqBx9+7JILZsa8nMrD4yCK2Jriek5pYTflGrPXHTQJq9IzSUIR1f6bpKOU6gl6Jxv2iV2S
M86K9OGalCH7CZis/Lp12LncAPaFhtdb7XP8y6eBsvUFTt98rvvObaREe6BVgFueIaltZRWm5sjD
v8E18MXXUCFzI7Z/IYF+Zp36ko3tnCCZRSUESuQhDg/KE6O5JW8zyyRWkGez6ersIW1VoNU0sYD6
tQlzG/FVL1oEFumNjMVXO9ZHkhG4Vc8f4uNbyQv7M0J06kGmSaRg3+k1ZhCD58K+iociMVxfxMg7
NXRww2OmLHxlDltyouq1vSMFOiHHJqMdC1hksODcxjdPkmAiaZc+dBC2t0GER2Bqh3CWoub/ULtn
ADMghxRU+joIp7yWNfFXCjI01hlD7LVCYWREZtAEjAsa6J+MbQDR9Vz/Rg7rfFjqyQ13hw3+4UTH
kO0ulmrqlnFJoQ1pSsgNP+QlJRgW05p/jvB1x4uhKUcsMNNUkBoZ4Rc4pNmopbjAUuNQ+/iC3hwX
w05dIm6hf0phdUy57z3Y7uRa1S5PQNDmq4i00ALQD/bUYG86IHeUQRNtu1+OJzYgTvgr/WhhRpS8
nxh7jfGE6awsI7zGGc3n1ltuyrDK5LIFXc5pbMVlJqrTrtOv8HJGOfNeF7wWkUt7VarIrOwO0gSY
MhWqRbFBwlanpQVfqpz29qt6LmFcJNFhGSQhMFC6G0Oul+IuUxNmA1Ov+7efBHWNrQpOAo4faIqA
kc9giReOZ4rwiS8vg6TLRWVNPNam/GO5fAIqkTO6616XHVn7zVc0EuIwGWtVq3IFF7M+8+AUt/ib
6qGx5ipFBaZxeE9x6DBfw1H8HSYHsEH+vWXAhrQrZiYbWf9qMtq8FQmFJv/9fWRQoXcE6l/yX/54
ZE5Vai3UC0kMzHZvnKot2nWxKR85fe87uAE2nUtoYdAJmh1rjcIov30ojtWykvhveyYK5feQiQs9
a+ACLtXvi8sGg0+tlbuNYt9+TKrEYNK/E/4Eazmm2GtU1EFB7rI232TOYzLufoe9Q0sCo6diGuRb
HNSFOZDxLKNmtpIxHuUw71v27Jjx2Y1+/lOBP9J4EIqTHPz8z6BL+sJfzHtll3SOS2pUZOCzW7EM
I6mWPzZ10pneTdOLy9VynpEFLmix2QXV6vPoUL5PaBoBCRoUZQHGzhuzh/U/bo7RvtuuWAIUQeiS
ydGH4NPImMnvIF5hXZDZ8H5hRhPfBfp7zj5wODjgkmJJX52lTHtbfyK18Yz6by1GWPKVzlrsSSMo
ftsGLgrpKscmR2eYiwawmNZ+E6dDXDIKhkFDLcnzpVjkO5ObV4zJymcMFe8EvZoL/4bPn1Jbzz4b
tkHtPggNbJwJtQsHzn+QsPKH+4SmjNQWMCLWGT64qq91RQM2Ix8mlOuh33K/Knn4Vf8jqyoBXCfS
41YzZm0jG2E7IB9BT/5GRetjjgexZCmv8atWumjI6fUE0PwXS8rYtyv4zrvhnG9PU6UZKZpNyla1
hcO1Zy486PE9SHW+MzZYIWJZg//YW5pxzsrqGbAmmLmcBSJ0k+UieWmHTE8NQJMofFPnv/DyAluw
16eved32Euj2CV+q5CT71m0Opb5Cj61QqOYEuTcmgPUSWRCZ5DLjT+rJYyIFaZshG2ntZ4hduxyh
zCQ3jh2RKVj79C9BsUTwt/XCw9jnmxv35R6Gn9TLuOqigqJWbpiqxHN/sm6vOxSJNFUDx3cjHPdX
C30afkZR4Kyd8tgrpflGdqEyMo1oi0x6WtDxZEmF17J7kme2F7dk4BrCnDZHSv5419ZKvPIWUZfj
wcyTI+9IlNV/n81KqIcLf8tjFgV6yRC4OyLsUvYN697n6bqJzFaUg9XkFY+BJ9CW7Al3PXSYwtg8
oWmvoHcPAkvdJxXFjoIhQyogJ8rPzaxqD9NLVTB6TO+3a0B5yb4T9z8Ll3WIHIQ+7SFCnRALrMWg
/sYmtW/wXQk0qXmtUSO9yYqijI2D2PojFCtd6U4IvSDriXWeCHQck/JWiZYYGC24wJVyW32gTbWD
IH0ywDOZUERZb83mXJjXent05EFnwmG1+4EQGmBp9pdTRDpUxIVoH2vTX6M+4v5CtSUEWgI5tVHH
aVapwlF1I3FGsL06QnUaEnHk1fLbyF0riE0mr/9A0cV2Z4YiPiYAhpJkWntVTwwZjsAYdMxpEcTF
y2Zs4SzpPgTxoBGjkKJGI9guPgfd7YUTzi2Le3xpWK5KModjYBs891F/Wjr3hu4uGPaU99AKEyHU
cPcsArfZnRFx0sFKQPLLTCA7VW1h7fx+6skCTOCXuCI4GroTW6EgP2TWv/S3bs3/1YXm7rsiYWpl
yIOk8Juk73m14wBLeDbcbAJF7TuaqGz9Vk7c993Kqj8r9aoon/2PKNPl/CnIoDmeyTrCV26e17zj
TZq4EUfkbFL0vHUd5lbusCHzMqZ7YJtC01bwSq1q6/oAu7Nu4W1w1VCJdXPGobTOtQ8wAsPH68mR
wPiXiWe2aeK4WFSMECX7urEFHgY7ITcgeIsqbnMVHo99EOuLfpBWgD5opJ8pV+pqqZgOxklHxrNz
9lF2DBSpDyUhMlnqkwwfVoACWGJtVR4YNKCaWB/bgyLaDNJqd+OUQ6/B4f7zGkF0yZ5fHPEnXttE
eqJAhYw+27Yd9I/dstN6eG3cFUoZl+lIUukhswXTRESoOfBnlBNT1ICNj1mtY4+1u6IEH/gEIP51
VOHagqzNKveWu4rPTRtWpRVcIw5KJVq+uBJEwM+lumrtDbe+AD3dadBiBjtyZcVBYB74BFT2ohJb
0pjSNvOMqPDfQn2SkaUfNPeGTzaqB9EZBp3XvtcxKpGpH9o7v7wHmQXwtbJ8huaq7yx9ViJcH+cU
wMnRgsr6xub7I2pGm/N+LByI041sGEFgPgoE3MqAqsLHFHvOUHpvh6PJEo2TR9iokRUAsPq4jm19
Ofjl50YOrR2iY2cyih9hnGi6+J+qC8xJh5t/OwzHfQqPW3phUXZOOwm5BbarL2TWMVpoR/+qwc0P
UvkU0MOzt2t5IZaus2fSbW0TF37RCJYBFAzTEAF3ew8+eniD1MP0BbY7NLO+lZBTjkYJOAWuwIsk
R+VzWYu60FpnYAb1TTEY4TuU1TP31V6LBadrJkncCZUAvuPURAeHb0VrE0Pl+8ZfVIPhRMYXmash
rXJPOoJozuUcL/xMdJCK5BJAwqctkmYvBmCDy9jGd0pUhlEnp5bXgxkWIVvBstiUOXuKv6goaV+K
ZnrEcEjdJSM9vyxL8O/gI20EU0j1J9Hf6Pqfahzpq6JxRbwhtyCoWmmZ16DSYMQp/FxtVebD1XLx
xfT9/ut+tte6OZt8sL8M6g7LlVqe75bu/I61wbZ4HxC5vxUcSEbVuKyYWECw6KBa5BVmX8PpEPzM
hqBzKihedDlK96fCA7FzgT9IltFwEM8sdZ3Qngxuz5Y5Mr9kkLiqAbOe4vJMhQCzPsqoy8fPMY6U
q8kc0jW5nd6e9B3dBlB/55MMOREkDndB7Z7bwmcVVxFt+YQrdApAaZMpZ+xSxRxc0Nd3Wcxmy91r
nQ+Qh7vjMBlRLqbOAnjrYbawT+dtjlwGvd15k9awXhzFKU90bmWZRSIVfVH6stT3Pp8NxXYGxezA
39t9lgV3NpOZz6n7FTDh0Clx0qmwwDWUcde30RVtboqWob5IC3CZeeL984NOQC61xoa4KvcbYsPv
oRAwzM0FTNhKlXJ+IjMZI21DYoJ+IwUsQPbh+0/Fx6Ba++qjq/SGasreWbnQAAazkc3R+T8niYYG
GQFPnmoocBsmTwFWEy1XRxBCHv5vWdcxCIW5309BLRV0ykefdqT4AL9DTN416d/RuhzREcPZZ94T
+yTvaZzlu4fmG4iwFs53275OWL0DH0P9m6g9cTsT/A24fdwySDjiS7jBSpvlogGKGU9sh4BN4JTC
Nrz20hVKdDKAk/IwkmZ2qJ2EG2+EsFQ7xxi0JFYSbTVWGqek5FQSic/EXhGl7w4gMHVQVc0XiqMX
0Euv2X7oi0fXxcQphbad35s4v3axEzoNmxAb/YdAk1UegpMe5ucn+aA6NxL9DwArZchrmuxbgPoL
7DSm9/rzYjA4OIR7IE2ndheFP5tsb4ezT8rklA/XDSnwyP9vAuTgD7cKUCzBVHkW/KXzI/gVQR0f
M8zZTyQ5Qq5O6mjybbrHb1owafARZONZ/gvYS+GnvSYGocGFzRrc22/nyIMTwQhVINZkbc86i+Lp
88BiDxVMN7yrEsI+wrIB0nF2Knipz2N0FHJt9Nv0HT0/zfPFNXDlkwo5+TMedb4tZ3g6qDZ0RNmF
W+7swV+Zf5QjjgXQhn/+dURO9N/YpoAdAjAPA/13honJ+Al8qTeb+/8rHACIk0ZVNbBH4rFV/ho8
Yi552VJ4TXuK+m/PhjUZFMIX/V/2KWKhfDAMR/UIP/6pL6PrEx32rbHsZLvnZwvyaqvCwA3/jA0/
P5c91SHUgB8oo/BURwD72pY580LpYSzbZnjYUiRSbbiqdDfrt3qq+Spu5niA3SW/SDM5KSdkhMsg
rRQ4O9dihcOgtpps/ydogxP+FuY5xQWH+cGWzmUxbfb7ZkXD62Ew9C0ILPriS3HuPtTl4EcQgCAv
4b7cQNeQ1Ng1c9nDbrBeLPQdt5/uXM4H4jk5KrQeYS/MCfvSqgtnFp9GirR5cBMkHQTBwW/Z9aiM
L8FF2TrVKCJoHqll2YH0TQp8VY+EUnIOjoNLX+iWaSf9nRAIvDVF26lPDpqCQv38JVlzD7U6M56T
hVui71751HWvqu3g02VnhWNk6EnlXYN3wSjV9ldOOs43YL2Qce8HLFX8++o7hAzLHk6UfAPfvHwI
XVFcXXOuSzqtkKqCiJmt8AkKJv2U4ZoNj7B2r8CyONP3PUnm/DtuVkJ6v+7rqP8ZexUKf9oAdmZZ
cNNha12+y4on6IqMYRDDWeSWO3vME7PxwwgXl/mO2IiUPcCTqeWcEPO6ts/ttIXybCO++ANpo+nC
ZEOqEHvu0wWNif2zHAo0NuhUDYevvEnXxcl1sPTKQi+RYhPmrcdcVczn2e3oY28BDcLIIWdT4iK/
LD5AnVz+KBijK4Xt7ZJxDld8pMItb7iJUNvcv9IhnP9+K90QpU0y6+/4EwDE+Odi65iTs9SLIvGy
i1J5BDz74zkWH+taCWsl4GCGrxVOaOrqU/YbPLUAtM1U9XJF49/vS8bofcAqBpETpbhrOjBw1ZPn
4RksNw0F7womdvlyhpq+8fNVSbLvDKfXO4C46kCVAevZ5Xz2Rb3ru1S94wiVhKNSfwg2RyWJ5dYt
nTMKDRAf6+nCYG/LOJ7Tbt+gWv4AZLk2GOpvLNu/2wJz0pc8FguOMmxUaGgbGGI7ZelxcI11Lxvv
AAAR8QEw0pn5OqlQOG9ewX0RVQLXvf8mnKuBcisBSWr7kaTUi4BlsY07ze046D1Y0lkLTH1LOnsN
F7DMxpexlf/Pflp0wud0n9YVwWipTpjfxdP9qg9rCOvbQ0r//Zcs5/X1dVOH9pusF0COlR766tMI
5FMaWUXssGdcsFdlTuTfHZMmFdITpSVf2Kbo7sZRy745ajrdhjMWCU2Eq4DTJmc0myB8+dCIYx5w
uzbxuaFygKb71faRBUFCQo/R8FwvBnOJ58DT22ibqqmeVzbR0WcUJLH/zLqqq6A8I3bji+vU7rHR
8GqdzCnpMcdhJYqrOXQuLcaPPXhVEV0G2mE8xb1UFOu1/g+2G9qMNC4aIZqGq1rPEofj9assFljf
RJm6ER1Z0lMqFwNFOowdWq3lPpwhFTcADjQyZdYEJ6cTrBoW6KZEc7y06fsMq1JQYf3TL/uDakCD
1297qdAGVD6n8czTEz9hzoRlhlOUStiaCbw137Ce6GLac3tty2qE0x8G8xHCscUpxmxx5RvPsf/y
TlWZ9YfAzHTzp8g15td2gT9HCD3MYjXYTL5fmjg0FyfKL38kwF7Q1sYah7JpSBEzuzIm6KlYeymp
S6iajXLYskQQQZ+x86LhnOEArddEx8O901pbPLzjH2CKxN/ENT7Su6HFxEPnW48CO519Jbzdvi/+
BNLFz5qCKUoXKlPYOOLjr9GgN0rIqSvYfZxZ4GL3yLi+LxppWYJu66Tp6x9ZhXSpps5guZ0JNZ16
dJ84jE93oo97B4TKr/OCUhgYGXPwqp3z5OP1mn/ODpkjp9TGFXE+msN5gDsSB4Wp4OiP1ZneCjrH
vrMWcy+Ff/gfMR+6nWUyE6NK1mrJ7hlY/Xin0B/I2/sFWcazJzzbF5ZnTbKTsmUwfAOgtifJkNX1
BPEgwNwkVDpzYYlNKCnmGLpRs4P3deY8wfLEJAehhK2A57u3kQyNmZXOxG1CmUlGHOKZuZj7USi4
hun4A7qUobCjWywDvqE38oevb0f4N3yYd4oxyY11HgmSM56J+UrgoAd2TLj1SkNr62hT15mxmH/8
UVnGeo89XZBRh8deJ9HT1rx1/t9wmXvvVdMlGJcpVV7ytn91y1CDykI3cK0ZWXPbhZDquEH5p564
TMAmuTGfRlwTz2G5/Vdt83YQ+CVFm9Vr7kv9uzarInWvvixAsAkPD1aTSv1+xo0xfFc1TDJKJ2SC
eGWVYXFo4JLjujPPozyuM4/3h7OVuyIZEQ6C5mqdHI6OGCuKpJ0dgfZvXEN4QewYD2hwO8Er78ZS
55F0Y0fc5BgJFF5ZIED4yvcGWc3MIT2oB3+l0cX4tsugAULvLWONXe0/CGRJVJFl0gh8sY1qpk2B
W2Rt9XGDEVJh9FdE/QPCsxZMbxWrNGrvwJyQCi6M9krmZsyTeIhZ8jhZ6rGtSnKeh0T/tQtnoicd
HC/62SqmXq8gUm49uN1tbpjba1ywyfBaLAMYknYgozfNRBz2F6VeTz0BeOhHzR7HsJg+lYjECQiJ
Y9hwa2hFaX5fkXOR30Qelxw/EE0EgDQ4hqOov0/Q7oa+ubYCpyb84BYVDIIZnVLx3UpbBasTp3pT
wR38cr6cWWBr+UhfGeHUylNB9ILgIAYLqFM55hfa5nRgppyoDL0SU0icoDrnOcWsbXeCvx7OX+Tv
I8ZrM/OJ96hl4vL+Km5E9ceMg722N29PmUS2GCpr4Qhg44W4DdDcnmzNzPCSVpX9WhYvIJdhf8CC
3fetUfpn+GK3T1+uH63r8EfCiJkNjfcMg+EItWCbqFFl0uVI7A5uYeeoU9elbH4bfXzKJKfHrzxt
C6Jb16/XRfrIviRKJuybxwk1T21lSaCC+BaHuwcnNh20wLRiwmjZg6nmjY6QRucDnh7XXYeHcPey
tHtPKn6l3xI4CUaGT6+vj5vjYEth+k8UvktWa6oUYMOEuYox9jkdlxzNpjc5zSoD2TCAW2GI1V7x
53lxRUJfy/scF+Ss9L/sK0JheASPDKk7ZIE3lG2m3MjAWLFeoNYlMKUnMkoU8J/Vid1TyJYEvnlE
cWiXdNkyCy9nGI4LKQuH2geblriRigoxViXhrcPvAOleaMShh17So/4/3cxZesfmEe5CFCNFOWMJ
mpuBOsS9+9Lgfn3jxF4xB6hE+YaCpimEnyQp4STyO6CB3gox3qyI790xVrbKSe0Sf27ZAPh3rvyu
yoV94dvbmlAF8Dr40LNYf+scnCQsDMiErnHEeiZduDDg3K/sKSOjEbs2voNhHQrJ0kX3rwVC1TB8
EZhDeVR6ZTV3pHHo2mFn4pBj2oXAcHwh4ch1339akkM3QSi6uf/2lyt6NNlOPTwZ8RUifC26cloi
HrSfHWDtuFTtQVfHuDU+0g7/WYWQh+etH/lKJq8g+zYKXBQDqLNE6kXPYC25eCAbyYzqCaeYWhEk
EzkxUqQGrLSjZYFXaUMh78z9mVipu2sIRfiuiEf6jx+ntnapfJcxippFlJfj8xklZ+OZOernFr0B
ZPiMRd0rqVT9Yhsf0+mmERroUh1KzBMoNnr80ILkFy6Wt2FQQbE7QiI7QXE5E0oW0ttqtlpyxDHm
9tP/hXCGaI2ySsxpEjKSOHMgkxqpWBeHNGYktvC7w9kF9062ZR3rvIazvDtKw/i+WYqpI5+7Aonf
5eJoqyl/Wg7X8Ys72U9G3/3nNuRDXM29ao/08G1UzGxZi16G29+A5Z729V6w22Mvu2zAEQj9BEla
L3W3uVfddkYPeyZ9BiSs61a9IHsX+mKTNlQqZLuO0Fn/6aa721RY1oprxgHE8i3h5+l/ehN0yPPH
mVhxWL4yiAK/sc56ay8uFWjDpaXrZnvuKxkNuNOrwRmQBZZW1To3LgVB2DaJAAjsTygvUzAEgEwL
+Oe0s6yeeFPwjhSNE1HTWWnBYWkzLbnVf2nRxUnFjJEIOIKI9weF7uRaoFrIZQG54JJudV8VPqSQ
CVIntPJy7HfnsYp74i4mh8V8+PDILSEeQfcohvLqMTKAllQj+gjFzYqle/p6iFn1QaUJks9s6pPY
uLVK2U8RM2UO00nxPNm82JT3SgBdFqTMoEC8/fgzyIH2Cs7Ls8pD52iDoVpfPywaCCZkldE1hNtH
+w8zLeh686EaOIHRQfRSL2OoZ2kaoHeR40dsT8b5Yg6egjmabhxktfqxWhZqy6Lh6xfV+kpfK7kb
J6f3q4kg376XlAJd45rUxY38h/F7PmXgO52EPIqCsLHVhaSZ5zDbTHd/4e9jGHnDWJXuI+i40kFx
IeJx62k9MHtT22NmdisvpNz2i1ZlnRB+6UlvOLvSc/fHhSIcLdzWXSzapvr6x5ICKtOs/z9rsZng
fll10Vg759283vxYNck9gqdUw6SjS7kcjDFhqU7ap+JIeoelV7qJoYq2MjaDvJCXjaAYWkplN2Jb
6gBqo4opgFHtRw6lWiy+rmWW+PvUWreKcXjFC3SMGthlBji+WV/+sNar+5OsFyGst7AjKlFCCcYW
dmbJ1WuEG23kzTcvpWRT+OKlxSMZvR9H4TOu+glcX/HYeMsQIEc5T4UIiwzo297MiqsJtCHErB6S
C3K+4Z6SzzK6DeyxjK52BzmHhkQE4lBpsl52GRrMXHSAK0wSosrG1akYdKC+mU9wnAtLeXT51rRd
nTph8iQCYpjeXdBHlChAC7SyQ/b8s9ZCNSaR8yHTMSXlr2qtwVN/I/Xg5M4yKas7uEZCQl/ysUg3
z4Qmo/D+oufoguCGNjGFRz6TXmfqxZ6pn9S5RIHm9zY75Dkg/C6nJZvzUhtEZw7MKhE+l+2W9YiS
0v731qVjqMQ3v0mu7m9bMWdRDeO6rOrAuuikCz8cuiFsEobvqXxlGdq6b2z5BWYT7hvcGnr5H23K
3IofaB+Hoykv1O59Raz4NIcdHF9VhFoex9YYz448SB4R1VvK/wnSWUHSUNGXPe1me9iIhWVYl/zP
Pl2sXOEQNkFubCoZifqDNXJvkWVlWhA6UXTTLnTD71P7C8qKm+nZl9757mMv1wuf+4LPbJSEVFd+
lYJkYuiJXT4afaU7bh1Ryr2NeiPvYTIHB8+WKT/Ngkqw1lfMZ5IeUUzswyyEjtkyVcaZvzvVy9Qr
/x8vPaEgeRFFcMFj4YQ+0nJNLoqpY09QBht0N+QQW+EtzH4mqWVtm4RwSdDVQvPAsrp1r9aAHYxp
iK6hp61/NK58LzdC8ug4syUHXGK02ZFDhExsc0JEUlYhhBdAyCVBzy78Fz2b+LYWg7ltGCvfgpfn
KIiBeuXGKIqDhZw9DZuxteaRb4Q2hwh11YqYbpLORY/jBUSBQ2uQo+ld6S4G5hF1TzLpESCeXP2t
NQ00gRehhUAamVy0O6Upyq6ZOH9sNiLLzOLTEw1u0881eQtEmTqWAez5AOPhvN+LAmEWAjvYJDer
gn6TO/1fs0WV544NbBN4ceqyg9LLC/41XXWO7K3A/f4aGYd7xlKiD4Sb6OiR9fdSqFkriJ9vj2Bb
87Qa8DkLdtC2Cnrh2K5zpLqmnHv+8y/z84ddFayT0OtApnNuj7gzOX2zkKadsH+mEozjN5K3CDBT
5l1QFdg3jKnsn0HZWq6PgPIv0SlrLb/mkJAyhzVF2HZXs7l4xtP0C5wuZlUHHYJJIDmn8iua5yDK
vZTCsSzWlphwGW9sgHyVTazA73+i8zC5nQbIhg7ZZ/unbDwERYrw51TZQxbohLT9MIjr1m3cHWNo
BSg+pU1PyrSTYbqYstmqqI9TZYMMpJ5Plsq7FCEEZv7Cb51+AgtmFhXQ1mFTE7aZhkIvtBlH7Uth
jW/BJfF/yZTv0W/Zay77OOIHSCDbCMYwgLoqWPkcXxo/v/8PgGrIbSy1m3AHGPcgn7PmgyjdpjuN
9URJetSFyFicBpaGl/7CCEpkFe7lzFIk5x1gIwg8SFsMte6xTfrK/V173sU3ffporRtWZnBSvydF
fLzMzSnhV60p45rHee6feNEgzaOlLYs0xARAqVXkHkokFLL5HZgp32FJNZlZsjzwp0i7AFvyAIY7
5ZhtbPi4Sk+Axnyb0AKkl83yE60UFaJ8xKo3aUZajjF6P8Ip0XcOHr04y3mSTzdxZm+EK8bvG80k
ZgGrbQX45mR7xuxma5OYKX24aAEKClauZqP1txxHh4cyjsLGqg4vwrxwRMS23zJ7KdiVrv9i4YYG
H8M7wQ7IDAwV9cXixrGnB0vqGTmoCujAowr4GpBtRKKzkTRhiiQ+XEtoIQ5orXSTX5tjAhgPkXLJ
jDqo9BWXSoo+NSl4mSt8xh+rOdcMqJ3Y2ehMEw7oq2vVTuk5jtQ+nc4YVzqWKb0/joM2RijSYPzK
vo65a32WoAh2cYziel8KbSClRWQABCUYZX7Wa0z5AmvAKjpvCJXch3GwU19otatu+/bFGj1ilVTF
7vC7aEwIgTRnEdHjyFOYcu/tvmX3IhPsZZnjU8DSYjyGW6qziBmFynyUMfDe5ZMUZppRMDmukHuW
MjueomoARUP4HTiOZb/knDEvmLmu095/pETZSTctQX9PGcfAuugdL2n97xHjqmQX26Q1LrBBNAcy
FBQscchpySMpxyJ3QVFPb5SjcxJnHbdLZy5FgsGv46Cq332UcxTD5WSOYOgaEym5hZMiJJgKMcDg
zQBBdJuIc1U2y4d8xtSZtpusoFYU9/BSb7Z2w4vjsTbX+QRV4aIkRJetNQjpfBOdFcA39VbD/5Yh
+nqbcULvOqZP6RQ4sTMnyY0jPG1lfHtPfgYfRwxBryQ9gU//7zoceTsplWMcobZN80KesvToHO8H
Q105TSUfT+ZbEQTtIZEHGFUaICUv0OUr1iUUBm+w2rasqSpo8zr60cTd8SYASjtRs3YlhTClREhW
gN0hqazGLFKlpJkbonVWrXFM3k5XDqulWs3puZ5Ehv8Bhash97GpzTWqJunmX6ecOUzsJVmixzVg
eIB4zzX7OPs342qMLkIwJbFXK7QPB8KbSzayvmqI1KpipO7o3K2rTY3lK0rcVWMNbf9A83KXJPZy
v/zkbxqoL626vADKUI2heXe4VA+PEZwOdU4iLoboZHSpIWh5rAaK4xfACpgYB8TzYr/XDT53oU5s
+ZeDnqQLQp/Nu2+sWqKNBPiKR7xPzX3JLgKbuuMSLdsOy45W9q7IskTfOMCc8fXyaCty4tSM38mR
Xe0jaNdMYxuajzWC+JqCs94gf9O9fO8upjuUlWJZswhd3ekCqoxNcYUjzezzKvz4N2tdNfcN3lRk
mKgXbX5ZcfoyOyI5lYm4LrOIU833W2ri//IOS5xtHr2UzMO95nY1f71BKV8/hAUYERtZIYU3N+D6
q1CzD0qJ7W/mBYMdOQpQfNCfldAkIcfqykthjQKUfPpA7qzcuIgSiAWQx63PIWxOPRKSLgNrjpf+
iFUBXYVsbQPYm4dEGJ3K2w2vHViGZrG6/cbUaGVpudvwDI7W+l7V6z/k47HSn7hcP3R0He0uqETP
s43V2N/ZDY77OlwgwOgsPVzuknrrvePkxbQRL9nIYuDqTWxe6eMSO5kWam65vWDUuigqEVgkCs+3
VNUnafs+qiDh9PZIINITMHkXmBL2acqvFA/cPmqru+RFy0YoZsWi2Xu4KmljFwqKtiQxeZbHM0F+
x5DBH5mjdRMabLMqkxrflpvgsc5RS0JVHk5ABaw65z155OZVkfy7QMudqKt1kjl6tNS3LzwsHZcU
GjOhxZXxCN/Xzfq4rVQNsv4fbII8sRxg8TwDXFn5g70X00To1jm/WBhrgFoDDccNNHvTAqd64BlW
JjIA6avHvsYGvfWMDe1g6cSMLm53wczqTZG0+CRPkQRVChnImoKiTazsBm7emzLEiKrInVyKLs1D
G9QkmkQFP7s7sj83W98Nc7iBnNrPeWTM0N/nv8FZyXUHiaxcAxcU8HXN9f53QHVjHiC6BfLRcjev
bRpl9vIIn3jbxdygo/IqtC7Kp42cku6KygIJ6MKWOoQTgcC84humM2gbdM52fYElUCqoFZgpFKzs
O5xT9/MRkwJRzs6q9f0v83c4Cpse++VTol4/wH1z9BqWdWJZAq7nmV1iWr+sgDmMbTB7wDQoxgbQ
6HSo5btkt/ZMUdXbHljclcbGWOXMEcH29XYzEo44Qp5IZgEYlS2VFJX4Cn6H0G0m1WlUstVu+Mdz
zrlMR5vL05bMCrI5UK+bBwz3Ax3b6+kaz8aQ9SSB9pcIt2vAuN/al+ymEKNNT555gbKxfzrjj89w
U3ViPlqyxuqsN4k7YBbMus4kumSzZxYCOMidIdg4yMKefCccOjH0vOvV4fUQHYd6RtvvVdRQxsqJ
wyV2sHgyWDJ7m/Oet02auw1MR3eMdwsdy8R338thd/TBd9ioVlQV05PlZtu5Gv6r/V9N0roYzUrg
rNNwzhYNqM8jtkc4ZOB9SBi+IS8Mcf8/S4fn8jAe6QgSPArvWF1z5NPANvk6bI9ID1P5zVTpijgp
WSqnZIsQNoIDQyjHI9R9n4yfPckO8KIrOlHydxDm4m7eecbGcc2y22KbuOTG0w7naYN5aJqOJdsX
nUuZZ3VWDO2kQGwYW7QozN1iqcKLdA+ugjZmDKEy2bGcNMxIyb6Nk2BquDl2AV0Ov7z6YOSHXv5Q
nnzwQywTcLfp7Gn6ZhYNhbz2x7l4+947kQKdwmkkoIvw0ubOgIiChCO44UgFfOObTBwY28GKSOzf
KElz6/mu4ZABi3VKX/qtrdQLxtkLlMdjOADQet+fn9Qhda1PVUBowP8jV7YW6NPzmTO+dCcbF5oQ
BAxIVZDeRrjLL8OY5xZJ4kYtYLEO8LIq48y52zhtLBykjAT7c3muftw6Gik88lpSzG1Qu0jA7O9m
ooozvyhWYhncXxU9EOncRy48pPzlk3iSXHYnWGXzDeRvXIvybXDAxxj59xjhw96BxJDmPP7JfUfY
+NzJf50CNs+LtikvOk1nuqyVPbGC5sSMDTJFutkKwjCZjws+wNgb1XGU322Yy6FI4Q2IkTnbhq8e
Jf26BRSANWtL1xUPLVneEfxyuAeF8pUDDwIXMVY8XA2FpX7aTrbq9lf/m13855nOcccg4F/xl4es
aOELoMc9WlEl6rCE2JCM3PyzQOLUV0sklgPTcQr1rYBbA3z5tvW5qMYT+yvatcFjHjxkuIfsyMrS
V8/onRQdYXfZPi7sR9beo779bUMfAPMoaf8vzRbApjMd3zzFpLBvIKhQZZ+ALV5snVOfYSfLea1d
jo6P5AmioFg2xgEFHh1EhxcXvLH4VKzsEj/OuZ8Vapp0USiibJEild9XKRaKL7VtFdYgCwrMAr3m
SvT0ia2wji/3wc/+84W5Rar4sjxqniHApRFKn/WHevlP+01tUXq67xAafAAMb4O3CxSav/xfKCob
T7bfRcjHWXnqMIkCNDkKMMdJ2Xmg7uvT1DvpKmWr+CBneGaPMKJbinxpw2siR70jrQ2VUIQCGAwn
G008Q+xkyYN8mEMY1I9xVIplNudIszRoo7dBSOF8EimmcP09TN7hPxqlg55ykcF3qnCctODoC1bi
tN3UPlnJ5IAmEKwg7Z6gQ2kYXMJc5yKbacgtGQnFirAB8rOJQTAJXQFA+Cr5ViLp2iFYRULGdisc
bd3sv/GE7JVIJ9mja2VEX1uKZJG+IsLhBo+tPh0/MZ8RRajcbg/bW6f0L9BAbzzxaN5gx2SsVVtP
69TzufoU2HoET+nBOhvjYxGZdbAf2m/Y3WKDEy9mSC0XpwlBK1ywPCs6NW2DnViygOep5PtpoUpR
4cX7yU7Wd1ynfTq02bh/oy1eFrmMCwoxKGwMkRxYcZagEACJbSHHnskOP6SBBpCndqdgO6TnqYUe
Z5tKZxjNElNB/dFLTAMWNKqfvW+Gj64mfbCvj0LMRZsTbES4LllQ3WepvhprnoN4NxwAtgGgqkCj
+KkGoMhWIMjdUwWm3GorUT+e48Fbab1I4DC9DMAgaPS6LqRk9qqlKySAHzsnUpME1jXSUpk5O+pb
hA3twbBFy+6ioij28E+577XTQ3eZU+KQsXcE441tsbpAX8KQrgxC27gffPft8TVf2tuivz2+Yxue
j6xpsC9Pusey6WxsME1E8hDd0CTIOT8wL58zJAoJrwE2pAeSYtXAzUcUnBzXZkarBDRLkEsICTMX
xYNJ+G9HIJZ4o8F+PZFuyxLB9lqxVrDJtrRYJYTFZnAsrJsEGWxFHlGIU8dxWOh0+wJXZuD/Vr7I
7UV6ZTsimhdCQwiykT9mxtbPjRMu7O1pslLdprTb4Dt1icnjlOcbBt9BjJUmYqNUlkfJLa7Ti+hd
Vy3v4WK8piXtb2yO1tX3+0+CkNii8KiLUxFIWeCiOBHYHAjLoFS++tPhg3kI7/CCOei48jpPOHIB
g32O0u+moL6j97Xt91AJg8+mFCJ5HuX1iDfm8VSS8pdJA2neZE8uuMgQqy7LXPR29+OfwvEMOT6g
VI2dlXsoQ4qOQBR53LyOm4vLr7Py1i7NvFRpaEBvSFLBWCAvBJVBeFBQ80zSVjD3E45S4isk0wpy
v5uxGrCAt9OYYjb7xYq8SDayT3elxPxVsOPkUZqKZhAOH8/8frsH8k0x2aDcklapX/xh9YPlsZTZ
CS+ORfv4mBAkpznwonAf84flrTylhLT0QeCV7o/6W4P6VvcZyDXxhaS4C5/DvT7g0Cl76M4cTcNF
IeVeQxQcXKoaoLVWZhkEwmz3bskcEFzo4wU8Ax1KXh7v91PfJ50Cxd7sIfSdUtDT3WAcOPjTbIfh
XksUtJlIS5JsorF6TVdP5ehREi0fScObfS/VYi+stVddXXRcg/iLdZyIPyaTJtEXd9QNcuF/Q9Yu
wyB6mydYTeK3sOJtm+F1wFIKck+cfXc2v4UL3lqJWlRKZaiXlunjgsqCCIMhUxmF2MZE10XL/vsz
KYgZ/lXvSKx3gF5evZEfG0Q1Vy9yOvFEdZHCtfu8T9bDFeNyS9D4M8wMYBDKD+G115lBwkmXQ/yQ
/qZfQTN2mGF6j4GIEIVnoznIVxJl0oYARFJTBYJ1xjDS4oR5p9GAu9zQk39X/fxhg/ePyEcUDS6t
c31mOvyAJ+BjaNJxS2qeZkuRrZHgI0nRoqVWHYDt5GcWn7lJUKYBdr/kOxPd3EP2PMpNfpAlQf6b
rOiPG8g2hGgZqg1B53bWmq70TbIpisEMoR6RV8UZvEN/HzWo085eb2gpuKwRdajmOjJ33ORPOMS+
L8UUq15wvccOhfrNXEld6z2hLfyE4sR9k7Lxz/R9JC6I3SjQW92daB2EMn51/snYcM23ICP1eNZd
zB0sj8PP/ihBwgxrfFb0QSPifnYtlKUA1vcNCV97DrIq0YVuYdT78LlAnBEhI6AF0GAy/wsySWcY
8efQmOfzllLC9gEhMOtvgO1+wiLFnsKdtmHubtS5roIpbq6S2WqfNHFLUAuBJLeyc+EsqeduvcN1
7a4MfMzdvgbLnoHa4+oQ8U0mezA+fvQ57VTuCen8Z4g+cPiVEjaXhHxQuTIHzdyFwjF2oLM75BSm
Xenho3F4fv0rmIjuzbQwERpbeSmXi1FgnI/7ChFjR/4qpEGAxYjwSyuz0uF0ZVbGlrP6baOa/dNe
WjRRdB0kMEwyhQnCa+OV2rKKURiAmxSNhjeOg7wGHZZ3WHThgUWoWiWf255e+46t235GbQMBSnnn
HQh+6HvmotjaBpxrXjs/cc3LPhWO1E53mUQXE35EDxswYeFjpUHzyEwXEOWd8t0yYbtdjUdWw8+O
iJBneAGRTT3SuqWuxujt7TckHeM88XaPygTQaCYRo3ppNYXC5UBhQPC0XbdqvBxzCuJEfvWLPkj0
kZpRbf7+2DYU9fPiTKdLdTwvy19lHFFnMlAzFkn8xKJ9h3pn4lCsxD8o8pO7TI0cJWD5z1GX5EQZ
UEAR3GAtj6EkPk8DwEodPQpZ15ybEAk7rLd2MHxdcZpUQFHwhtWM78z30Ew9KB+YbGFZS0AwSYfa
nTTrga83OkgDodvQXlHAwTV8tH+QJkiRXyf471H1kVkbpatHY2rf7bGui71dRVYBoGFW7TtQ8BZB
h+zcqrBysf3+Dya/oq0FRsoev1NtPkS15O5sE4PnOiV818v3HDMknWbmTsMezGWPcFA+euxQdMJQ
vDYx/SkLxLwR7YQkxj9eWr9+5AXTByph1E5zu/A2ywvp2zySGsFUGROsUXfODoO4SdEn8O6xt9gg
74V3PnbkUTUC67Tb0tm28jvWpSxF4LrdsZkwUWJLWLXqZCFws2QpvDtvAL7IzEXr+Od3zDFsOiRk
/703Xl4olof9JcjSYTytYZKqCTQqDGONzDUyn+hx3IG8d1qVvVMMvrPBKenAFgT2bZL92+HyFlGO
SD/GhH59Kg7iQfRyCOfbGiTbs+yl2LDUJVssm2roUNwwyYCuo9Yl2CS3SxtbFSWy1cnXNGaiTgDB
aeP0wdCoSDa0zDlixJw4Nwb/o6uZTT2uZ/qQXzr7F32eqXBoTgLqAwD8yPqkJYOKM9+w2V1nwIvx
ShT5UvcpJIujOzkMO6LelotNgBkg4qWSA34GID5ApQfvnb5GrMUyp9eDWZuj9rB5WhyU74Gukemx
jEWt0c/bDPFyLob9QyIr9ZdzfXWxsfftwAKE1uLaDRKB/8IAopyoPw91c/Lyc1hDfTckE8myFrlk
jZqecm3qD9WLPa7ushizEPWnZSYWarcqEee494yJdtwcA4FBOBBZU6KNyLkt93uArvPBmjLf2ycq
OoRkBsLFDhaqHmOoi80AMg4hAinT6cior0dr9YLVb8KK1F69CjybhUE3CIDDj0ulpj9NH0qKR7eb
t2MZxrQ7vwzlJGFfuJov0m5PFP5sGzXnb8q6x6/eyA0LoFQiBSxBcnzIopDQHk8M9NMv2/Yel/f8
rlCc7flqS48eA7stWM3YApYRlHAQaxoqsXezKrl3b2WbeT0SozxItlcm09HHSLnt+3jeQFwKYVcI
Fu5tGUfpZMS785ptu7Gi/pIUlqcqvVOdrUGmzhtsWg8gj+V/i2rw4PJf8+lR+Ma6zJmLu/RIXfbU
AhyJkBYONzbJwzHXE/0NFv95kl1i5KorMHNiOUqjaFJPa5XlkX7y0t5NtO9zfOnSwPAtuz8Q84yQ
cUmYN7AJKiqg4/2tgJe3raxN5nYZnzIkFHb5YF0MgOlQOa4sBkzb1zSIXIYFnIsQlsMthdGJvQp5
irB1+5OH/rYPHlAc6BZRXyQvSTn+mHIJNZWlpXURrgOowxautnp9fD4Qrx+ZDFLI22RqkIASdFPX
CZISuOIfVHkgMrH6U0rFbDovLPdy5dE8lygUnhYtRR+oK7up57XCcZlrrLH+sJXf8Vx9VTFQtXCR
NUnbZVjVJgg/F33izBbisj/ajLkOSHu5iFFAoIxwSU/0YkKq2mWTqjOVJQ1s2goYcUWrxdSx3R8b
BjvlA6REjjWU95F/Fkz1pyxoTOVRBwFIJAydmDHx+N7kPPY+604bSZtjsI6e0MhP/R7+cBXRbZlV
Bf6Q0fRdnXYlFIdGoZpuJgLOdZZ1j3Wsl1dWVsZJXoecQFdIkyJhIVUDETgRH4RmoPI/fmLejagJ
XCzsow+SoT8UMYgG/iGzhqt9Sbt84mcxW2i5tg3El7HWxoMXoYyiEe+ctrxn9VfAmc0yIhVWqEeE
wltPGBHZqHBzyqGHIWXbQcNUW5+lg1q2jjHGDfevkbljgyijkgkPBwpoyvechqjC5xD31n/qrePX
k/nMQ/7cnuYYbO6X4VyWqQiUf3Rp2CCYMHdNG64Iy9ScSpYM/1NyVAtSTFe2VWyzZ3H5xb7acStf
h8H8p9PjfESTsp1OJcmHICemRP8h+n1ALVrGHOA7eTfasNWXNBeUc3JeW8F3ZbnkL8zMkJ53lDat
VrNRL1bFnh81kiyfIZNA1p+wdOigMXihhyaExe8DXSTGuHwIQOGcz6grpYKfvxFo59JfbYbiTWqq
LWxyJ9cXCg44rWPuFG7L7COWTRhsz42OVZIZDH1Y1799hnM+yb5ObuzDM7NoTKL20O7CbtaGtb/4
8LD+MtoDuFL4gtW4kiMrKBU00AG1Gf0IAtDVaIpbJPCxub5d2x/dVG3qsQVVCaydvGb5CZxuJRoy
MM8qj9ZjWppwdixaihGBZXC86LS7T4YW5rclLNcpIqJIum+aBg2TCNgZCpBCO0+LFUl+/COFKBV2
GSfF7/JhnBH9L/QCvwJfMBzmHikPM+UJo5rn1sNo5QDm8WW/mdLb13hUeh+22ctJA+RI3UoMaFkV
+pBwOpLWLHFs+LUmzCIXpgmkKp9bIvH/8bTicbjLjLONQmtZ/dwXmsumTeTtDRBfEpxX2U+v3Xj1
7MN/B2cLx/EFLZpJdmEK2edigT89pPZDLxmep603u72rok0SUpnuGZWNNas+HMiG1teyMIQ+Mu41
0JYzW3iG52opODzFY0sEIfAqojnZcL7ngli9roz+MzRjA1kxa2nrFp08ADHuHB4vnamYLqKSIkp0
pkMAGCzDpYG8MPCPla7vUg0cELWfpWXW8/oGXg+lkTArvHnWEFJaTS6OrtUMeJ26BYJ1HcYl8vQE
3eD9/40CaMvdQpISkiugOO3DJkcpLCMC/o18mS0/n7hHG8KHz2avtg+O6hy0tDd1dIlipMGeAwFR
Zv/ZALsV8wvGowAEijCFqQMl1DgAkzQtcYXtfSt6DDXF9IXf+9bO2k0OoTRkdkO9KqgW175Ml7yM
/+WvnZiHU+EMr4IjioOzZQFFiZNywtvj8yIJoVBCjKkcbmbjRB+z5qSTUpjT+8oEBFxQKBEpCJ9Q
NsmK7uloeKbzQMZYgZMoNMvtGfsaaLdF6FrP+efx0LZ5XEX7g7RD9hO1GRiXGx8wnmaoVsjJmJum
Ji8QA+3hrsL6ihCIBVxc8AQgH9BrgPdtiFD0MQiQVSJr8rl7YGQv0d/pWUXTRNxMTdFD5MYMYXho
+4V+tifPrEGHMVyEqoiR6aFFg+9LfWnXOaDnbzqtbus923HLHiFYGQqUK6b2wwA2IkW22d4HSkOJ
O4wfMMi9yJnPdy82GPKSZwZ2mYvJB09qPWH4sxPtzqOPGiZz3wLpZav49C4Tj5cysbJ2ADoWw67D
N3Fh27+4LerTDPImlw+BrkKfRmI9Do35A/+gTIroGgpx2w0IoMz1B7T5BVh+lE17jhnxdHLssLdz
tNXaU0ffl5p63acXBLtn/bk0Nadx5lXm8fu9p7DmiooWe9RF9Ax4MlCITBxG5VBUxKS35GKejqxZ
1svZQbL96zt/2SCmzbE7fA6xxswTkNStBjEKg75QEzb4xG+7QNk+HRJpAOAu9iv3h0J722a67s13
VPUTx2AJO2slkKx8Td9IP+Y27MCxBuVLvyneVSJCbLOSl8Pj79arnx0/1NRwEgEevaRIkveX20kz
Pcm7E/vmxZunNJBD9pWOOX+ern+hKk68AkJyHhwaJXXYwxarKtuhnqpSXOVOfVGO5V19ux76wR8W
LAXguYUQ0ymBSu/Ajhc9jXAEqH4nZNMVHSNRDUpN33gM9niKXEbt9MdaVBDGbTJqa0LP+ayuMMI9
npvseEdBqSklQXBAKKnRzZU0YLEdEvE2jWYqaEh5GzkjVJmIvcEKpciUmmA03eeiQf1FK/G7IdWX
9hlXKT4fN9zQ9858Z1HeVmdwkHhbwVD/ihqR4deKckRqnHt5sV4xrYHNO9+zIwoGzcXC8tL39Qx3
IJ/k6sf9/Cr3JchNX3BF4DnjH9e/Ldc5v+UfQ8kduoLXD/MXW02W5iyyOZaRAe+cZo+wIemT6nOt
GJRCNhTLRLI/bH/yIFFgN7JWNayTrNpzaxK6M2Y5M8Et7ny80nUOy0bShEzqatu9nRzHcJotIpDV
IW4ehANDRlcF39DG9NIlOFdxj0vf+EhckUf+lN2ckym3TnLIYqTQnPBoibdiwPwnhqF9alq+Sk6B
4HQsAEiz0sUVuCES5Gak7+WMrRi//DCAbEgwwS8TIh8UTaSUxHgYVvGAH0cw0DxhjX4yhq0JyndU
/1BYG/LmaAGg63GyekjApagC9Oo8vcJ/sdRfG7KgAbWWQ6b8J9CKQCEWYWIn3VS15manyxn2W4Hv
7IXsngjBM71dB59blVsZ+fAzQWLwoOnpGAvDqusEyn84clnSPs6BWewzq3A4QixAYpU6NQCUY1TB
ta+ymhAhWA5lLoEghhGXUyBZzmda9PgAM0tEzWgOKFUCPEl+SsPtiUStByncu8fJlKQB+YcLSbLd
zEYBTRPJ16z7WAMFWQlnXIu8jC7LI1r4yzRlf3JnfUucSjMES0S6l/iKVkIbaADWT0LgtXrSD4A3
aEueCnbwdCKkmsaXzJrW4JUI0LBQ/gxfSUSPPSw9QL8Onzfj7Y+PF86Bb7x2HkpxDyiO6KgsLd+N
mcbfyHWRATyd904yrkxcjbBC3Ay7ZMnv2OHPnTy8XtlqWhTcs9RLbayqIz2n+7inF3Fh0I2WzdB8
eJE7TyKnBMSg5FweFJxHhV7QIof7KvqAsUR1XxtJ5TtKcllXdWpFG3Xt5rGAPsML5pieGc73lUJV
kqyZlpo8tdaShlqnoeWaPK1OhD2Q9Gd9X2Wm4bRAsmKCNnwoRnY+c3A+TYqefTjELKTdqZyNa7Oc
hTMqzdf+oacYXEzIM3pZjTacOp77kkciJ++qRiSv5/pSJ2keAmmVohyAMesiPJUcC4G5eRUBhhrV
nHzpPAiy7/qNhPdKZ1VWS7GXXZ/1kbBahAGTLw55jakhszz6axDiW16ct/8oehprgVH5LyAluA07
j5z8YoId1LtZuuWEOlOWLaID50PBC1yM1WVDXqFi8YOVo/+9u7q7nAdwvDukIGLemr04U2gaDbnD
qfbAA5ahhGpLoREfcKygsDTQoBtxGmgFzGBpXcSc5hJcXHfcUuEiSXAUqncNULzcYTS6lUu8InEx
g16sXPOJbTIrD/Ivle1fjBggIXFxQn/iAKEyY33MSsDjhUygdJQiyu0qt2Ujn/s27P3JwM883aYf
3G7Gsw2VpXv4LbBr74WlWnLN/j5h/AWKBa9ND/uStvsAXcJ0t+cfo+wpw2Z4VlqXmRvD+TvrEjMZ
UjizCj9LmN+8DvRuTHYT50TccG+Pv1jylt+wAdhWn02R02p9gk1/jxJ5fKwrxfW6z+NzEiYWN/3S
QqPEXg1YRds/Lj92O5J5Ue5tmlnj95bPlAjrRrR6VhPDgAuxogMHyP5pAJe8Bzv3gVmZR+DFmSAS
TKEpqdQZGn1N713MSB5NEAyj+hfUmIe5ySE5CDc7FC+kNOTKA8D6p1E9Fk/32yDs4Uz2ELUdcFxA
iNYr6ERav5F8JhlVeyYe8QdfkoYHbRP/Q8gJxvqim+14IbQ/OXF3zYxmOWfjwhk5LB7QR3UzwXEr
wS4DKJGMsAjR3QElRpbiT76e/zDUgTWdEYIhj01JDOais/V76rpdXKVCG95wEQofAMcMIaowb2FL
BB1hZfU7KoKxv9w6ZXDPBPo5gxIN1lN6vwde+D9gCkperLBqgTKsBP1WTfz/TpFrDoc2dbnAtYSC
u8Gom0iNxBvieoT36R9jIQiWsN28pkRZqfYtaW2ZPuNOI4Gg+R15glHuBPIBR41zPVWBeZ+BqKaa
sRfPUrHjq6E8Ixv42XwM1FUqIpU0mE5PrULSzC/HGjaFlWlO9GfQhHGS2eaIq0QLvs2UUhSYUhue
39Wap9xdqHmHD5II++sNMAOAWbhE00FOioUH0+iXyC5KQXen5fKYM1ovkB2A1s4O4yg9kqd4grTR
fxSNK2suMoE/XJGFFeyvRp6mVp/Uy6pBhORo5acL1NaXqRNScDY9guiNyo6RY7v2QxgBqnQ7xR9I
Y95GeBM6MIMjtKNH7t4CxoOwKFeyFdSAnwPcUWOm+zG8/0Fzrxul9HF23IynjzBziATNhqSvH+n4
e3CRvDWlUI2x+EnvnKzHRoxq/ttuTSZZGF2Q2uQiki96CnDA6zKG4MuJigQ03RurUPGYqGYRgy4P
9whw+nX13xv5uXHQUqzEVI98tGHBse2XHT8byE7BnpTWafRhb9k8XsRbQ9les1JhdTKteeVrXAYB
kQT4GP+tDSYpVsfYb/xICl6KUHhvUBR25Jxfi2qr+Tjz49SayFoDi1/3+rQ9M4pU6dOydF4r34V/
9cSZnfJuDNwgSzTOPC1BgACgqR2Dw9dP48NTj8T5z8RWuk+vLs1XfmY7Xw1W2kxA2Fjq8NbRLl/1
+jUuqE0EVTP20Vi+WHkyPi5Ha74qFN98KEneNjL8M7Doi5Y+c+PkPZ6RyybYDFinyScTERZluUNy
a7eLZI6rfN2+6QGHWQza7QQacF7c+CbyCYTcE3tVbnfV5bi+/B3iZolQVLW0zOCqCh7KS/FKfxnT
ViCN4JKECIHUMO4FRWffRTlmR+r6V9iITmcii9j5oYYMEUXtYsJsQQw+36cx28J9ZescwgAi57U8
N7JzRfYd3yxg+L9imJJTlHq6VsbdTRWNd/PWlFYeYMT0KX4Vfn8BAMecOpIRb0sO2lLwXxOeRkqg
gZ0sLSC2MSHDtbtVhOjutARNvZT0PN5VbsufCMtRp1g7OcDlMZcOfGjk4S+cra5V6HTi9aNTTfq9
P0yr5rHFGxS/ZGtSfaB11dN1yPpv5Fbfrra4/ukJe221LOghgfvvNZzfWN8R23Xs5sdsSQAAJlFA
xo9OM/8DOl+4KnNRrKhlyiR59OIKsJQzS6XxRl2Kk0Jw/x3h9qlCWSHyaU6dU6KyVgFfmyXSCaMJ
f/FXZQau/efJQEyPOWiwCdz/tSkAu0nxziVryVz9hii+9RkeSyeg59S3+/KV1CgRwjl5XVTOAG+1
jCeymIFpTyMc9FVzD7sS+UrL659MRNHLcmoktGTObTfRfbLG2BGNPM9R2SLXRJn5JrXnB0VrCzxE
Op7xAxb64TQDttYzOhH636yf33U+lsqd6yGF6GhhxfkOL0u6fy1+q0R+/3ZoiiOKAFSXX3iSjhok
IR3VbkLbFlf+6uWYKn4CXSHoOT6NR6b4z/PiwhqW+QFtLmuFhhyrpxEvM6cfIQdRZrpOINakNTnX
8ZRzvXw6Hv7Gb4lj6LoACyMh4XP83vIchC6KrbCaCPMrPwD6BKD7f5oYniClYiMjPu9lGnA45pfo
SM9OH7B2ap+ueQEMjy9zXnoo/XqTiENQdEawV9JZe1irV1wL8lYfZzl6yYkIKt35Txkh+HNaUlcc
9+lXquZVz3uagjI0Wt4odX2XpAdfskbXuAsQACu2DuGROKDxIu6KRSLKLoUAtp4HUZwYNObFG8JU
sokhc96Y2Hz282TBWXQ6QrUHaqmpNp/TIpQNT3HVOxSud2nMZ827uXJYjnJjZhDGjMKcwm6JC/Ws
Q2ah9W/J6iaOQrJDzMMoG3ezq4YoprEkZI6XtTs5yJ+CHbs1x/pCwTeh82Cfp3C4eBMwoDPQml9l
GY2mQRCCTK4cjrB9+DnmBm+rPDJXVvUxam5dMJ9iV7LQGPIO7di9zyjl/KPwnieMAXxwlNXN5FSr
nhaebchVkV+/1On3bKe/7WEI4sCxmqt3ce8H39LP/7g/bnyeDxsP8D6fxcdSoDaNHpI+7VyQYBWJ
aUkFaAH00PCM8WonxfQBxC0nWSPDnqQ29zyOCrAQrpTpNzCfzRdT0ezk17PWNSAkHbMhBGNlOEzZ
+rg6hMxFYrZb1+QaTt7Ir44EyAaoR0cVeYkNmMZnmo2XfyHfgGI4a8PGRmGfNGxjiRyO/8r3f2g3
YtEspz56vENqWC4GqdIwN6oIpPcMwij7/49IaMSVj8oBSNKPMeUXt3cpOBYFcDOLqYAAIM7BJD8P
XUsK27ZFLilICX06zAzl2JIpzomopzJiju/JfY6uG2X/SxzPUgy+JIEGtwpJlrfXMEaSyZXaYXC+
ZVZJYKdYWATSEqGmYCsJkiqwVDBryMFoZNy8myVD4XpQ5Ks8/LGEi91YUtFgm84cUTpKjbvOtZni
bvfTDQ2eNWTZhlrFU2U8XOkm3a4lJxEI0yiwamoxzRKhg9Gf5WyK6yFQxDtiL2Mxm/2KoywHIbs7
mndr9giH7smkycwVT3i2jucpiMzqsZbL+Ndp6D4scGbowcuiuJkgANz3V6EE3FQPjNpbHPMgaISq
v39qExdyJyeJPG/c5WvOHgRj1Lh/KVWqdJh4P+M4Yg6TcKxowKvfoMU0We2XyDO9y4620XkYjZo/
rc8wpBeVvAtTubojYGZHo14VMDbBuMFyIM8Z6ymWVnJji/4nts2r3aw5Fs7JpIHfwffW0Yrexcc2
iQ6uanZkpxcNa7H2RX/63Epk6pfF5f8v+GZbhfv3nn+XH1zPKTGxU5Lj2TpZ2t4yTtsTckgrLqKP
7qJAe/sJNRRwdLstTPSCa6yFEzuVrpU+XzLO7jrmTdh0K6MCvh/gbo/EyLU+z/ONaE+eRsVgMLmB
lkYdR9Jdpt1UocOjgOZ7Z1ijsl0TfzaeWkxcQkq1QVGRoBcZB6+U+dofjWK8VRMYqIzoCGWYxI7J
5KSnVhFrloLUKDGc7JFRWd0zgg/KoGNeWE53LlqVO0paALx+ZwPIogDuLcwMuOAvBRKJP45sFnt2
t3+aZe/ntvAm5Ax26znpwR3RZVurBnsvgTPUCTI1C34WQCpZsOjmE8UFRPPM6mVpxJhFHWSJoRia
ANnfRRLCCZ1MOn/mnXukZnvPmIjVdgpNxEk3yENJZO17P+cQq/Xg1aWWz8khu5DJK9xhO7JNBypf
g+ESZU5D/6T6YR7+MoQk3m1Vbi8W633wrmVlUcpQM+tLk8737HXx1qvD80LwYC7knGgHlGD1nqcM
3dZFmFCxAfoTQmxotocWp+TY8+AZBQJ6fFVdyPkbIpoMGlZFG0FkfHCtsT8aFteDqwdEW1ezSfmz
wWfMU28X066vKVUmf7K14dUsDb8lTq1wKGwBwrM2Q+LCLKEhKdM0U/9pnXNzAvUldGjSjvpJsUkS
ve0drB75yNPICeFEohFgCgFpq8jKbQ+052vLD0YvE6wtOM803BER9MPzKU2KKYAvMawxmTnj8OxP
0sw0Fe/anrJAM5Etv0jDDnlEiTpBVPO75eKpeoonF3egCrar085Xh87oX/e9QS6QbKfHpEAegt8B
A5YkuidFtQLbeCOxSyFwd2ObwVx6roSVWWGQzFu+SBlf5wWB3HSCGuS/Cjcjb96OPCFswLfZmm2w
AKIuUeQQfq0XxHCJYX2hi+go9BwzDgrkiYlbic8DXPd+vHJ3I5qb8G4HA/8tqRAdqJTJrmSBz3YQ
qGdOUnlcX2VTAyYDjoQpnVP7nfKJeBfeJjGdvL5TEF/zeZdqk/HohRYDc+UjWoSKztkRkUQOBIrY
xcwa2f+nnDrospDDDzCwMPifgHfI+2nMCahawAgAe95Ww/6OgxGsJNbR37G8p6yy+q6RUA0KfB1m
pwfc5s+uboxAr9x4/whR01zsElt4XzwsrjwwpEvnePSYCN7FTZKZBEsltBFa3DKIOO4T+gnYG8Ee
7saZn/AGUjgVDB57dIGjy/nZNRvkBZcRtPQ1NV8AXeL5f8ViQvmw8p6GncgWHXcIMNrSm8XgKEFF
HnU3eAEcpH/K0/ibBkDuWHH8bc18HLQ9JRCb56jNkR2t1+w/RM7TwMNEjjyvqkC6rRNMXf9Y9LDD
xIDidtAC44u2ONrYPX24oErbcbYL/JdmuhvaLFWTkvNtFPlC+eADrJaJL0KFZHZGd2Rajh3vBlu2
RTyyUUZgr+PzEQjc96Oyy2TA5YfcewHPauIGflVbmmh9OS3dml5rCkx06wwtyadnNwgUBcQ0zau4
ggTrf+jycJd42SD/7xEv+bFcDjidvV9WJ/wLWwHlDerNfaV4VQI1IywfRtrxprWx+UjmxFmVFp++
0/6DaSFwJlPkDaCUFrt+IoZmWvpjTxMKWEwe71HW1vv847Qdo186+c2c1TkoKRmaYiI/GyexElSo
vJJpONGyjc1AUt373R3p8j63fsPgvxkz3Pkb7amziCCsIn7SHjCjZ3q75jpIZDHQwKkG7ACQIkQN
Ydp8fxX9L2dHSvWDlsu6RaI4Sb2OoeemqQMyCvgCcBwSanu+1Vpj8fbHujHcsBJaKaDF5DQY7GZV
1f31hQzsH9jJhhz5poNUWXmf31vDHCgFqEfwyF2Xfgg7K3gGiBT2UjOX3JKUckxI4E2eNAkmlnoI
Z2i30E+3IsmcKHPaRP1d4sils3JimVEMtlk8q/ZIV34+ranjX24X/BCCAirV45aeJvCtR3ggjTzW
5RPn8RTmUhWqJcNFBOEkbuYmTlSLcVKuKHka1YhYZU5dYkJyGu7QvgtZun0qb6UmnZ6yk2C5/Y4n
/QlbVgrXo+o/1fYvMQ90jcbh5MTqQnPoAzT4ghfBzTSCkzkTA6Jmlta2g9zG9OxAQvU6OogjJgse
cVcrSval05rp8U8sFvSInoUmtCEjZHEujC8kWb4Oydt2i4mETrcRRsTFa9wSqGUF0aItThaPrToz
uAAM05r0eIdgObl2fv2jEaZvTU5JAtaXWwo6r9XfPHnqMbXm0m8bhVLfbpglj0FPEhilukV2/3JE
dietzwMB3O/mCALQdxlm2UJWqHJ6P1HPDlEOKht55PFZUDjADrqGxn/aC80EkRxSFr8/rThn7ytp
Kabyj0wswmQHlih+1ubrHYjV5WR2V2xiDYcNLPybGePdyJKKhAc3Cfe5VSJpSDOn6FlgSoyaU4Gl
f5vKxRni2+pcLFR4fjB3hoeA2ybwOBc8O9xNVFYP9x1rsQaCktScZqguglyjgmF+RKzJ2BKXJJ9s
RByo8vReyL9Wdo+CpFnoU5xI5G6uRO3GU93ZeqV/8Cq6zAKs6ntd59mbUsG2402m0IMElvkSzL3s
QOio28u+nMjQLhl1wVfhWjc5+JKN8UlhujQa92oJCXlwD9GxjAzfiyrlSqq/lj6HLO7/eW9WE8Vc
T/q4IBoPUMKjTgwTJjQVjB50LpZ3e6Eor58OyFB27+XRmxTlHBOnlntba1vUMzJAXKUf8zuhUwE/
T/r2Mvm7XAQhRsOLh7pUusstiktjagD9qe/RHqczp8TR1VxP9bTmR73fMCHO6w3C7gZu7hH+TGTo
65/J1oVidSQhhdfqZLt0eRoIC/iwcP5tl5eubAkW4p2XXXrNrbeudFyztr1dWdqoMg+s7eNX1Coa
y6h7FM0LQFSuSTptm2I0lJkNDdISDfmp5aPQsIfXIJDeACVHezOfbVSrTC5iu7DtHQiczg3WcOiq
1U1m/Q6k/qKKmKy6QkuZ8Bphh0LqBZuLK4g+KzN+YNE+AOxn00XlM+UpSotiOGFHVXeIndYpaoIz
wa9zdxrgfzs7vZ58PUCCeQJ8xKESpSn843GKq6RZvKMH7J29NTh+Fvyq2YKpw3Wb27JKCQeL+0uz
789u0z1EOzGj9HR9ZejANI1NYIOOjMaea8slYtu1feYCL3Mp/2E0pMkyAZ4ZgrT5knxAEtZSl8f6
sw87Wdul8UgthJ3JWx8/HVK+Wquf/y07uuKXapAKqFUXWW3TSiPoSdMsezDTMfuIAALUBIVOzSO2
kXr0bxCwOhJ/ggcbQ85j3EAa1EK2Jz7X9s49aAJRnyUSYBwvaetb/9eAszlA5ayTzI16V9JdKrZb
v3rTHihXj3bARxAzGBspegPj/Dw7INzFEQNX0vszdw2L6Vvuha/uyOehQdbAEB1bfJsM90OqXouy
aC1SHzO2cbbPNuyM8s9LUqJx77XyeVoJw1bC4aPne8sBze52DFKUywY9OZoIvkAALeFMjaP6Grg5
/MwAfjW+es3239wAeS9qKh+p1Nv/oWuTXhSeedy5BuQTAJSgmqjgf7gFxwyNwr2EBkzjOtoFQ6P3
v2zCnOpbL8WKAdrrHCCWT6wEel6MbUoiy6zBvLUCzZ2ZyFTAidHX7XrkLcxsejLMGFaqsqP2bvsL
S31gPY9fsrTn7gUWIExA7KaUxdi//5A0XIu4fVGs7BmfBU5pE8Ud9JndWsNgJuD7mkB+B9bcpcGV
pQ57MmpRDWj9kt/7Hx+KzIMv304F+V4BaGErRNbxJ3hhJqYBCYPiEY0zXk77aUvlRaygby87QrYi
9AmAAa2ez4idu6FPY93GGR7FUNeaTc+qkwwnoT//8WhsoBd7XbsTDzH2D0LpVr28nTKl8UFNbTKJ
hrL5tAcwnk6jkUygrSN1G3knSQqkANw4uVwj4qEKWCJlYbcFm3A8t7Nnc57CWV3y4VXsz5ZQGxxQ
EDPHWSaJGoKzK6fybtGnv4otPffE1drPjguZH3UoDXnygHi6oUkIwVRV47KJR+Enet5AFZwGoUwm
3ozgWOnpEqbELs36ZA27FqsGnjLFepUebwfEG+/S70ixcZ5tMQbz/hP9Oe1VfZue0ETK1j37D3EH
O8EB0WneAzq3/TLNWVpRU1ofUmBKrcso8KeYnfoUWzot/0jS08p51+lLDAEwmI7RNV076wvTf09d
S5GqAA9KlwUEXnk0i/j1J4NFMOu4dx0iiuZOshPbHDsbrBwHa4Qlw9SmqmS12HKk56ty8bAFmDct
uOzgEuY1sr6Pn4eQIUo5u/QFJMlbFaO1L4y/UARzcbgBmA5Vf1rzsKnDha67GAM31vTBmLfYYiNu
5/uWwek7gtrGP+QyOZTtiV5ppSC6qNPaLuzfqJuGwdbiCjsP4Ff2H5FiyDjEtNbnBd0NTKDh4zyg
H7N9DCBtT63Dz3Mw8h8T2PmgWHjQOpupWH8HYQ5wc/iZtLzbAFm2m3HogkPaG3XhqlmGN5vEXsaX
anbOT/6sM312U+AXhkR42HzDXcrkAmLKi7ujFWej0Y6wYQcItgcizZDP9/dVIIco8SkQVXK5bChJ
ovKG9ir2AY4FfcqxefiDKH08CBIogDb8g7tOIdOWcm82+8IA1yWdP1I83zRpRt3xpXCSz4QGRTuG
eodJ5J4HqWxHl6NIfvcNMzgK1Bg2Ik+MeVbL42kbiorMS+QjCEyNUJYctsQ8ON6GneS1GPU6DEh5
Wy+YZjAXK6KwgwIg83daKs7RTjzVZpIiOb8KRP8B3Cqgzp2iQcS/Bu3DYvhYhArjRMX4SfhrHlNe
gsCW+ODcySP7NMw0e/ProNFjt0sDr9FiUtp+Y8coQrrFBSiCwd13xv+56RUePZoHD5pXew0/t9Kf
h5jiW0ONFJozWmtSt/I1t8EzVQGef1m9sWa+FI8W0s838PO7E7wGiOSFr5YcMklkLVvmQWWU9MVF
C3zPYoACM0tQfg6T8yhBEwfbvYeoIkjvUHFvqDYKGRDUEqe2EDDGXZMAh/3vg/zOljGxNMaLeqyO
o6EpO2VrYIkhQXKUyutQ8a72D/U8R/4xN7ABtUd4Yr6be/NcWyGpGarEseGCj6ldTqcbiIcEDUVP
78vW2P3+Z8myWXGk5zr8SuUw6IUq2xKmTNFfU2uDFlFgyxUr6gmosDQd68h66oTglC93hWqmYxeW
wHy5/EVM1DAnl3m0BxQQi/qTUyyVtFh+viNgcyqKv2xYlm1fvPa0pT1vw2pxIeQGFKRFeR9ViyUR
U8P3+JrqgHi1Js7WtKY10gC18MqLHgx2hvjmg7nhC3YLLtz2lPD69RQYC/5DiA47YQLPHJQzUKRm
UERERRQZYi/bom5MCC5QFYp3vJUy5NSTaEz4+7AYli7JGWAnLJn6NNSHys3ws9o0wbcoaRrZF+D0
baBzjeemXlUXblvYYoqWRKoa8Pibieg4Vq4y2M9yP1faphnqewD90AWWq1oH94wgmO7Rl/eJ/nqz
JZ+gXY8RfPwjZ7N4HsQKQNFPcwKSw3QxT3GSobFvJKrVjlaJ0JZndhWK6+IH3H0oi43lrbKOJix5
W85YvuSYzEAuvMzOIZZ8y46f9qwPPKxY1bPhsmWblKQnI8pvTZJMALPEmXv9AiqXqzyIT4VI4W6r
NVMUV66Pv9L+ekLuucvUKz6rR5eeWtZ36exA5QA+xQCZBjwq20JV2AVIQMgfN+paFRc7bgwKqi/A
ChsUdtRwGPJNxkHI5hHnrIasWyraXyAw5LTmhS5Tzi5csA8LuWKVSBFLh5BiGTq5zB+yJyPVVQdh
c2Du89KdM9ivWqbd5NcqyKAAob8DNM+HZaDlkWRdNohxuWzrNziP6638Q24i3CJ6yAdwuLSjAP5X
fCWlbPB9luwfobeET22HYaWZ8e4ZMbZJwBP1034+den9V94zL+SmIS/wgUg8YlTNfIDdqodiao46
MHMtwXbV2J+wTULupwQkWQPxCC8smFfHP7i8w7EW9Dg2RxGEybGHpefGp9LardGzkzXmFP1P1RWH
gXrKob1XZVzZo38y5Wv1hKKeKx5jv2zhkzsA2Z1cII9X4kfBv+j6cm+tDdIfcJ47Od50wh6GNgCR
6OYrUjCn8d5ZbrIMR/UPlSzON5y3Va3G8N9HYCvJOO0D+zHqqrIJvyjI9NZvEsNTkjtE2i1rdFGp
2IJ92GgNvNCmT+cjSgDtkqCt6MVRBQKKNh6cIaAWStTqJtsoWJgTB+Fhln06bBnqoZi8gRmb6o2s
Rh3trsCph+qGEWhCQMZH7FKvkYldmZDXxTWWCyS8wrUilBVRgPK9jQU9k7xCCvOGQBYC/SQwuQf9
RD181h30jD0pczvX/zq5aHc0a6Ilo4FEjvdXOXiIbx8nRyEZkk3qrILlXjUAxVs6uEYSKKArcfUo
lQeX9p9S5HHikyOF1AZNgaylgPgLOTUq9Qqn/4HG2MtjWm8V5REcwqTw18LBykISeSDRZcKSs7aX
yu/TzIhRZ6ZS1KNKp3ITGElM5Ymyzib6Fr3PurSnSMLCY38iVuZRZGN70ymy08kUdd1cILAyFWsS
NgIEdmXFxhFDGfZ9/xdtVW2kUhuw/FzPR979Czs/FqbOxR2FO6CXsT8TcATYm5mK9rr2c60YqkuH
X7QBli4ehfZUVUZ54vrrO03F2vJ9lB7fhK201b15zLOcAyk/FEBmE2bLtw2zPaYmiLqqAndZWXEH
MrDXryf8q+1FRX/7cKIwbSC7ZPm/vJphiWu2GFQVd3dhfmcF4fVs+y8ZlW+CsP8tr9Vqf8OGNz6d
yotQlAULVfWsyyxVnuKL1QUoSrRbQy7th1wFSEjo5MVX6h1aE/DMfyCfhlUKWXFPOkdmD/HPEMY/
w0d3aqfFPht+qf2ozIDUNr34DrFIR5wH0IaDJ/7aDRUF1FnhKEGJ0tPvASWC51V05wnMGkSufYw4
SZAf27xt3LRZLGiuLaBwmQrRclpZwsWNSZZA4ibbu4NvXiCXGLlykzvaTb2qLOUmqKYnmC7STWKb
J1H8s4Jq+cboWIAFxeqyfNG1PiA4/I76BhSlnZEPpfaWgjbg//Vt15d58F7lZhVvT//Sw9NM+3Sw
QIeV00C+SGfCviquDS5Q7LT8N8naHf0wGWIzKZJjDEVhXt+Bp97E8yqNWISBf+MHUKZS6Z6gVcuS
usbpksvpSqpucwEiaTr941Z5O6tD3GEeF1zCXTCWSVkLJAPrZ+vK6mgImy+c6AldNWbQERpIxXdh
UV8fxIMDksKuZba2jyXkxx1BtyecSi65U/nu8Z/XGY4fHZ4Ckw4c86S5NE9ZFA2w32RyMAM+1lwq
ZYld3fXgP8L5muJuVvLjRm2Y1PvtJEuCzg88W2Ald8Sy8GBxD6xHbGH0kMwFcJ4N+MN+Sa6QhpkQ
+7yZh1HoYbl5wKCWMflOAKncjGju9g4aS4gvfeGKDYGXOjq/SLtUPN4O39aV2Q7KJPQwybtBnPUh
M67kAyEOn3FrGMQp7gFTY+dvjd8gdZFpRnXzL4ucAuzDqSXdiAhDz7suSneCRE0iBu60Su1d6Wwl
Rwpf4QMLeYdkW7kA8NYbOo56jOf1bPdY9pgkJNL/00PPL2yL4uCKKDYzll5+DBkUsBNTK6QBHr/b
MRvK6Lbr+PIxNWkK1Sl9ChxnI1scPZvTpQr6IuipP6nm3UOyKh7D0eI/JG6g+7MhmlhKopwNCfMa
nVuXdWegyzJUvJaOHgKDhJdyddWvsCUOjixHce1wURR/r16xe46CVFOEbUbIQlF6/Uyeeg/ZPsjM
SuRpfryQB+sRfN8V6F6GqAdPUPYJJodboY3V123IxEXlzUVsuftEp4UXjtq1qbIzW0YbO+cytVqe
K7MjGshLLtJRGafmU5aIYJbDhbk15BiCEaeVc0A8khwy0Bb3oLvIQr6LIZrxchJOy24BmKQoL30Y
yP9I8sz6FjSb5CUZcVFuhfFCvpPODnnJWO/n2wS3a3WeKN4pnPQ9WMbV6OtH0CJj2K9tnKtMUG/T
b53FjuDSy2SqiHoYqjVr1FwUH9ixRU1GWS5fE/4+05Rl+JSWP1G+/juaOE/TFnA3ZXmz48c7+BUG
llIIKy2dI43IvQSp+PwMGsy9rafyvTqaoLeu/kf6oe/6dIRa5a14lsKpP5CUAhpt1CZx7+KMAPZG
si93q3ffY4mgW73JsQcl6a7IcZ2WrAFMlniq1aQxdrhygFzu43TbJsj9Thn6cKfKnxqWneHkkRqF
0f/r8/zyXPkghA3JZE3n71+wpq3eT6TWK8ADbdgwnGEg7AbteecnwMEH5Ty8MyP54Bm/1C/7PdF/
rJNLlVqSKGewU4rbEjai8LsiTVZ401S2hQYhQOHRDzZ/YQg8OWwX7+UT6ZTTawq3e28BnmI2AnfM
eCmGxnCCMYG/AODqgeeJGKXfFkz0iEH0iiGsO8XXO/FwThiag7je2/4NPeAqZcrBPJ6xB/AsqDzu
KdHL8jajdWeHBInDVNSdDiBihquRp9ftV1/HdQDkbzZBmOfWJd6ANqx6AIpdeI8aarMbtMeDyHcc
y99zdNF6kRfcdTHf3vCtRi3bb+AZEP0wdjnGEyMU8ijrRob2IqS8hALbs92H95jndabOJ2QVClgY
l0KSvcE0PpLWh/KRnWNulehusaaV51zXViLfWoibI8PPmcmHQfRb87O0JJENZF0mRjBm3Nbgn72E
iBIqFpDRVJ8JGNZbKxwgse5RMmhmkfRCJPKIGonrJc3ISPhCjHzi+sj36mF9l9tfvhL6/x0BqGcg
b3hmY8t5hfeE9KO3MvMGL9KBgvQluhYuFdUPZtZ9aSFSC4hdNIFTciLmqugY7T0aV4VRReW7bsiv
W0cSj/k17OmbYhIWuWEKrCZlfnd4/oWOOd4sp0OHpx1mZjSasyAAwIhzoUpHCsLdp0haJl82Vpzq
1G/Lyfmgt5F/sU9nBtpifPTNeFntsoXCPpRNeMQKkQlmZgtqf0mDS6mWi2nEX8sK1rw7fkqHmvv7
P0L2DKtuPMe9p7mxWQkn2hE2Hyt9ImNjsZIrfWUqAMGwBHgBOMGbWgTI163NWnRlUt3/ONNsyoMw
eq2s+kT2MHk88yzt+1yB32hmSgma20LxHwZZMmJnzdZvbWnn0yMX74xULFyLhoYQYXvio4M+UwVx
YOCrG6ygzgsMAw/VXB3lE1DejueUyzkV4zn4K5IOM1eqgCiQ2EcK55vkH8zF5dmmItPpPwMpN749
W5Fo/zksUoy8KWJHl8KO0/Bng47dk39cHlXLFrqolihSALgOcOTm4++TlxgtEaT4NGbwvwMURcaG
07ke6LG8Wcrt/e53jdS4eCqFy0yvvHV1qZRaXQ0IWHH97QdsER0+c+fLqhU3ylBeUUJYE6pt7Tg3
8dahi1iNW1WgVdjoEqW8GS0JiIC2/T+6gYt3kORQ9+qI0jbBjK16nC0zS/ZZP+S4ALyBK+6gmgK7
VWHtwzSykx+AJ55hPr59iXlT0MzmvECRvloezAH4mKKj/lr7pIxkQ+Q99ezBq7bKE9tJdfS0v4gR
1AFYCcb9hk44NKMQcCib9M2yjZespAWpE8zEMESJyn9GdHNNV05EeVNtWmMAH8sjuxVZZtSsaIIx
V1CPmiWXW2W3gBgxtpvRR5AqVNG/URhQSuLUwtIlL+VKyg3tmYCDJ3grOnzyWqBiwQOuwZtJkdn8
3/3/gEhbYtEtXQFieIBVMkM2ih/sILyA4Xmm1seGCbqvOTss6N9xIRBUckS4s+CqeIcxX+bE5MCt
3Jh1MTzFN3ANDwWNHuYsDOE8JKzJeHaAALBntNvqj5jL9f6N0Ec+5Hfu9wQIS/w4/vW9kBiHjfe9
fOLH8TWmLhSshsTY/Me0TMCxLiEZDH9QIX2mPV1wdzs5zPWVcVY4e1cE/QTJSK5GNehqL89iYg1M
0iujIZdfr06RwY2eZJl9AkZi4RfQ+DDLRQkzHACL4ph45+ArYm6FZMlcpEIJeacjDHIfy2txhpnf
IAetzqyfUTn+EgHMuUcnZzz9GCEOOecm0LoueCcvu9Et/B+HvTQgVY6CoT80vdrOaaV8nMopJz3a
KqFy9rQ0hfTyzSXGPrrq+jNixj4fiecB3WdnMIm5XyVqC5ztaXKUJIYu3BacyVZgBlO4uj4ZtMhq
axyeEQNcJR1roGMNTko+PfYRPrg/79f1NKAAr1tgHt01t9/Xpmg+3LR+r30GLWaYyhw0Npo8fOT/
aQFiU0MfAk1tQChrJeMuSXxdKhblFcLdvYiHwP/jH0YtzTu2BIQlAw36OUJnKRafvqExO+yZPmiI
VtZwUuniIUK+BUHlNy4fAAdvlO9Sph63eoucy6u2YWaJbsLj8WafIjSFV18UBaWW+u2fX8KpSnwc
ubdWFlWE5mejpIJ2rSpgehnnsn13CXS2WUOxdtuekId7ft6XeRsNr1thfFAL8XXbtuUpxe7+FZ08
mLf3CYfjfYKM/15JUKIMn9/gXrQb/U8N+/gmHxS8lZ0PZUA/ZRFUJE7BlWWG3ZoNAzEtFmSVgpCc
JNIZMHsMZ9cYflwzREYId8qw4wiTxsAp9XiIRdOSm6oB62sGe4NxXxmqlFlXLtzfCMmKLRavGDvS
czc0RvN3W0DOkXa9lFrQpkwvGwUY4q52pVNfB/IvFadJv0O/QIP+QigWe13U+hg7oEJ4iu6STZ3h
pPJHHXHRaZYc1JjiTncqblNv5OkZEh8msJBHddU2aSxllH590QccxbhHsrhR9SpCDUkU6A+Et/iJ
8TKJLX9pK8VgWQa0gmcf7Qyd4go1PLYBtIswms/0KmXpxW9yWLYm1Vyragtu4b0a6H+2gkWhl4LV
om1iWatcNOUtriqy3pcO+HPqID4yg9VoTTexXArM2aaSzh/nO4zFKA6MdX/uPlwi2jVQ7LjMPj1J
ZqJSdSBIJmbxpW8Ua8rfpjRb8+f/9Az5JjK5aMeyqFKeOEtu1DKsVFp/5ruOZ34/ljh7zSLf5hRp
vLXoCWaTrs/FFmmcjvWyfTD+eCdk7hJMta74VhM71x8oGv2GZ4TTizcfl5BzM5VxvbGJeiXC6dFa
fURf1Wmcv0RniHN9XRPmXgl6rymuyl3N6D25Ri2OQmySIwpt7cPGTI9eQYEmQ2j3K311HYbsnwYg
xnY04UA4P3PJDhoPCf6kYSvjWhH3vdIwxCUcwQ4Z9cImT5gpuYuY1MucifM6YlMhB7k4kPLwTw5/
/wpwbpP0fWwnEFLxHR1VFicp3B5oNPPZljzX+rRxUf3cxoR9HRrZnFTji/HMI8hrtcemOZ0r7od1
xSD2B3vysVueHuXzFbfaj4quE8yq55m337iymRRULdu5ukBzblwRYgwzfNL+NN/xX1cjXeT88KYi
HDe0Ck9RYAAGxHvKUhraIUO6VqizAFeYrI93yNWPcZdivX5wfGSMqwJdFEQfGn56wGLe0Tb/a/xx
htVAcFj2CWM1jRTTK0Blmxa7/spZLio3ZWxdVexE7ZBzk1mrDBgIqO6QxTY5zcQ/PYcCIjCgQ5QE
OTxmcORZybbqDxhbdB1qT5rPwJWzPH+TdvAaXDmugB+rMOgciNw3HRZfWODSIIpuUuGo58LBwoNo
u6g2KW9xjF/I3saeshZqCNJD83w+MTXgl62ZBvMGg5a1srBbXlSiDkGQ9BMsahYO0xFgdfPEvOLm
8vi2CNcB8Dnkx7w/KxgblRXaNOcXiZppEn5dscAjdx+KgPhqQdIj0tUeVIJ9bVhf3uu204DElqcr
i/nfwtvek8y6t/ROQZ37C+PDBcSqRhLuCGGXBTatwIsLE4/Th9kX+iWjdGYJKAW3AH7Yb6DujZo8
i51L8J5VTxmCFKvjr+owPZLXJmLyQIIFFTYjLXGytoTcrGqForDWrAQF+q6YfbbOpzjBXrBAAFtC
G1Xh3PPLuua57FNrf+P9xGKZZ0uLpYsmni8uMIeHYsTwUg7HBbagpYJf2WBsKRguY6DZXr6rMl9R
b1LXK7/bIHZUh62GEtzNHigC4te4L+E1NU2T5HTGy+qeaQLWfqtwX4pxuUNx6fYJ2DxD12dOfNM3
00CrO2GzNCsQ69vaRZeEPi8w+DjHPmoR3zcOeHDMBHnPS5aSZ7eUQLeJS3L1RrceN4n6f05FtzMs
B08V4bfeUShJZAgwA95m3mCsKC3o/LwHfx5kpqMD5YPoO0BQTeP2ro7vcyFNF1h+4oqtj7dMGtpM
Tsd03gbFm6RRIcWtreL9eadvrIggkhtOYszY331j/K20y/BMbMNUmiAMtWvUQAdQLH5g+8pt7qDT
wmEI9pOjNPvbvUtv5Duq4LMOajBP57z5Ux5zTau7JadLgbSmMm7WMQ5Vs8JSqh9kkKdmCmqGHae5
4qDhUcj7r5G2cS1aKBg6saARry6oato2YkJuYXawnG7M3dCgSvqtzdjrpQAP044AkIsrwu6nma4R
vHqTd0yt5T4WfsV13+eYlx9NHNGwEC0dpOBl9z2I9sobNZMv9hW+m/HQ/vZiT9PwWv20WCr7nu66
wFmnxdS42Vk7iCoona2VaX4hDsSGZOxrRuDZVtVMuPS2VtyLf9ar2OpnKtCxxdcAFVyCMm/K7ri3
vTc8vHy7gutDZKeK7y5sa4/vAwL9KUwJJ3766MzSSvXMRffpNXlrzBQOUnW+3ASo85QcXEe2F5yE
lZbHJ37q6mDdAe+bZTr8WD8z+E5L4KENMDCLOtbiWSl43pTzAlggWhTZ9dPctmAbkXrkfkvrC8Yz
CKMyB1MJRq8+AEq9FrIGOxfSAO1UElmyO0Ak8EC6j5TgSdMzwzbTdHlX2VtOm6bZKAyveadOKZ+X
uctw57/qx5y1xzIOr3exkLYdbffE2ul5zZpuJ/OE31rGOCXE4VLjNtrdLoog/vPzCm3adQ3HKgx8
7O0V2j4rCdM0oPu6MvurM5Qn1jnbGIr4Iv4HKxfbfD28mg87XDjP/j3rvEnqDcfHst7PJet6qaUe
XRdNFpIpZ5s2gGeb1AWDptvnCDwgKFbz6U+R7yzN4bWOvr47JfCehCRpNA203UYooIagoNrqljjA
lLGvfdj46VA7sjtjPcSTjn/D0P0MPJOjA7UgajG5KaccowpFTqcwtM0PpzbEHGUDBsNJ3TCjKlm7
3pRLmdqJRu3JK8iqflN4gBxaLyFCzy8w0+hpa10O+ly1GSBFdGVidubppKu8DeddRIQa5UuexfGt
V0Er6FDLvx7Og5dHlbMlG2kIqfQ/xH7c/rPcve4SgIX8xYetm4fLVNCUROTYxeMem3FAKTynSF71
ImQhqVOYr87YVy10dxGxgJz89tF8q634CcJkTO82UWWtZIoqya6nCCt1WHXGQx9fck+bXomaf8fm
FbAIIF+wAtw9NM+5u3BjkEdMW13XGhZvO2EBt+4+A5YDwYUB9d1ZzaL1NxANY/v2MCmOQF1/JA/L
mPSi4T5EtlQJDfTdNMV2LR0V4Y8cTbERXGWGVhC8Dv4yryBKY7jXjl0pGm27TzZzRQnTFjOw7THo
fWEZLdTUkzcKKaFdRDnnq5lA17oEPC+vZH8s9TmApswWsZfU4gm53DJACVO0G5jcU1EyE8oM0fhB
vtsz0L0zplsFDzNlH1VTRv/wv4wfdU4PNfwrvESyV5J4pTr7A/rNv54Nl+OI5kDUh1lu/lnX1DB9
S50SR6W7lgzk2FV/laa0OycQl5bcincpN+vBvB48LEq8IFSAfJW+4B4MF1x5uudh3p8R6QtLC1xv
NIGBnhUk6+b2mSBMr0Lj5TnqFc6FEkfFktINERD9YKR1vgFMlp3Lkhd/TGTqKQBQ8AJUE4KfgDpK
L+dySXkWEkk81bSfLnxvcJCK/A0+pi2TBwtG1UjYQ3waQOl7r+rm5v5rY8KtuLAnW7CvAQ1n/Qj2
JhA7yWlzM9sQqgaJ8Z4WF20babELTOYYHORJYNx5+smqaSGA++yGah8BZ+sTzjjcEb5dpHAREzay
0WudWuUrVP1zbLEPKyAcc4tRruVFUP6lNQ0PqC+hRAZJQYyhoaMdBznEQQ4G+E5ZeTB0/ibV5S9p
wndscGAnoAlGU93a8+IrgLCDpOoqtmBuJxtd6UQklAmX6fV1eDbbe+fM5L8YpH6IUuzpWh+SumNU
s51pPPotHEmlNQmCxk3mi7/5rMgvcW4ETEB/jJyWzg4gTZ3Ht+vI53wgp5JcVQDprlPUtA56LIem
sXK0bD5+P/MmCGXJ3nY51BAIeJW+m6W/uEF8vJPXNS987GvAzdbQb2R97VSpRE5ECOWEPmj7QMJI
jwh8Sc6Mdc7+u0Q5/zj13ah0JrymvF6EDJXijvMSZDDNsqkQLE18AxirnTlLFe7fyZsceaccdWHV
E4JcKOSgzP0kA8qD0eZV78MajzUNOmFHQJHkWGT7KSNm3MBGPKbr+NUTlwrgpD+dQiuPt75hUNoe
3oBHYAfwXcADkESETmHs99T4FQHI972kJW0PTN3rUdG4rVsMTErIVz6IOoGavUi79JghoX6c+n27
ixDCWPQ70vMynysJ4SYXHyF7gSxDF/3NheXyBkKoAt98CVjRSglieuCPurNGZVBL+urq6jzaGTiM
GmRgT6wwGrI1T6Vh+6kmxgjJB6fMZUQvzbo5VFbGJKn+AISGZWjp/FZXfuSOhi2mMvnWYABk0zJZ
/dqsVz16jjCFdClNfjDxu41sPVe2+FfYOpsfz5Garv8M20iXbbC8xioVDxKGK+yKLK4PglIz0R3b
ZaJqzAMOY4drsH8QNV2KO0YR97OqUDdKbFu6q4MtMyA+DJwn2JWv+x8I8f3j82geRWKCTEBTFZEl
1bEVeW+64gEFTSugeUwiXYuYoyiBaa4MVhalFgITVQz8eUHS+zr5GRGMPO1ex81fbhejCgqOQsFG
cLZUvE50CHP0+bKVGFgFdVgedIwOSENBhuwGpx+VJFe1YH1gP69WgfVOGBtPhmgJykjPs7geOxz8
vbeRiGpy75VFIfd8uLnhfoIR9vRLuD6U35g5uz8pQGZ55UR7pgYYl9lpB4Ti7PVTJadPHchELO8W
UUR2S5baX3gxHAA1wE4ttlIZGRWALav/cRSf6ctLsss9lozQZH+ZzMYQLX64W3GasbTRRd18QYlC
OwHSwzpbxOyMI63vyoFpz71UBU28I8ZB8t4RhJQovvAbyuDteuJXlVe+JcVYK7cGEWeJhQazn2L6
2JP+/DlTbDtEB28urAR0Wnd+YgqP0OM8oLApwcg5pMQnU5HlZ/5/my911SNOww+X6R0tSrS2qTr0
oEvn9aHmqDrnsGvTopzAux0BbpxF2q+jV3D64TH7InNo/U8jKLpnQgQ0HLAIqfN0M5smO0+sTMAU
QHKJ3EOtnh/gGcd8fXFw4SuA9Q3YNqZPe6BQncHWjjQnnK1u4L0cfsLLjTk0Dqi1TQH0QvwNVm/4
QlQbx0e/cCRlaPlcsWf7Sq1WkTPJqmspTJp7qRkMq08N1OX8+SO5gwy3pTsojl2ZxhYRBAt7kReg
OcW75FAWM/16fZB6+qrAbbpZpha9VjpASz5NzakbtYHOedDHKSZHimDssNhN+B1KzA3U1hQpvffh
sND51xTtTD5ij8J1zMT+4RiZ8xOHP5T7E4ERsVg3H00NKOww2SImLyJUK5z09NtjhD3q2XycDH6c
BfgfE/GHgqydWkW/B54pCAmEQCVNB6AJOr3F37q3hOjiHJAYpDdJHjFFObFarIfwWjOQBlZr8Y5b
fzX9aJRQZoYDeuhCh16k/01ykbXYW6MDF33mZIqg5mwOZQxLWS/T9yje0bsw1clkNV2AznWCy1rf
eYGCtlufrXTAf5ch5jmF1zxqLEfTWM95rxdSUirVFQgDGk/RPQNMRxyAaTH9sCndipsbGVBLs51l
JVHiY7Imo1D97gpGbXSUVMaFCGK47O5K4xGTJTzAoTNNHtrjKea8fjI5LsvT9nHBLEuEe8Lc+Eck
+/7sg5+2q3hf+T2fT1vz1tGj/TUMWCuOjhU9fDTcx0r4oMlNC6EQb89pA4STrDe34cGjRY38pTfZ
JfWfWU60S5UHfqMj5KNd8kwx4RYqIH87MAhpKOkp5yqIzW7LoIYPtRJtJorTHM5JdxS9w1kSXsN5
rU4XwYuwH0jaN1t83rezCaQUAG6rwzN6nH/pJGQ+bJPcFQMwSRDy3C+Npg1HvDs70kuCBzP7MNlO
PZVPaSYjNvKgwhGqXimzKsiat9ot40g2IRI3qJ/OuQDDLEsdAskzKrPIlagDZR+WFiVmhaMMNz+1
Bc5Fg63G3tCl0Oa9oxNzxr0B+meDX6WgZUcFm65Ve/pk9zOnzwwWWJ0rIdnG90uflbbHlkR/QXCb
W8FTdDIGaFDdSj3D1E+gSRWZAYkxD1vm2Mt3gpuPBb3Tc53Zji7XuZNmB190SmvXRmpGJ+SZf609
ZgXhZ75wGSzAsQRv77BTIkthGnyeIsLArvaFLMaylCFnc1VtAz46yOEM+yN0Nm9ndMFzBq5XWFrG
3LVl75xz9qOjvnx9niEr3axTDxDhiDRjk+QOa7FG2YvSDjSpfgXKRvTLC6Y4z9xUbtO3W5npreP7
VK8isiEZ5nKnUqA5TT8m8+MVYqmwaa0J0qtw6eI9KJwaXX2aGyrnZb7PBlqSlrQsKLJuQjOY2D/s
Ju+bG5lUCKPudxGhufNleFp3s5U+dY0DIGcWzhywCZsk2ZfYtJsb3xtZ5T3SHXWLHpBLm0KFhMeb
irFU8TAD6wMRRsQIkP78DIZDL/OrCL2k5Io3hhpEz6BKyJ1RESm6BIRvUuK2AVerrraQFVKG/Fd8
Wu57iwr9UKyamkL/1kzEg1/6EvNwqkR0S/Mem+v88/BiKp/Vun/Rv+GG7d/utNkbExf6Gsfw7uwR
8XWdNGZF8y4eJNrJjuE2mbSt4edudgzn4LAlpfuG1tNGhCBfpSwRpkm6ElGCIAixtNmVYrwp3JSD
r1wIoL1VaT4GlF4g+3WbplUX3yZuAjXqwiLqsSZ2+WDnB9mENRbe1QFqptVXdC1UQ69XO/v4SmDa
GZxZ6dploa245bHRdjBK9zFthyUZ0Y/oISvmsHBXWnuGaAt9X3jjsXnklyCG4mSTcJot80pEX8cH
zGSCeXomf9gQa9gjMxhL3Pho9wEUrfsQQjSLUOgNA6rMKYdu6dOIf+8kGLNn3pfXTYHokbggXqU6
4VRfzJqSTrzs0128fi3HXshei49dY0y9RCaWvifVY9BMVTltbfQIlHu/EVPm5nGqcOGupKdwHBP6
zfJjazXuwBK8E7ezUXeDW9diiR+hcpdIJVInaqUbGO2AqfWNpeEjRRj8DRyFGjBdPkFcXwSKk+xe
amQdB3Y9v5zplDmhkNowG5CS7nDl0SUlDkq3YQKGMRKz7Y1rJROQaBnBtbI1mnP6FajD3+01E8OA
83E0Dfu9aFmz9SEFZCs5KIgps0E1o7czGHh8KpHtjYWGECZinYKzYCbHzquewJEjGJmE/ZP44rKI
AK9j7JozK3AUy8/Rp7oUq4k955999V+nXP90k5pxjZhu5gVzO3N9Z+Tcr5z6ff762ossG4ki8Qfn
ATMK7LxKiyWT+yb/OfK7+KychQHs0qytvdiP16A8Dq5+YKlWFde/ipSK2/Q62mgYDhgV+Kn29auk
0FESk6CyWc6w12QefHKnyWeCMIM79z2wHjjfXwcOAsEUONw+mDAc5KkkhKBgcAzH4PC98FYiJ+TL
acAMNuMBMBLMe0UvMpuyQ0WbLBS+qfIdcEclb5G80+LboppFHUxM3D427y/9zDvz93ZlnbpHaObf
JI83IYuMiiVXEeYFJR49uaYeIfAtc9oItWUJZ97PtH694QsDFFJNhtzZuwcYSow2/yE8hT67w1RM
ox3wJmFTYh0ZyvV80uj/+YobwUcchEHtn27ffQ5Itzz3JQlefgs0BlcXCp8qZxAqZh0wkfrHYjHV
DCrK1gaqEozJ4nLVr7nxCNqJKDP2U5htsSJlD3UNKC2dMomiO+wXsmbuFwMErhSp5jLbH8VxxTUq
ZAdDolmoVXtiZzjppfBadePKOmbIHRKdiB1royDkow0EtYLyvui6giSF1Ho3G3wkxmk9HOMVNu72
iCIRvU3806d+9DIdV83I3q4IJ1DWs7z/dQpJFYQmi/h00UKMJ6fKfndZeoI+hHnD3jBVyAwXJaQx
axyVOIGpZvxQDf3Yvxdhy1SRVibXiDK2/GdIMLRQlyCqWNhATc9m9igbj8Y75jXufwtbSua5lyyu
bneyJj16U1RoPVm2oP253Z8Gpj0rOO6L5Z7qGEr9hB7zHDotAZJBAWhit/g63qZN29udQHjH0NVX
FNXIMURhu7G5GKEFMl/2/e4C2h7tkj7JDdK/ZMsAvc0zCmag8IljVQwDuVIY9vN+NOdnyBbyKFqc
0kVjxoyk8CsNCtYGxm4CyK3vJyKdkVCSNRdl2DdY+JAJbUk8tsHOlTyWv5qzXGkT8RoyMRvMIWo6
8QdqT2PAsiCfO0bNiBd3tRtV2Cmbf1pOAiB+VY27aRrJRgX2HXHVMlbLHfDYlvvMNnxH7CQCTRma
/N4hwHwBDMqCxDC1//cB3HlFUoxA4h3pLNB9o67z+R2DlUYl4HV9WveSsUYMTDOWRTL5KTGfVvPc
absg/3NGLywrsXYBSZdGLY18tCyTZGIesQrI5qc0el2Ca3NNL0QiJhlwYHPmOyttvvV6iJu/LoCB
5QuXFnQ8ty+Oq7xM27CGxWf+4bhmIHoU2SOquQvGHkGxOCUipST9FDMGviqIlpgNdBDJh7O2LF3X
3xqwRHfw8NX5YE0YInCwksCgbf7xLh1vOAWweckXgDtrCDIn+ZzmUFeYpGkUrTFmPcC1S2YU295w
YJ0Nar3ZLkUMcPqpBEDnVy2iWLRkRY0mJDMG5LYwVz84bFJSB4nUU9t+XOusvqiI7LgQkUZfwE48
TGQy2gDsd/hBitBRI1ePPP+qXt5q15Dl6DCg+U4sq//uQs5gx7/nGwb6elYAj/RR+syxxmTEYpI2
ix9FZj6VZzjmsej4DWP5UinOb4ETKRZ1IapxE2Fgwpxuv98Itrz0ZTdXVIcTft1wj8p4z8zQE3IK
AdQfHxoy6DOuVc6EoKlcsnoe4TBkpwsZxFN2RvzDPzGzi9Px9OD23CT0m2KOAtfKZggM90rGd2XD
XQ8X+2Nm0QO/PODD3J6NzwnlouYRnR2Po4xYhIbQNmZUl5Oi+xtCTYT5Pq8GhgGlZatcfXYpN+Dp
l++gqKvCUl5mM0HkYRYhJmxm6laF97BtjnWG1yUP0IjZvhZmxkejA/OR4QhQ6tlGf/7NpQGQDli0
BKui7ZlF11c4pp8DIOBBejE+xdkjJ34NcbmAG0v5KXKN89xI10E7FaDd3T6sfsFhZbQu7U97bjj4
fgVDMExc2QTj0Ah95rtgW7E8EmiNSCTMXoEALECahuvPl8wt3M6z1ceYI1CSW2fYbc2K8zwe4W9B
kKvHeP6VhBwyzXj7g06Cr0NQO54AJC5a8RUtkgsjQEZr2vS7+WicURzBcYNt1rcJhfK+ZM22tjPg
IHqfK+4Gbv/6VR16rM9uhGXllLp6251bAtpt/p3HyJlTOKDVOsLeO/RAKgCBh6LDJyG9OpHcTVKp
wCmE8oLiJ6nEXTjSaYgUO5sdxSTyJJABg3Gij3GygbSiZXGcRX+kXXg1YDmcstqjdKGdJ679c1+I
JUoL785iOOLp3OcOVTA/+0W9Ch27FeuVuQeRRuCQzLRRk1kc6z5CqYrAQtB5XDuFWqX64NalMYPQ
yDPFTBxpdCbsKSL2EocxdUzqXCuOK6MK16Wt+R1CXut833t1iioA2c4K3z3GRU2wz/pKnIbUh74N
lydRhDRsr2aEfuVSXFZKiTtDXAIWaCpfqdzTIe9Xr1Ogm2EtcRALsq5MRsROwcQeMdKMzqvaiG19
gnXwuKXSdwz6Tn4uUZ6mpPftP4Z3fJrjOuOHRtFAmpAFyCbsxlve9T7vRojISiGsRvqGjfrwCJaG
rch/89H+0JJTf7oxS2F7A/sauM66CTYwPCCKUDxgU8le/SJHuajL63bsiD1qkVjfPbtubLXUBHU/
/x63SDmDRZnSrrszv61RHbIQoS3N6Sx+OCYoJJvL/KSREJm7ZgZ74oZyajmF5dMlQNRlh5FDiecd
OOQnkt10e8Pq1bEAXoCAJOFTBcD4u3+varpLzTtAp2HcJCaIbRqxfSnJqEDXGOHdtFhPwErfBe0C
xI2iI8CN5TXSOmboMWLsmOz+C2fvVIlVd/3Tz857WmHSkNAmh42Qn6oC8EG6aIRkxPN+VyrVcuXa
uIRLoCVClAy3x9kyV9hansaxk2WPhYoCwON9pUYKLMgpLgCetyKJzMTHWJ14si9vPoX0AItzOnzI
9zK51Er1/CwsmVLA3Ly3FYEJOcYHEV90ptnIw+pEamgf/UUCL+pcdqXEkdlA/XUg2wS4074f2/bX
d+cx9BrgSb034GbnrXpdFhTRVvfmwtIaz+ZJrh2ZxarAZKifl1eyHUHdCjkNnHLnAH/oOmJWP0+H
+XCgxxwbfgWoh44e576qEC2wW51NpbWKZjJiROeNXhtf2vv8RYpY6VYM5Psj2HJ22GHwoBXchbzB
JH/3AqT8M0wC4oY/gPHLwX7CdM0CKLNa7fKKDMM+9rAPUIRHRN9Nowx3Nm+dM2u+jAbVMTR0p3tK
MvzNOKrx6+2PLxxmk9vUv7vM8qX5AEtIwgTKjNOQtEtl05Ps7j4i0/pU0Bx7+BDv2iiAjCrTWDX6
zfGKdblAf/jdbxW359sNrDr+Or4l+EK5jkRzWqhQ9RYH9j1Y1KUE77bMzmcTM7SfJKZaquZr3oRK
K1IaZf+lfZhJm46k811qDo4LXcLm5PJjiEf5T14dYh/qQLnRPWoKSoWo88tlSjFnc31rQ4VFIeJZ
y4+gPpFZQNyOBwjVlFN4BwKkAOFbMQlvimrAzX+RRhoAM//3VklKjwmPzZQTM/1VRkDg5vYNyewG
T3yrxL2vKTKEDk3SR5Em0drlGYDGHxDoVRUKr0wb6DfaE8t4IwVcEsrRM3YG3JhITDai2edwF0ry
aHmSWtgieR36vZW2uPGc1Hwnvdd9B/kkHa5H94SaiARABQJ9RYfSrYm2jGD9rnWjQzLRosR9b34z
3TiPwMT2QQ9pogdxGF2ph8kVIe6llMTMJOlT3/a9eTqX1RVetdlHLa796yXNsn6GDQd7fYi2sTdI
4aGrBHRhtAWXttqc1nt6XXNY4QHSAEX5/wOTKvGx/XNgG85bVtkpUm4p6pnTB3jyvyN+wp+riERu
sQJ9os7AqmojZX+AmXpkUxRLa3zWJ29Ls2zr3eCWU72P0131xmnSdTQSpnI23dq4VW61ce/nWVDW
CsMIXSU71e07qY+Yx43p9W7QZ2rEHu/kGdhBaQ0rYw65YEAQeQ1FLkJS3ZqfojA2EM64DICcheq/
XFtBFnkSSkXNu1ps1KaKSLy5jAWnMCKd2zNwwUVcleYN/lHfjhlOCn4WIpy/gdjxoZST4/UWcBb/
X2MvEPCoPxzitHo/UkisYCpEm5acCTAjo4/cPcRs0lWIcJjebggeSf0USTgfYYs/wmpDDcKxBTK4
XMvkp+Lax2hZyZBzKC3G+aYJWr32J8+UV2yOJEI3Zt9q9ELF6TmjO2TrXg7AiTFQ75E3Eu5WDNaW
HG8BVtlgCWflEIlwxh36koHtoCfpI+Pm640f1jAhe1TwNcAG3ewwkSVR5FQgPMxkudRRu9oFeATN
Mq4T2k7mV8V2zMiOTtRSGtFb9t08qn+t7uUaqQY5OqdpDwbqJV3CBqRtySjzYfbf5YeT0tCTW1iI
uJQZ+4WOhxrZhz4xDQ9ssaJMwiYELd5iNkfO/LQIqFaCij+8BLUgLnU0sptcIu/Ytyc2/cM3b+IJ
QhugXcISXljQ9kdQrmch0qsBql11O03/beAvUbn6CjHT5dV4N3Z3Qb3HHiNTuyDNghqdNR+mSEDq
Sw/T2Nvf6CYS69ge8wlVfKtbTTCJu7AbLbnzeMrCP3Nkgab3XD1XmcTmlC/Ots0dQuFG62b84kIP
YPPfabR/8tNTXCb4z7pcpvQPGVLJTbsVsSwaAktknl+IxFLb/HMRzPKVZr99/L0V5ancehN9+dNe
xfWvaYVZeyake/U7AyhEqggPqtsL9wcaYM3/ZPSEfdsW8aThN47p1bquji4nl649Vs3W0DSEUMqc
DLailXe1++DzA73LHItAvNlf27YCnmMSJ1eGoSflgrtjgdN8IjjUaL1UxlRr+wJDU6KjdhcckAk2
XzepcjrWe94591U9DPRir2b18gG3agivt9xluVQ3YFHUW2s8+ExhMBWw+OWt+d7NmKtiHbyG6yPu
JOIzqBh5NNKNMI2qCK6ktFyJ5XkIePTYnc2WBR04wKGsHx5FGlbLT+0k6zk864A7OsD9ZKeFIXCi
nSmZCZhnyrbWmpwcZ9fJYyuz9n+MUHwsFye5PARlFzETclhXgHKVpsZHIh1GZQhaWdrm05UaSKN0
dxQkyZLdH8XSBGx5I9i7dcFKAxc31rlAUfHW6DxvIlaraSc7IaIXVl7ePhg3xtT01ifa5/Co4xzp
ZHI9bT7rnusnPbgT5lMah+mvp9X7xBtCOEvdKY349F3JMps2YffZadp8+lJbvTRLcAggN2XATsEa
5cnhcO0Qh+IH/nFmalOW1a6xGzim8UyEDVtF/EX/i/KTVquyCBlN8jf/H45BVG2UXdvF29+Ofj9J
YAcd+5rM8H/AlTVLYD3NW7gN3KhBm4f7S39YtnCzn3ql/RuN81PjJ+y/cmonsXn60xz09UkijYqN
DZTt7arP8jAjHAzRR8eDI/OrYHGSuGkFNN6EdTyVUqt7UfCQ1tJuJNBypgs6D1vT0CM6Hh28Zl+Q
JMf2q72s4Kx8+SM8V2Cu2+D5yD1uH/QehO4Bl/wBQqYTpoo0uxNY/epf+91TtShcFaC0B946tB4R
CWFrP9s1uy6yE/XWZCbcabH26rxxWpHsCso+VuazukqfiycwhSN6Be9dKeoLNZBhFadL4NgJeNAK
zSbH0FMS9V7HwNzvhqyVi2wgvAQq3WSfVALfvNWTmcqymQlQDOTarF+hg2I3k28+ZW60u40m7Ivn
JVJOrfdgQh6qqNC4ETsdE1r2hcwlwyN7LxnZvg3njmEJ+jqEyZuVDgRUK71aNPpvwcN9XhtU82jn
tZyRyLzg4mWRfuTBQBm2IPNVZyLMW5j8AK4zc6KKwArk+I97I2PT4e/Fnh7wI0O4HT/A6QY8fVJ1
I+QWZdqsDYoknb0Tpn0RPVvc6CRp9YadHf/BQpxEIVI8DMyS4ttubibOtZsqpXaF37wk1+TgnyVE
OP0SmAlr7+SCUdy+G6g1Nk3+aw1W6VgoYcWAUFmyp7kYIcmppsNkCB4OLma9Tr8nyhVvIrm4Fcbi
o1UsHkeV9UhQcrJeuyaMr13bBeoDWzNU7kCYTm7BbRafHxv6TC2RiV5bGWRIrn9grWWi+0PZaFA4
vh1nYn/gYHPoau8ouRY/JManZ8rmIupY9RA76PauBi/ybZMA1vC9OL1blAT16YvHtVOHeLZjI1BO
SqBSzaPTn2/gZGF9HRSp9DKHcTGN5Q8Sfugfa7jKc5uDvJSV0WDQn2X4S/BjsM5tH+6SkU0ccZZI
yn4IRaBOc4RETssCHpeneh8eiDG/+q6W1f//uO1rjh6wkwaPGaWUoBguiZjZMCTQblHeREQsaZSP
zqtDrKsSAc815zH2j5SKct7GujHHa+cLtXhq1nXvVRVPqyP7JktFdzMH4+R/XQGyEfqMtZMv1lP0
bFJca67d9IH8n0lEbMO8UzlKzHKhUwmVpBWxrg2iQqSYqF0ogFnmGRVlGfZUu5hHjfkhjGAtreDc
MWbIAzVLGYkVDiQXBj3dnPkYwV2MRVt9n1l1uKHGmwRPZ8ujO2Z1mlgXLVGgAyIuOazXIg1FFTsj
yYtu+4Yijq1Vuzvaex5To4XdIqLlfXpTXWuRo83KRLP/5E8BKW1O4c35P7Yvmpjmr/p1DFeaNR34
sjesoBSEVGSCk7Bhsal/3EFoQYVS5OPn5A+QIS4HaV7Y44xqoWdu0oBONo6cx5SquzSZw4dWfuvU
iepzlNz5lYx1wBiIMG3SvabP3Uyzu+9ENF0hfsJjlnZWmBebXh1ISErCgtzA39HFgJfVMkV9GUNq
6DBATCze7yyQazQPM74Gt1Vg/y1Fk0KaTxmMQplT6nQcxaPu/bjGZzbEzC6CnW7vvY2ZJQmRD8In
asFnGVbvzwbJ3J91WgTscS+meO4uFYnzh6EktfqALvH729tkENt8eN5EONloGoT3nf6suPF6l2g/
uuqLE4egvjmsJ7oMKmfxSmSxz+DGVXwtPpXTqnjvbEJX9iaLoUTDqkHCBY3rShfeZj6o6ubDltVf
fTomWW8OkI4/DuSqRA9kmaV2l7m8gI9yfVMNhzVocOCkgz5AjjT5vhPMgu67uTO42epDwfJ0Ne+X
kCpcJK2X6Ye1+xh+4M0v0MbSv/s+cksfHnED/toK1lE9wQZsrtU0mZBQlHzj1N21MY1rqpLsh3C2
1l5c2w0IpZijgLl7wf2ZdWxb5xSwTKcR8zBV76oSVAR8779UealwwzWfPpGzBrJT6gvp8GaL2/9J
wr0er4XCoGRUP5eYuyWeaIiRCnw1eq2WEVALJw/0pjHT/vbZMEioxfSXiPYsNOYhZcZtEXvakt7/
5g6iTm1+rrGnpqmbhDCcr+GfR1/M3Lf57BXEcGCYlaPsU29hxT9Obm3s0d5yVlF5R9LvB9x/u2ao
OdH6rBesl2d/PRE2BaSbFHLrlAPw6hG/f9NJUfbiKGmQYfumpXKmYl13eDXgOCy+NWNDTfjsi3En
CCR6N2CkI2ubpCzZ5zs1sm1iY9/14Jem8bmaHkLikh3AWJksLPsxI+ALoVoAKy/hTsxaFbIkiBTH
yk5OI3hXPp2Oh8A/DHSKw+ps/h91LAacEgyv6XSceQPWfeQXtV/BG/TXuJcmXFdkhv+lMtBURQ4+
p4O/BonF6IooFCyJQsadMX3j1GiNgRVEzPZhw937Q0RNsOJihuSgSKdbM0CPIy1JZ83gasPDEnuo
G52GoNWtNtol+IzhMKy93S5MxNz0iKHtzJsrB8YGGYT54L/hV1PB6mqi2W0OPJz6/iZWnGmAUgR+
/HOsws5MfAcuGnk5kHr07HWdbMWLAQjeYAtnc4JouhMnpeAORaC3lMsYZ3mr/ZfeQjp+BWNmdPhB
fivWsrrudBQ8PiiHFxKTuYjWUVthz+mWL3Eutf/rn9tUtxaiF/FbHLqIUtTC5Zxxk1ieen926o93
/ouiSOUxA8+z7TXMLyG5wbfMjk9bQ88wqH1ZySM7H8lWc51lyVXo1h0nBZHLKFQMC6gNGo0aohxr
CMRFFyLUg6y0vpVuO2sQgtUL955Z9Dp5lj7Pj1gn10+sIvNfRgosunaFyplm2KcdiB2hpoI1/N7a
KTBH66fs59BXwRNVADhGe85Gn9VUZE2ojGOk3pTxmrz0nQdwLCcbJkgKAhxZucYTozNWbCMnBPpp
aKFrSvTbKKVMEEwwdz9CRMAB+EZeH2i4lHT7fORWWq3gkryoLJWRy9w65eQL1AiYYOn2K8H4Crxt
/pBmUZE0wGBoHiMOJ7AUllFpfMvcIcy5E/fbTP6v4rxL25zV4EbT8PntwOXkMuP8/dOiwm/qU5sE
/ThZVF2qWL/D3ajkHFAG3TjR0dgtdaQi5mQiRebJMKDW3C+0S7SQb32ZvYNAETnl7TcfajDcEw+D
ZOFmiOT/redYVWXL4BUT5tL2F4t1ZQQmUuQc2Ur6mZh+X2ih0EjOePybIYtpiaRnQt3Prq3oH9/M
BFr4qg/C1TGhYVGSW1Q9kKFlGgrUsJttwZ5fKV3lXmHAJ/237HQzTutOr2R5/Www9RFcSySjD9uN
ETrWVBOjLzDBT7qQqyUBjrOEBs4qaxV+Zzd9KoemyjFMUEnFUXf3hw1wMKdgFLj0tuF8ouujSq65
ykbsmJNXgyphbDrXbEz+ZkVaj556rzxujS0lJ8s7xJTaKR3at13FZ0ZDs7hzX+mOPIywc6cvqcuu
KRtbfuEw9i4lMHnpu+juKFDVIfcft5hmtKAiurnCHrhvfkkongpRNepgLEhqjUJ18DYDKX/umrFH
pWerMMce8P1ZosP9kOb6xy2PZnXPCPYkBqgv8wDBf/ajYMwIxg/XGMZb+mH6Usj5BZyQBrK4bPaI
t4l1JtrLnhSnctjML5o27NKc43haNmfs0O/VfuixYW1rpxbgcwFQFzFNGV8l6eP+OxIuM/Lyd1LP
tfQU1PSuIjs5BGEwtdJ+jhvBiO+QpS4nbfP4lIN3JWpnWpeAfn7yDtAb253JKNDAdRZu18E01mTV
KALwtAw4B6gLKa/CcVfOdIBdLCd2jJ73qa9hzVdvkLSJ/6hzrtlizQStsHOPqQA4ar0cY56xcw7u
X09Q9x06mLGUHo68eDt7G24mPSeTNLTnH/PwU+jlI0wA5VJJprpYhOMtaup2f8DRsci05944puSs
ROhvO1Mo1s+Ot6v/qhMFRFj/RC+WG87jwGA5ufwoJa4gQOIZESvesfj976EaYNiJaWJ7zYYCFw/F
bZLaqYh4x0ChAOuC2KHIJHI4BrRrFrVhB/fZSVo1a4yPf3pSMeIJWQe74eATcgf0REeFLK8WD604
gVC3DO1zBDpICHJiE5WWRnfvaPofC+BHEYV8YRH2huRNbzaD9kfJMi5NZL4nbaIR19kC9Sh1Pp1o
79KDVL2EhG77HbmBegBeNQ2MpiNrQPL5c078Peflr1RgcLeAaxW5fgpB62o5O2TFPN4fAUi/NnuA
hlNRv199/JkKjUGx9XkWYZWCRCY9LGeyGW23jSDSzr9ciVm2nDw18OqKZU3bDEcjiC3GO5IxZzka
zs3usyeZ5raZMp9OQWBb6YUBb0ZckIsaZd07BHONR4eRhyBWu3Eg6HPhZKhImeBc3hA8uPNIIewU
K5tjysqvm2DrtUcYF4rj2MbDZsNbVn5G2pOsbv3RlOlJUXygxGrnQUXj3l9NNq88Kw5rNlhz2dgN
9+iZEm2/NQwpGRIQZbgw3SF6nT7JG8V3K0OlIGI8EwK4J9U0qh3iUunyWuqntyUyS/h9EV6iMwRZ
YEszNo/0spEpKAowMDFIIu2umgRS8SO+wLB3P1nexU5hKTNlHrruff6YyjgQ05vln19l7ugorA4j
eonDbQq/JgD0+VNCeDttLobsWXoiTiHi1oiGTetVrV+RD5OAtxNqJKyENAuzoo76JtloJ3q44OS9
2SE8ZlOuwVfzfSUMBNd45gcs9hqSv5RC7+9rcghcOAYPhIm32zB2PzB9TqS0AIHD2IMIRK3FDfHC
0lKN2i9EoZQ9KanqZk2JwzyZhBF6HY59ZZ/SUmi7q9VcGi1Q2uXliE92aTXTy/c78p8anytrqJRb
Sbgo6Zx35X/F34lzbMNBMy2vb4CdteUXMpxIizWNm0z95SIkL3TWT1P48fDokEM9d/NYk53mlNGm
zrjAD38wZwgfGcgjdDAtLl9yTy5CraAHXKwSo0dyLf91bbVLOyTIfgGgJNyBqQT3DK6OBVjR4kKV
MJVnTKS9X1im/kJARAGQO7RGU5tFgtkka7QB3yMQQrfZWSW6EtcDn8QB5bhmSsGl9x4H04b1lA3a
7tp4pJc3gAkQ/2mdbA0h5dgmDgJneY6nIgIxOrpq2NcwmfVMHjfQ/A68xZGF2IK1K4k3p1bVEUWT
lkY1FvqkzwMtaeylucv2OSlZ+RNDBqoTePt30pZxytGPu9smo0OHp8CiR9nJPORpELO3hV9Jh0Jy
s/qadUDR2unI65QmClhaR+R08DGARKCMBdjHqlE+nQBJH0cIM8Hk3KWSRZ6oj8BsgsDjqDAVCMgZ
PHsLLMhxAHzTmSUbiikEOMBiJi5b7Az3y+fkAxSNRurTxo49djmN/iWv4LBxa1lCyx+ULnrLLXUH
EKssVUiF8CfL6bWZKVt+x15yAROIMs5uX36hIlGCKyqdSFMLHeUErqTMgganJ80wIvbmrYr/9RYU
u8kHniy2RtN5jttWRHtvLIKADEUtVMcHagGrFIQdXKTrMV465hCkKVrlc0H/kjG+mxtHVNJbIclU
SHduJcCmF/cthpr8+9xVl+WlxFPPMzPw0ha4Sfq/Fcw/VkKvmDqWp4GvCpfRKvDldez+OUwfjv57
K3I/v892iZzkjDb+ykERYdCtUDwLSyn2kA72mhsEb+oGmwl9CsPUEDARwKDg/mKVb51lsrrS/E2o
gZS+YtFT+kAHc+FWRUcBLv4Q8iYYJD2V96NH9G7xL2B+H7uyMTv7qBet1Nq6+HRuc21U5UZXNxG7
hDJneeU7LUJUkrsMis6srBdWlrnZ2fnYv3w0eJi5PffJFu2lpnvkh1A41xCl2EtOgx/icCoLuC25
1/i6z9UYAEZJVJGtb7FeMQwmx2J50k2ItlhywH+zlun9D4rwQt+b3det32uldidvzme/IlzSA2CQ
qkYFlOMGW1mwnGXq6ubLM6D9nyg+Rp0GdnJ+hhCh2kIGcUkLhgrTU/1OFhQ/kG6ld3C066FqK0Dt
Qs6fKUcoO3ptSwYvdsC8ZFg55iJ6CFB1HCsoDbR0x9VqU/MS6dkTksXTReNCHppSMNcu5XzPYg5t
vfyK3RIBGYn1YgE87EYbAkXxF2AT8q3YAJXlLg0vclp3VckW25qDTKI8IXZveXYv7ijJzaGaGqhW
3urLQWHZ3v9FY77BcFgpZrkcaOunmFm+3dd/H/nJ3AkOr5GvE7qb0aT8mW4U52h6FNviIYMzsBDf
Kzio0j4WR8fKbn2SnkNxdZ+iPYT3KJJ66/iwyYSSxv1IC0plV10SQl1E41IJnWqK/ni/e/tFmtPm
gyfsqXoS8XdEUCm/pxpn/GEf5mZ8JEtyzluViTdpDbrEJmRX0N89SSVrr0LTmD28x+mBFAy7iDIx
jaWNY1ioSG9PJTNoSYhw3jUJGPkQwCPjJzsRZFk2aULuEdzcVuUb95GgOPLLO7vvF638hg7pHAc/
UmzodwO/DOAM7nRMqzYWDZfyReYACfzrr7yEnw62OftiocnVYIELXOa8lRk5qY7XRS1ZImjOWBMF
hCfxOWWoQRlsjSUPBFSk7xjfly0UtkwqlabG9hmoeszLNT8cul3IhjkenS/PlQ4C4wxLEotN/xbv
TSkJLTCu5zSmN8VzEzgCf61aGS0Gk0MVxf+nB4MByQyiv5hrkSMEWqyz+XyauEr649iQVjbiPm8b
l3KOWfX0nCMk1iO7E1Xu1lM3+rc7SbOruETTF0d+oaov81zaxGNln0cgJeZNH18S23iHw0seHO2t
zxZzPHpVEsh6oJ6BxHEcQHSPUScKtXwqAevATMZMQJOOivzFnrW6LBZYI8TC6TjlLbVkVZhnbUg5
g8ghhLBI7YcWmcL/6Ih+qYIwx8Ui2GgwBCJlMpicCCWS8NgDeXoZpV723LiF9b7oJbJwyxI/4jJf
RJVZWs56lWNW7g2JC9gyJVKegGn6wMIp8xVxze3qQi5qCdkSAmNM92Jf8+H/OQvOMDrSX25gF4WC
mczpmAt4BgXR5vOHxdXrA5AAdxru0Nt+NW+8xjEskcC6SDllerD7/MLHt2vGWQRhsvCdnpq7edYh
Kh1v5IYMzMH5VIIB8l6K5W061x5iLp+CIL3VNBUg85XIPBBB8LacQ6HGQ6BxhOINK2w3yFVYJyTv
vHSzIHletJiNFNHmrq/xPDJyaXh9urTXVRWv2zDXGoCxPq6ko/25PuWhYeBM177/zLCTElMTLZXh
sWopNoscviTJ4WD2vBTyWZOarTIO8PHMEgorde5qN3vos+X55nROxvFwQS4QgQ3dZhh2vP0MmSaZ
uOWZyBAFvh3MoHAPm5mKM2ZLqgrTrMC/+EGxD8YXQXMaq8LDT+J9tjh9yWEE5NRDMZpxRdDYhyoQ
oPM+qqH2HePziH+RBx3709j2cd6fDTCdmOa3mW2PAna6Ul08IWCuWkQBW1xndHpf7ncyWtw2CL4O
/qWRRGk9Tu8Mu1akqb5dlUzvzmTBtifs7Y459/PalyDJIyWPvVTwKxrbMLb7JV34NE+wwuauOYC2
NVli/tTQCzZ8tSPLnTGW9pHZ+OF53dFI5ZAJyYF8mvGIzyfa1u+ZZeBJhyqH6T2LN90otgrZXySv
+00q5G0X7VhHpND6YaUbz2+dnrNgViPBnXbLoJam7Y8taPuGaWCV4IpGA3ia2CSFI9XzCpO/C64j
y09nDV5v+u6LFK+x9W7hb2rFfB748bRXDTJzgzRHwcEqY1VHMdTBF7PsoIJNm/RQ3JmUZO0+XT2X
yn4hqDxUYBvoq0dTT9X9ofaNvGCxqUlLHWrjFS0OM1Nd6vKr8o3OWJPliPyDvKIUxqdt7AnI/Hqx
xUPFJWne+T31a8RjZKhSNUUzj3C1LVO+l9Vu9t0Hm5F5bWU6c8UW8K3oQHDaAVF1aH8kXbAfOptA
IgcgWNyG0PI6i5INlm1isrd4ACdpQlQUHRwynZ+4lVaOAujZMOJMI2wntSktr0KrLfD96PT40EBz
qsAnCxMXGUeYN0mEOJP2XjnwEv7dhRCOmxApteNA2I5VWSu52YpX/0o12U/HC4e7RZjk3peX3bbo
j/sJalZ6bMU/u1RrV+fpdRO71vC0VFbp4xyQhBzU7Q883AlaBcu+po2KTUW7ntyCK/qtGaU1UQn3
iXy9QYR335XbMzYeali/iXTkIda31ip+t8uFy0CeBvnzcfRgTp8KxMwjJJwvlIV50UT+pJqILa3Y
89e6Xip3YVHnerYlQNLzFXINTT9Df49kMbZpXVqJkiiRXgs5oFmZh7w0peE9PEJE1XbOTEqRGhDV
fhK6su3pVbU1R4+HlFBDAC8tD9Dgt88O2gNog7bBGnt7wkEgKkc9jkPPJvfkZcbNiNde9b7ejOcc
jshHHeRXaZ3j9alASx6JamZcryL68XDXQAlI+3Eo/RZcB/EHseV8bwvgom+ZIEQqmXz3CXLQCsFr
3nV2obhM3rCHNinFklfIfbhpdSa3J++hgcy/uf9E/CIWe9/F+bj3OLFcyk+6IlXzUNGyA1KYDPky
8+cIFtKzfITRqXzPAeo6iGAOxTrxxeN0F+Rl1yShB8tkf5aUaykSfRkzi3tDCRnybzyQ3xlQfngZ
QDaDsqXWCbyU9UXfqyKQigeD8S+jNo/AFwuRUUqqNgqObgQr3uoCZ/6R/0vrdC+QtVxyuOdh1y35
cX7mHuUo4305M8LXrpbJdJG1rlyCA1fS76OYV3aCbLUG/XtoP1YFz1q+HcK2ogkDorwy2GDJAnF1
TtPkNMtVPphpgMJWxNcPT0BxaI2uWVQmWO8zBihrn2aLz55A/nOWD4nUoNQ907KAvo1JA+nSJysl
oXpuKQIOfVyvkqQI19lCKndC7PY233knr0EGf4YroEQri0L3HiAIkYH0M6Ef/orQCVr2/u7qkfkK
/4gSc+Z2HIe055Rs1l1P2nCK9xCguoxYO5zw9U5wMRQJUfsLYNG+RKIQQD353o/OLBDh1Jf/r2tq
S/K1zg3zcCjYa/wy7u24f2hQFmMFTFCZJi/Byf1mWj6OonMPq11Q1/g9dXHZ4GRCK/TiUYb987Qs
+zUi8HitbkFl/r6eBjymp5JjYKHOfnhZ4XrBlScvrdtEJw5xxYefQlKtSgS8/jw9QRHrakX3fk5q
bZ0DyxXGAT28C6i/lOfzPNXSGQxpvPZ8qd3+O8Krzp2gs+2jKQbECdyHNUfcttTdq2l8qf+wCjps
+buI/po3SylnW83S/0LjlU2vB/4YkwhA2XIipppAFovA5qCle6psgL66o5PZeWl1BXa09qXoGF3W
081sVSZajEkezYh+kIfFjCKIK1QarG87AQg1ib1MptpIIIjHNljc1udchuXKlQcJTWu/Ksk+DXEF
jaek4/jJ33XdD+L7o1SpQll83A2Puu2uUg8Ruo1umueNKOX78oRkOyo5/P8gjBfzvcCrBiFKCM7f
4SRYyy6WYxFvRFOZv8o+kV5F2uS9qliT8heR16UQb5E8FbSq9s3GIcWR0rUihIdmW6V5U4kHtP+9
u7zA0nrxggg0BW6qjDFk+nTkbYR6MkTqc8/Lz87+wy75iaYq+z31jOX5F8P0N9Pw+pfxAPHXrQyq
ZWP2WYsrWwdf8lbLKczGFPAY7zWhXK097WuvYKlsmkHgPETvCQe2qz97eBYvk8KoJwT+LTfWS15t
wNDkTI4Y6nR/9SahWB3lzr9DKnw2yYJQweljrkN83hawPWgMWf8r0ust+r/xCcw/5Viy7NiT295u
nkQSAHrIjjmJnhwvTO4oVLFFeUPHZRvXb9vH0fXZdlDI3fhTFeOf2CwI9HxtUNAI4/cfJiKnTfH7
kSqq4iUNe/QE+mzGalUk2vymo2a57l3z79cRUmYKqRgy6o5toAuqGpvbtkJyjKwRzAv3JjTfxtk+
KDD4xgvO5gBqkJFrdgguPqwifs69IK12FlPyXFVurq7gjqtcy4uXNDU0qVRFhx17gXVA0bnyNcKz
8KYhp7MHNlPU4vYB/goa4Nw4aTPJC4T7+87b9rTOoNoAcUr7npJoE/yPz3Ot5HJ27Br+tf2B3Hsz
bPkKaUB8MG4P6jS+T5FBFC4SbmhnU18oMFZDKfxAf3BX+baQdsoUzTD7oToZfxTCy1B6+7+y5290
NdcSouRpg4Sp6XxAz5FYVZ8ltSJBo+bFDoRW8achJqxMYhoa6gOLW7Yr0or6dwBXL7Q59J/+Xr4s
jq/UJlKVBIlr03+r070tN/BzyFQ4gifMwFgI/5QpSAs32qwbhPSHJAY6wPoTWyCrAu8hzqmMz6Z9
xlxYXRrxhi/vg6QfvmAzvC7fMt2E+6L+xnr7zCAuUBkN3I6rx9lGwKi9WBWMOo8iiXaV+mRDRKnC
5wb0oTfmgNZsKcDIlBXknamr+iyCiN24Q05OSQu3arXu61ioi+d1IrUCP3rwHI2z0r+CRx0HK39b
mRmVsr21ivx5QwdjNa7kX5bSSGM3SFkZpk3o54AEBd2CVRuBNuJY9+DYUuD1z8FHqkHhi0piSqL1
CeAPfJv7+mKgInGZ1yN/ZYFxtRXbVD85LolXjy/AAOfuERmiR/IjO9RGH42+2aIGinV7OQ1ZNyrs
gn7RwKPJvod9C1Hgyip34FdeqhwC5QNvhNVr2UVSAC/XyX7MwDWzg+4/CmGbbAnXsajQVAAuUhVa
08ZmHnZYGbWoMISVdY5zHDlFvNvjbam9xyYGj7QbQicNbPXr84mw3y1cinAimaysny4RIy+Rkyd2
Mx82CRDn/2DF7bH4ddCOeFncEoSP+uZWNTbsB4Lq0CsHxsW2rjkG6N+YQfLwNIl1dp+mL7OdSfLq
nPohBHK115IxGHhnezq4Crt9IfXJOQGZFmSbgCKqkMImUqn9xb+8/Un0isOMBCGA2SDw7z0l32UH
pAnXcUc4EgXMptYJ0VyJJss0C/bDk2CTi3D6Psm3+6zVjx7SZ0/9PwxELjW1sky0NAMu5ydvmBuy
b+RUC3/uw9P3Yx9I6sMzVo6rbmmyEOBxx4AjFdNwm7pR7KsB7asM5oRjIBtWkbhbXomo/0XuVmi4
yaZUqpPJ8ioAn3NLekKCM5Cp1eA+JxscVR58/gQrxvtRXjRB229LrboUP/0XhPiR9A2g0uDvKLL3
J6gx/Yr1GTYwpN/Nih+dyOcX/KjgaqPV3J6ms3C4NaCBPRDi7S9kh8vOQZvVQkgbQK6EMLh2yxGX
oDS5sumjXO2dfSrq4aK+g0s3VC+UW+UWZ9eoPnK6nNqUsHjamxy62Fwxm9a4rSFulXd1uHiIaHPF
AXDuh+5LX6CACgdPdb9i1/1YKmZGgx+Yp0QSi1vO2uvax89YZ9Gj76Z8sVOR4cjoTOq4RKzEAanM
fIP/2fqavzwJm65VL+QFC/fKbjQ15VtlxFh2jKo8a5ZAXwlFjS2f3NQaUxMfG40kFAPkxxRH/HyE
avBQrczJvGiDYRXmQ+RanpBwDt0w4K8OUXgsz8eH3av/FAph9SkDpw234ohLJeZBgtVUxVwYLxmN
be5NX3lX8NrWEU5ojkzOVIJdHD9s3I2cMcget76FDLNYP7Lf49kpY/bGny4LxV81myAzrLj2z5iR
Juas36FM8X9Ju+qAIoH2naj1jC8tZxZ+uMzv7eZMpR6Z4Xp3qs9P9cyJyrYQBJFja/C0/Grlke2q
iU2emyZ0lMderxNDxY8ua//TADJLs9mSQAoRDG0a4/ZoQ6QGlHGkEHW/D/EPeg83RBJL832rmU5D
0Jzt4MYTEDfJzJyBZg6d/l/eFdqNI1+/CMSRN4uGD8HSQlO1+bRiqqQ3AKo/MmyRY61XhiYVpqeq
VI+hNDcVfy44Z/7r25zqesqtmMGbfLF4gK99wpMPwV4Zz4cg9WV/YFUXu+Ayo6GkTbnTUsHS5Aaa
o1BdIw7Xqs5/M+EhenG9hu8FK61sTNsgKEr5G4N0KrhZjdL94+cCEUB6un3Iyc5VsBf58uuU4HUb
2aOcHXWB6NrZgLd8pV1zmyTJYeYSlkHbGoxzv+GDQJf/XEALE6WYIyy9immL81D2VmhkeOSnzwV5
WZe+sdq8+AFWUpS2lZmmNzWLhqhz3tUScGAzX0qM9HJCE2RFFcEXupL6k07UlFEvVbtXEBvay8jS
6mRcpgavC6nApX0PeK+TvXT4niTi8ulpMfhq568b8eWKNN08ijzrOzXvkMkP/QXJKUz/Oa+i5opn
ViXKvu6hDDRTn8usZ4ya4BRCbFnuAC8s9TzC8y3j8ak+4K0geiWxlmWyPcAmHeIgh3dXscsrWxla
YUzdn5tkQIHMHK9GlfzmhdplF39ihySkRFartSJgG+g6pAbuwLxFtNLw2UytKfyn4FXd3PSEJ9Dz
b72usJnANGZJMdKX1Txld4S0neqGSNiWIj2ocIJ2MdjlGfJM0blUkvNsDhn7MHenCh7tKDIk0x66
e4+41O2RjNyH9b4cz20d+ofpGCoKDqM5DITnne3OShAQcz38J98hGjKcXqDQcnVb3ZdaZAoEPjsv
AY1kqe560G+J/yP/w8Tl19LVmSpzxEeTf9tA3kkXHhNi8r9suqRcfp8oJL0GPujXkaxtCvbbmyG6
tOh9ewTN2Mdy27fnhKcDMTaHZKYM3urzylYjugYmDZdF8HiG9oU6qyhvmgUSMm2SYLwOFi/d6Zr1
bwhxRHiUpQz42HQigjBO4LydoHjIkvkPUufkBleFfzmQeh0KWJEhf2I2IRrzP7n1l5H/TrTIuv9R
tWxQIViZTXevFHt7qKuXQ4oOfYL08mKI1TR8xbkzk0HFo9FzY1Q1eWvnZ5hSasMlo0DrjotNiP8+
x6ZeeuDkeRrBx+QX1MmjNMREzcwraRdzRkk3+SnQXWAuAopY1QYOaEPtYcv61iHjDynULj22VGW8
xbzkRDqtfAdyaTLmyknXqjRtb4lIFLGNzG0t3ZA435+L/FhtJ1cHgL0bwPfGO94DrzloCCU7oqqq
s2WzfW/OdDc2ME/eyMO8uJYVcIbIe1VKEq4zBcR2puqPZRXzjHTX38inSnTH8sl5Nxe764ZiVGFR
/XKzF5szVpm/lybj+RCHwZihRPvl9NJYMQWZAXotTi7wddCxHxo8c4lSIJeEDKogVp8kCYQB9egf
0u/1++PRdWR8NLWD9DbbCq6AoQahV9ln3P3zAftHAVtmQjFzrPQdeMLaug8PJlu7JccIoJl/oViE
4rEzdyda5iUVKCQHoS/QPog+/WeJXR56q32LGxUog47yKogorcZFcQrPkNxaFON7rly8Fr82+m8H
D6LOetJANF0ra3q9oPVdC56rvMyanLurmrzvktkZahr285TrRMk1ttQEtFUnkmON6gpt3MKmLElc
O7sOLWU/mHyMMGkLQC5SEjbitdnVeqtmqMrOtLWehIVWx2Mmg7dWRDbAQHtLnqPuwUe+qg/gDJ/A
/9bJgqU298WpiHXuFmeuxTNXKyqjLMEZwmdPX8zPrR3Ra1JNfLcHWPPZi8R/NQZ1f/91V7zaIOF9
V2aMWOvaiTqnxHLiitYOkfXSafpzyhEJdudagrb3YW4D8MPvUBWIQT1ds6mxzYsGK3bLoZjGEseS
Tfx0UULZHUJp3KDAdIhPGcmOt2kdm4q98sHv4t159Hr/+KoCrQiBXqnTNTqFq6U+AAyhhuDz93fG
FTPZWbPaos/JBdCGde7cutAMuNsQn1hfFvSE7cUfaORM5iY8H7LuIM+CUwflz5fB0AIg2KoGdXfx
RuF9wtC13Tyo+Mc9LRvtsNNzkDdJqc/njMudobH9lnwYiKkKGOD4HOehgIG5ePuQrHDvaBouFBLQ
I4bea7hdLBu/holZ81w2Z/5WxvCeFgvFmQWqx2LIZG4+Wku0V/gA2V1ca6KYqOU2jQ+M6x66apCe
hY6snQhUL7Wxa7GJgZIMWvqQfFw5lX4yP7jG0Ls66lYrGgTI8UavQ/wuCXvcA0Wgx5MIKkMwTxts
XI5JVMz0SNFfQe/Fs6qJIMFX863o2sldKuC0ffkvgUyR212AUy+RXHJEAcqTd4RjlyxQoJ8L4df9
R1gDr19yJ3Qa2cDmnhxxCn3kow4mIiRmCSW2t7ZppsG5yuSB7wxdBUiUb//Bq5Ig3uaGzhqfkSWv
/D6t7fhI8XqH4gmiyC+BejPLtPlsMfyV394tTBXBnElqaF97pK1ZUiJoFRg6OMe8TWwqjB0616g9
u5LAhhuJKp8qPdPzSgNiiohI6YcKDc1bC1RtavW7G2YbLhqWP4WloY1CreaVMkx1sc1+cm8vvx7P
23ac+5WxFZP5KrRFR1MV6kuPjuQiC8z8zXlb44ITjKvEqgsvCYwWzYH0Vs2rO0gaLme7M8wd83Z4
I+KiNJcQadDeTYcYL+hMVN4JQ1lquQU6a/YeFV8EfZObJVQonZKrMdCxq3J/iMPFe07G7qO0oFmd
zxnycDMWrjEriSxKHXsHen0P6EGxq8VJ4LGNH5PjzVBiKhegokNkPqgRIBH0IXHHIEbNWqoKfVXP
VJTv/ARzo1tSF3EEDI1Y0OErDDBgr0QRD1/ruE+8KyABaPvNc7f7CTIc7q4kvkMojsBPkHIgA2Pn
pnD6yP///Q+k+Qxx87fCh+ClSTouzvu1UtA04hQyzvvLSHYFxO4MgLrSLQNw+ywk8glZb8QRudVy
Z9Lxmacy4B2UCT5hNtvsr8luPl4DsVx5vPWP6WvWslH21Zij6XEZoRTDKMWNCX8+WmBqCkssNpRn
CnH9WgzRNMKV9f5D62a3LvYoidzPdcZ63jhHu+0HxXvKBiMBhABpLse27td94PA5/iVM0G5aTg7z
K7N0m2kqQGnBAYPfE9J7wup5DL3M1SKvBm1s+OtGgprGokruUZ5OgOKTXVv2IQKukLZCfmSA38Uy
y2Pmb+DNhBNnOKQlUeJFRk4C8ba4h7FLOcQi+YJC3fHkj1No5C6i3Y75sklthukoBx2W/KerO5sF
PwGdTodAhxaLZ3UL7Y645dNToPU1tZSghQ1bvUmlWPrBecf8iC7nQY5YKWEtuWgrB6XTyJbs2nPC
Rjwx0fvWwrWhuNEcNsZuFtbU3hrid7HRXUNoZU8QqVxoTSGi2fsnPeda8ytQEIfOiyxuQqtFrRU+
TBd2KX+3DDStbRigIXyu1rBSXzCW+p0OsMPZ+3VUppDPhnyhzd4V0i5LtqhGEjGkCfZpfU+3TxIm
tWZoxogn1LMs59IyW0ClJqMg2kS77N+DIqsT2lBypcQXHXThgkzfi0n+317UizSedPqwYzhI8dFc
RKJd1InJGfrEq1n6+CBG2fhIJne4wDSOxkynHD4irnnyokUnt8UIe1PKR3jDvfXoF/0GSuAbmWzR
6YU/dqK+sUP5u66uV3K08fSdkjvXyvOtf5F5Eb6dNWG1tdGxvWfkX7yHDOmt6xoNQb88dIwOH6Pe
/5KJqLjR7D0b01yR+yWIG2Jst8PeHiPfg3jqPh8m/UZ6Z+RfaSs4nOKi8LsThMyln3w0aR/Eh4wt
BppYjy1sSscU2bn07wiub5z0XFzjxVCgJyzF95z6DaZjJtvPLngqM0UC+NYilsWuwg1FWUCYIpo+
IcuhTFwwj38ZRKCx0ZQiNCHvTS2QDbBuo7/1J0Z1BspKn+NRvsvjz9+UDAmpcS3m41q+GtBywncO
z/MLSripFtplcHLDMNV/g9PkvGEnCla/8P1m/A+xPqocCVOVysXll4okPllxRZljyCn+PV1U8/e6
D+ZeRZ64O0yQK7XL2Vkc/RWOLNePfFntT2r/uAUznH+FC+BWgqQRIB0KD0mbErmqDzlKxNUloOZU
dxb5lg803GSgU5UnWYE6o4SiJXDYgu8B0jGq3Y8ijvxCxHzBajMK0TJ0OMv0Im54h+QhKL3Mej95
Ac69ZsiIX7XP02gfmAreqL6e3fXI1gWJSlIT2e8+7NEBBdQzKSdymO0UFL/u7R42hR9+WSUp0ZBS
4Hfv2e3mG161dj4I3XvE7zUjolFHCv+IYz5Dl7isFBu+tNB+dVsvaO7Rh969xjc76oJ/Ai0bkpYY
saC2ev+48FJ1fw/vlbAhF5FwDmIA+IV2JFpJ/pnRdkHlu7TblToiOxx01NE1DMui7YQ3gE617fhd
sNdY21jWIvZQUgWTfuA2sjb/EKhq7E1pHIgp5ygFRutU23cCFT3A16va2779SyCEExIIIQtrVeA1
QFG5CdnMqwEJQN2z8XnsbZsK9s+XIPvdCh9gP1vO926vLVLjMEuOtPXuENuwmyeC4XoVwvGZEIkg
loo2ZbpgX6Jql19MHdwzQ9xbHugkiqgz205QJH/Afm38N48owWOlcfRra7bTmE+gT4HtS69Hajhu
VXjmNl7rJx8e7QaxmMcelo7dObOwO67NuH1AsxgPEEw2dThXDWPWD8kCTVh9NiG5UJZ3xfDOETJ2
q0GlDuliEC/o96BbPcDInGhgyJNzdNzY45fXqS/KM16IAbwZdy1KNRLceoaGLrIK5nXv9+7eHjzV
lCxKJESnxUv9bU+TXM5dM+N5/oBIFJIH8q/ooXbL+3atC7RW10pAmeyuwSrFdjbgplscihEqw9DQ
kOWG5T15TfeoELaN04tPdDeyrg7ht7ENcCA1qK2zpK64s/TeHn87VjtpGXOMYsm322JMQOkrcYPA
29rQCeUtl8SGuru73kbztOw46nNsMLiHmKWccJQ8qSM+WNdgWtA4RVa2TwDcUWXg8VSJS315Odbs
Dvl259RGIKhxg0Zq8XDpMXCZoNb+GP0NFSaMa68t8Y2EcZb1IbNDmh5l/5mDL+yeaNL+hoo9GH31
OG+QroWcaCOpVS8wU9A9XUg+ZxA4/Ciusr4w48HUX2EG+1PWzvfVyDIGZk8ahPeP4qgvUa0mgeG9
xa44B2N79bwOz+SpeU8uvJnoooeoqSOQS3ZaGCwqWfH0VAKXFOzpqcn8sLhaoFmYIqnv3NihfEio
CswpwslyPiHqQK/RGcdVNTiHyGo49/eizSdGpUDbjDC9v3JxBRA1FCM8bBBfaS9/oqWsgPWZ/leK
XtdVPyxNS4ZnOmabRsJ8QBHOsKLqK1E3Qv1/joiRNJXYW1Hxj+dobsfJZEb6KRrlpVN47nvWidby
iVcPdsc4kOAIR1nNk3ZfEHNXp/0/AD33DQaoiZHvcSgAwZ6Rwa0isjIdChAUqVYT0nVxTJB8LRO/
mZCnwTyi+n7czkBCeVivtSwGt8o3d+Gvk9bLdg0kKNymEhSOKjFB4KxZHIygxtLBdMhIraQNNTUo
o91ekIj+W/rTBTinMNpmKNlCaw31tpd88op/IXTZFMpO03yHqb+3JivWCiCIu3J+qO7OjglaJ75w
S0RoftxEmM5D1xt80fEwTDUeKqR1Wq/XGxwz/16MzCjlqo0v8X7u+ppBUSgnli3uC4yHCy1DHosd
hFlhLkopTloZ0v8Ug9JtwkijX7IlXLnAGWupiNPknnX8b1l/4l3j2tsX6+9x2/x0COaKKflcXD/+
KzjPdK+SOZvMVMeBQ/y1oEw1XHRb90ZxdCaftuxXqCH7XbLk2Ho4Q/W7ppGsmb1T8/1vXK6ELv3c
LnpA8i9Nzn4J7+49sXZdDMfkH12BcAcWoZIxpcu7bRVkCHn4e3Yszt1M1/4djymYSyiY6ifD6D6X
FXYjgPxuW4ecKi+zMBoFzo9fs8CNLsIbv9nJ5iI7dDNJizb0w2pv3I+hIPtA/y7YsnNNZeZnrsEM
ffn8Da7heBZCaGcQGF1l5mUR0wCXDXOxjUK1dNDa5J7nNuwJwEXduPDGWelfWWpOzdCKymkcJzG3
YhEfmfBH3G+E7ihCjrR6+EN4PwuZh11Qip/Y57cBlg4zemYNgrbPPsdppNHMhDFZi5HJ4TxT9Bbb
xsOUWJLNLfY4AwUmJkP0jNvjSX0wTEwQszMeHfVpA5jd0yqfqMO146H29ugoEZGsnfgCIirgAEvG
XpwDmX7AQKFYBoElyr/DqyHXWZPra9YiNuBKJ9OBRL9ra496ZO2FHx4sMHF17p168SNvBApoYz8D
5QE8XYZFU9NoKxzObHDEuUsdH0jPXON/OVFi4sYof284BUkevjs9XYRzSoTwkxYRPraN+JQV1ear
PSmUcK06ctJVeObf1Ibehy7xhf7BJQn8tNgjuPOqZ+WKzAvl7p4DBDm18YEWf9Hy8BHygeDKsLWv
QKa9iVjKQDZ+qqyskyRLxtc/My8V12cDQpPTJP4Tg9p9bT1ekLt1FAn9uKu+xmleModMjDopHdQi
4w4LRYvdg0OpRFWJZOuzxaXXyjhOwZLdvUVMJesdYWObffu7gR0jeF6yN+1H+7gS4IgpH9rg+dmM
GkihliOzXKijNoK6yzYZ0IZn5nXre5+kb1IuAfW8OLJSCLjj+dAk2b0winZDITINrMDJf8OjrnFf
kSHMfO9vEyZcy18grbYA1llZdDp7XcIJz6KFmqm16f7mPUZLQSwYuGx6QM8QInV7YdzXPhvney6I
KbByL6tjuEpc86kzdwZfOgyUwgoGkiil2OLhl9oYXOQ3qws4CFTSYkUF0OfpY8eZGhgtPAA9gEkn
cZeyJA0HHpJQICkpS02xyTLylrdwlgoZqg6l625EmN74aD97/Pfou08hRH+0K5VuLujY7FtAT+3J
DSOrhbCQ3NXwwdbh4TsMZR9susfa29brAMsawFrO4FcXBEIn++bqosWfMeWaHXkCMcvPg1K7Ei8a
4KxYQkvv5K2W4Yxbc0rDDt7fUxI/PvufVbiGiUW1a81j4WFC0mDQknyLqJ782hYtMnwQrOYN9TB8
RYeiRDcWWawckvJcrpkUM/NG/jBQEMjJl1b+aNmWGzl0KH7GRXigTqUWnJtL3wIl1JT507o+jYXp
UGo096F4fcKGFlDkiwFE1z9hvQLitPnPeu/tQBWSYy9W4RCI1+bRsh62nVO/1bj6ZswZ+tq0toYu
prEHr9aU5zq7J3gPwV9TIOjz/9Yie7wd1yBpBVgGcXD/ZJsUsr0b96H3P1avEh9jMqYZA0pZ6N8c
282pnqKEt5Tg+iROpQtEOgLkP7EOxT26Pntz+wUXfDyI8FLrsDSkfz2IjuLsd5uteJEIlLuvgWGv
g2TI+VUCdTWgYudxumj0/Jctri5LDCZsPe5RPcMaaz4Fb0PxW1gv1zWRanrBZY3iPgom/8HY+W8i
9p/9z7Z0KkeLckNIxn1aDHT3r6unQqGYw+wQ/ggQMe5OfWh9V66CvP88BwaBL4wcjuTx0RGDZtur
PIoRj7UfrN4IVygDhubbiqSk6KoOnEZLK2KB63UvlKpezUdnqzuvCZNQw0FrYz1RMUfAU47TYqX+
QrhfTsGIKeQ06XiVapHIouj/09Lsdu70zc/g0PS1/S2Y7Ce0ssH/FoSNAFlH2oGh3E9v8OPE/rTS
SGrNETjXX97O3OAnWlDXLE5Xd2D7y4R7LLftaD0jbZ/ZgrfxZJ16ym6ZoUdMaPlTwa97mUjwDkoV
pKO86cAuO4TFxATR97AEDU0I/OBkPIRBabkBDcVrIi6bDcc0HhTpM+mMUvElb5OZfxnqQn4mwHKG
Ir96nTyCuerBJZnhxVr2ZZg1ZCGGNyAAcfff1M7or9fxLs52GyMjX1usCfxh/v+G8haiySsTWYf1
lkQdUYSq4mCeX20Uq83xEMw/iPwEyXXoRuueD9WwDBJKewQyMGN/6F41e6PNiFZWILa22aMSfZ/o
LbjZUTLvXsMnbnLrUCzjO+TU758KLv2VeT1IhvqQpr1s2YiV2LR8qTaOT6eD04NAkyIQXAfeM4ie
SoQH1Rkkw0fuRr60bhf9c+2PR6OGh1ZXUVLaFiUek+bI7ZrNxt+jzGP9ouwx4OnxPHiZpLSUW+B0
WA1XjED/haySZ7XDBCWgYrWRhIdbJ7fnSJKOgvVHUDm3YPjZw09NQ1j7+Ka84V5Tl/5G4sArCjyJ
gnzI1oBgO6JGrYaXgZbJxK1BBs/P1hydPyebTTMlOmFZxxCIkaNpd4sz/LWLj+tYbqYt96ARCMdT
KAk9BXt7NvntZJq9igZERpuu3MazybWUBYjcW1J3p9D4TWbPLW8b/Gvb88rg0/PSZRLzCvdLYCvr
X2vExnjOWHGOTRizFqr7xTKdH+XvcIsBBAS82i0fXIJTE4Dhpphyi3FzTNtf3hf2kaE9PFJtR7nY
JmCg00dXu/gnZEJxdV1ezhOjTTAqJVPV1xByHyrUU87wCppYB4imgrGZINtNJjcBsys+IQGhpZQh
YbcR3duTZ74B+bUEuECNI/Js3oC0NDbhEK3YmIlKn68Q7moNztEBg7hdT1xSECtatyRUD/bE3+hZ
siENqCQU6rUG2guCkI/BJNBFDB2cKKvx6Dr+YFtzUvIZuFP5DBDqmSaBuiiNPdroqUOFw88v+Lxd
75sxAsPVlEBdjhI34hojHNwCEwEuxn3riAJGC4bD4ehc5+N8dBu/UNITxVtDMH2sxVWqaF2PDmHe
sr2LzJ29gIfvpC3SW+HJ/x1Mopq6r9m7GOIUvzy+g6RksnfazbFACqcQC+e6eBU969SdDRlRRLYl
ftzyLQulvXhq0SHsQfKUwCTKl7hAt4pfGl2rY4QVzZzxfSkUD/WbyO3ET2G9ZhLlWSrFwcK+EdUJ
Po34/Lmz6c7/NKGlYBalGQstzG+1svRTgdl7D2wGoaw4FQOZDYo+O/ScDiQVBeUlQ4z75mV9N/5F
bzi3QeXRByiSJ3sWkOrsxYfxwahXbkxYgE9Z87L8u2iWltSVcmrpn+66QO8XA+6s0s+41XT4lXfN
d5nVOmZonUbeleINti6g7+iDrtMvImBJuNtkBNTBkxBo5HQh7HImuG0N9VnJelpODdUH/t6/p4Ze
1yozKtpRHWKHSQRB/rvRxkYEAht+LufpE2rWwdN1yZ1Lhl1G2zO6LUqvIFFD23z4XvWNZ7p80krY
MlMi4p17F5FFqRu4p+WVsVaKqXK1IQWhxOcMCoTAXIR3j3SJOWkmyDM5hRpPmGdl/WCvsrHhKFgj
nmxSvdRTJRXVrgwcWK64u5Imw/wHuzbzUiy6dGQdZRr1+LFuVluTE8G9AK9oCSgSHZ3TkK6Sue46
NUlxL2Ky87UsTEuHNbxjzZ1aO+l/KPy4gVirzljhiVfXcdPHreRnWDmSMg9etAtkW8rL89sYnJzD
UnCS08Zaitey/9aqPw2Io/+fzTLbJNYJs0VgFd0XoLjCqlGo16SCMg1ptzhVoBhzUOeZi79BBpsl
vbktcANQh3CLEepv5GC2DJsgDsIcce7yDjbNorr51v9dUu/Cp7oEN9UycsecBKtZaILKtRoC0LW5
1mrZ+4tF+Bs8HO8Oz8mEW75FaE7xT+LXvF0UlhaGTvG1SmJsogJ2ibSvoJq94qLDoB8GWpW3N8Rh
QfuU/30BD87ooUJAz3qJxBQ5up4IpInLc1kjK7EvvOcOPC9BtEiC3VqMhGp9aPCY1UCT0gOtIgTN
lQJEFrTFAiQIylt226gtg0uS7tbLmHWPIw+YyOL/u2R/JT0Dj8jIjh5vLtd62jPfwwGzDn9MU992
FufXDSkr7okEHeRSmpiR+0WQUK4T0Fw3Niiw/yqDn+xZGGEFjhtyo34xT/spgbhHAxQZ8z/KoxIC
dMB2TGrlJWHGqLElfKbxn//HsINR9u4PynaTjsSifv5rO4q9f23yQAc1CDzrXbI8IzR1GrC7x1H5
fSljjCjya9Rs3CqgPEL51OmVtRIPXg5yeTnKUYZLsp+uW+dhgHHzo9gDjnnQCqGLhT1Qed7cP8Ir
1DH4Fo+LNXBJH5tB55faI7gzcST8ogNLUNd+kAtImb8JYU2VQPz9tcw3UcTwMkKUcA8iALWVQ7p+
mmzZEWQwH0qwq8gxywp3E3e+MAiaAxjbMK1OLNoKxGKTXD7M20yEs1/hUfl9zsqYUReRPn2o+R+Z
xrbwNrF88/vKHS0slWQsYF9d43yPbVy0MAra/y5IHnj2cksyi+ruz7aion8FhE20rZtaoMJMKdLF
g+rEZeaZI1DJI99Pfit3eogYj8Z9ahNRiPlUWtuly0OUl+4fSbrm0KrskYdsx2VL3Fws/nh+70za
sXOXIfnhRzsAuWT60TtwZSGG+mtzpIf5tkUQeu4oECwwzkp5YEv3NXPBzhg0d2FFp2kR/UseNip5
nZ08IXvLroTu0wyknuBycmkK2+/zPfymn5uRmSGw8EbsworNsRPbb48P/rh8k7jsEmK3OlrX2+eP
hy5M3WxlfJD7CQSTBoBa0ItQacqDZemOUWFJ3VI4IcsrpKtZqAM+rt+CV9Xd46bOnSyXaTFEOlUH
ah0C4em1CVSdn0SbH2L1pK65m1yTPeFEuOdSH6RAH61AXY+eTXlYZeGNXvT1uxkAriHAsQ7vpdOm
mLzKAbbpHAHj267SN7Y4dbBe50Bo/1FzZH8yAmz6EXpY8nmIEI+YxChSKWohXTuNU6Zi4HBEpV4U
ulq8NzsFvEZ20rQHkWG64wUQUY1t+tdmol3ujrj5+qRIBl4GBs3bzZTdBXnnNxzkzninXgBMkiOD
kU+6/tR0ieYYT8cp5UCZVAs7hBIfBOSUAp8zqzH8m7Imb/MKGzfUUIxe/CMcDqNBb98KKMqhuOLO
vi7/hIegIxYtHnbOsvNIOHgS+y1YspZg/0kbgmJNuuSP+koaZwXppRyuiORUtkSGm1YCscLz55Ec
K2RLYSKJa9JEnPW5RMibII0NYiZvea1fWYWYlnWKlvW9tjWb+jDMuGZLsJQVqKCoXOPAcT8rZo2+
Lr/8OX5PIKzlof7vlaXgThn2WXrdS6sH1NYNTVl7s3dM3w2uoKE74XXrGA7HKFTvdNjU61WPmzko
YJWMMXRUQeZx2BWO6cENgBpOVXGLdzLG9dlr2+MT+hvcNhbjIoo3i7wvjQv3FHe1hi/DLq+tdCOB
EwUG+/tnCjZ31Yc4Pmt8uQBBXHRgk4vw/7UPwGLxFVmpL6HvOgSjQE4PS+bZXf8BU0MRhxPICIHt
Cl419d5qt+bEKE8PozbIg+dCfFLjCfn0lyZXx4wHYiRH0j33OxqUfbVgpKp6dGlAqHgyubn6b6vT
sD4uuloDBhbOLt4rlRiHEOqBZWaaXqGFvPyavfmopbAsV5hPyAZSi76eGB2XMwWE4zSJZ7QYu4zS
ylVDphp/y50dAs6hA1e3lRgaqKYwzFbK9HhZoZ37Wt3upWU5MRy0wttHECGZ7N3/wK5rmM4g3JEK
Nia4uD+6MJYf4gyTJMnx2yZAyipEy1pbZeTRgNiWFAZqcnVmCKCQqMWAZOkruTY5HKt7UEsZwkPz
WlPevG1zaToIrN/XoTHeyG307YLyC4V8pzSzccHa/o1hVL1hn6p8ghbALZwDSPbTgSP+5a784I18
bSpvEZ3dtVwQLsw8KjlXrXjrFmFqWCeigegaYwCgod+PpDylhRXRe+X96C/K8CdXoPQ8fqqMMPaN
OBecwggbTywR6rf4I2jaIctW4O25p8Gcq/jiAuYviQU1O4Qm3W5iu3jhJJ9ehe+eOOpt37xfdx7s
/NV670EvQXFMzgVY83fsZh4s1RsO8gslqHgE7R+i8Q/S62XOYyywCIF6IMeeFStVHiQwdTmu7Z1C
w+YxxFUp5A4x5avP/+03tlD1zBqdMc60IDM5obMZ4SsZrut8u/Za+NqBLKb8twMfpKT60o4zIQaw
/pOiEP8XPDWD9iuNSkvQD8zyyUjELD9aJRJHN0PtpVGnNK4huPiLVrje7kIeDDlsiCIP+TLG5G9B
xREtaIoJbAeLkHeAmqMI574N6Ud1UcPjOh3n+mV+ZX3ZYPuj0+PKTQ+0V5HK8fnpWGk5cH6cmT0/
zEQaVxyRE/xQIaE2hS65V6VdjnuGD41uAdiso7PI0NwyXJYFihpqXP6sOdafXUOWb8Af5d8r+ypI
vUSnDDazm0Rp+62a3hUeAi/w2b1dHlBp6KUSgVPzEepWCZPXo4i5qHcuC7ygIy/U92PKqGgGylD1
yARqHjqlHWLHPDcN6EgB+Wo4pWcLuAo7/6brvf/xUGAPm3iSatxqZvl2Euqf9ANzyLTQQNR24vpo
uzurF4ITAbFO6iop4CY+1SBrhqXbWS55mQEE9jnrGrJBg6e2ts1KhxW0GCDyVp3eIKlPCYEO08BC
D1ru9lta9hAMSmvHzzjhjWfIBSGav/LYGyQxmWBeXTd2xjTtO7tNzXEDQoCM6EtuJPEXZkTYo+H7
X9XjshCLwy2+wy0khrbVfcuK1IeoZmgi8BuKnL4wiWLArJxGeepDV1TAz1UynW4xViEVFTuhytur
LG5BF33EkrS9MAOdnUPy2DrC2a6WSzkm7auiVLxOz6zFL2Rs0Q+QXfkb3P0e66JyS1vDAfsz1ASM
ysFR7hhRoaHx3Y7Gvv35vHMtj3NbpK6byNjUQ0bIZc86qKDTl/I/WkDq1ykt4cMvrsWguGwMbj7c
lOpgjJSQcxKMQe4dHNltGrSAjU1fvWZGxdbvem03J9gSfxfjtFXyVwb9dTi8cjvxpZNTQEV3rTcb
pbfTkIonBA4f+EQafHNlIKk2Mbm8VB79OnDpFbQiyw9usvGgWwC4OdD35vxHOESeaDaVkbZ3XjUa
HW/dotVw9ralHrWObYDvAjwG2fLRy6irMBNuK6RsBiDwH1r2zyfTnBnse22LYLxG65PiGqAEvprZ
/RqZB+q6bi5ra8wfCXZhXlM1SkYiVKE/ud/KrEbMMosDoLC4TGufKvMPmQPfbirahwWjgOWuTfr5
FTHQ+JQqy9EJuLZnv4QJyh/4E0mj2QfHDOM1S2CXjo1HqIscGugTIMsq10l5CNAM6EmooECBEcXm
ROHvtwpF74/kwCzYImdYyooksEccZ46CbjDpek2E2pywWTIfZcWkB+ePILCxqW5EmwZNEZ61irEV
AZxhia0zwgZF4PRQZbr78mZnyDaF3Kq31r1/FedSksVCvl65Ppkwdokj8T6QZ5GAhqFFkLM5n7Xy
n5YBppnuizq7bWKzkatrdNl0YKdJthYVPNZWCdoIojTEhV9Gy3f44lut3A5qyqtRI6Qkld9anaGg
D/ZH088JJuBIU4qf9JMjya3ayLeYQDYn4reO9WV6QXvtl+VIGBsfI/DxqmPS4n1MMNZVHjIja1M+
VB9k6AMmmS3+u+0iGnXzcWQBcH9ndzTBv2UQsD4p1QWgmvQ5LSbQhVn53XOSeoEp9IcFSq0aqwwM
oWEfTsu8CTxxMye8xhYnKlK6Y5NSq1zvuZJLe8lKNaYnGb+1zu7b+ipnSC1w0sWuTx2YCE8BiFzQ
siBt3EkFL7lQi7dL8oLpMD7VcdOidk33OYdrBjBemYUJ3gds3LJWay39hjaj/YnTvhNtSRd0tXZ1
sV+IVj3nii2vSY7YS/iNLT4JJCDF+T8IpcBK5lBNmjsNzPU/V9h/6/KuPiiFdi4TbRPXUpsZnJMC
gC+Hc34qqtlcVMhq+c9VZroH9s60TwH7fPBefxvKohtDpeXGY9AH1oqVf/3nKeWE8Bdq0LDgPCv7
ykyt4FolvwwrmCGrwwtcR0wmkV4vBBn7PEWNqCHG8lU4ZY+EULUSZrRxnDLnx6E7qOKuD9e+Jqyz
J6rzVtBmiyyH7Qah2LQcOYV2bLtE5am5CDMg8McLIjn0SNA6juLr/+VPDqBdtfAtOGnj5AyCpOsD
c2ZgFQiLdIb1f0kI5RGsQn/nLb/L9XIUtYHcWkBaUSjSPoFx/yeEqkO850sz/o/eBljbdBXMeiak
96qe4Loj4U6kz1UPbjy3Tu6gY9bStKDdW/UJuQNDPAz1YEivVVurrHfH52Dr00CdQmwsHJSpRWGf
+hMN2Mv0h9fobLpgunfPrPI/4aTXXxnoSVpq6Qk8NkPvz+1124/LSofv1wsxc9r/J3CAPrzs+1Ni
QXWrUTIOkl4kvHiplusOpfvRqhTTxG9laJFLDTZ3O5vG6gPAi45lNlDreuwdKwhAtC7LLWS4E3E/
327c8NyPF+aliE0T8OHRqzDmiayTq/LHSiFnBt3n43mGu6iezH3FfAlbmClyBoL5JrGZbaJEwyxS
v4iP0KQ8GJzYq9giSVlDmnfcmo++IO4ngus70XWc/iSPpNPHNyS/39kRg2LuPzUdhlQRLbbOvI6g
Z2pMtMN6YKQfSb0kMhPMmTXKUSV8Ave3Lny1BXgZ3ZG4Q2rqTzfFWK1i9W0a58J+rLOGtJPDQZXF
4DmtSKs85QBxI+qfwk1wT142wjbGO3JGakpUCFFzIVWONxkgp+L8sNp4d86yqIgcBnvSADdj8rSA
eN8W0DICcc6XSVxSJ30a0CsAR2a9iXjm0zHrsbdZnJUAbk4Xjo2IxolKrGT2eDJPppfeF5qPw7FT
0vGcImY1n8M5UlgJjJEseYVTRSzj/c1CcA5juMwMsi3wZJVG2nucH0H9mwkmamhU8AEXK1Fdydma
r4PgNkVkPqPV3vPrWVqno+tRVw2amO0F4ROw46+m8izgS/6PhfSzwCyRb324gmFLMLcYP42r4u58
3RBeyoCLcF0aKA1qNhFIB57XytDxbjkg0szOp481m21TESc57tmxYh4CUnr1KQBwNUTKZe4lXj+W
vhsBZlTlyXyhbLEzxnVtkwaBjrGA584vVBVvEBGCz/QfgKcpCcKHDZVm42FSV+69mmL/mdczwHPF
BFCA2zSXb0UZQCBiBv6p4xFJR1hACHIsGwqOiiwrIq3vH6sK5fKbYwVkLfEUWECfg3lik3YjgExb
F8Ba/aMJcdVm+cozJndWIgxQZOKlYbMtEpEJYzaQSznae7ZtJkELbcI5NQWWBRzGxA3fb4nga59y
B2mXCd3c2gsD7ZIT4AY5K78nP+5VQX+EWiVyK/L0QxikmaFRpyUh36xyGJAzWSnvM+mJCqA9l5Nk
2nN8ob06RLwsMz1pwmn5JLd13EAgUyEyH6yGf/aK8iSjBHDAITh/qZgmIoWX6n5uglBJ/+gKc7ZJ
qx+4D0Y2D7YNfmDxKVG3yUBvWGc3fsNykEg79DjKG8MUO/Jn2Waq4ef8aMPSEl4iwF53CiyhW/uy
q8rlTsJ2WZpLzrjCKpUZ+aJzmF1J+q8psh/639Lu7K+yvMnfvnZRbLY8CqDLE2aY82RIGhJD8Q1Z
llqXqZmi9EkPvgqbzvvrQhvsggPp2Q9XPRaB/sweEk7SDy5AaDLXfk+RXPx6tLFRrvl8NApNGJ+p
Ejz8DC5L/jPBMbhka9Z7RHV2F2CTbtNV4UUnoM9CEbYD4h0rCJwiyYPqjDcKFk3yRvs84lpZHGeo
Mi4Gs3JRk/MKvqeILRJushPbvV1iBFxBrHkEK/8D78dbccTEc0nugukS1V9TutDoXV1q4L7BY1YH
XTmtpe5jzYNrlfJbX+ZAm2R4/+GieVesgRgskGKHC7QfUaavW3pxjRViTPvpSF//Ho9BFgT6qJMT
BodWKUN8M8o6g6NCtlzrN6hegabR+KcKfx+/tITt/8w8pOfnRtj4SP+KEwtOrICgCP1yyaEQLGC6
iTsjIKUK48QgJn5wGbYUqa6OdL68nxqzX7CHsxb1HfpFiSWTBQ8RazFKwQeGwyg1WDUoajslzeB2
CUE/l67fykN/PBzW82isbLd/KTaX/de4xnw7hxpdpBs4jn1sLrGPNH5sFgC/3Vka4qIohCB8ECXb
jZ8ouuRwnrSvr0arkQJAbBg1XAwbseWoBXYUfd4pEzhxd+sl6/aHNN96lFjAjKdcrcQI5vvNNVI1
go+1cJmyj5QW5w80OpUofFkLYZWwVOQfeDcqYAvNXFXWhExgP+HaiEtXrEAsGtCgANZjDlTvDRK3
yBl6GdOEosneGwkI0g4GR2DAO9MXbohkR6HIHziF5m+NFaJYr4oHgJC1DAgRjgfzjsWRBMsN1BDr
Z/UZZ5SKWLzKgJo8g0XENl35NeiP9wOruevt30HIr9rd9mGkF9JdH4kVM0PWh4W+jJXEXtzcqSot
H/RQp8H0MxmAJ9EWECmZUmWiKTuxikTiyjIc5FsmkSoU2+YOMnlsQrPk694q35uR2c0Ej8FrqEpt
FhOXGSzn1/lrwWDdtfxDqL5v2brnhGBKi6c5qqY09y7Z1H7j656UL3gRm+r+fcQ9exQGYl9UuMU0
ng4MDrpNYfFGnGsIKzN/icDYkFIfQ35CFFpKcWPEL5p4hLcPYztRmSLN1lwTlXHUkM/f6zuFxB4P
god52U/jKgOaJlqI0p/iQqtT1GrOg5ZmRvrFaegq4b3jjfR4SlxeNQArQTusA/y6ueh/CmA7PZIA
OLDGsYAFGfGWogTKivSMJK6wVfK74XB82C2ChWsDnXMKL/Pkx2HeLiu4xgOcI7f7j1KkZvEDGVX8
KlKSWnYtd2VJGZNoATX+Jx++3v34i+22GAykJDJDos4EYO7xgviMi9focN3uvRNmzJ+cDRUFYg1I
15Rb3l/GMik+cfbd2DIKQOnIJEYYgvh6CoYccrffWXQ9duwFZ+2XbrBRI4FEAMw90uUXCYH4fJOG
FFoWTMglAUaBwJyvf7bLXuSFntTZgcKgSxOlUcGnXB5kvRH1rjGJ+L4h7yG8EJ308B6eou56Cgq9
/rYD/cPm2jb9gaRMva2cROvLpzWCzMFylwvZJl4XARZkQY+5WXTLWe4c4snWHTNfuVN/zp5pfnSw
fhCm/DIU7oqvmVvIFtaZn4y8Iu7Cxm1g/t3WJ0gnR5DyXCyxPNX+daS+pEWy7yB9l/rtvz+BPHO2
NJDgc0127ne/uuyr5MnFU0dXmT1wzVCzJZaCVcGiWdJNlJo1kVHqY89v4xGQzKkvo40f27U0tM7b
k58geJxqAaHwQwKSQbM03ZJRsmIYgMShbR0JSwpBpemDrgcHKzzLkMTPafR6MNXAnz5Sqk56hrHw
m8Ck9Z3XqhUjyiFPglvEKjfQvBaKbkopESK+0HC9aFjSevCaNkTMrTTMwYuDldSf9i4cbfAI3ygE
NF4ZVZeCZ40TTgz28Gxa4eoJX33/awydgQOWmtCAhrAPDn3oAeycSG52SB1PEvAMdshcrBr/fJtg
BAJdruLbdGRq6N2fDmSCOAFoxBLCmcBvgIMOqhYVKDG0YZTFbLucbVmtl4I7nGVkfEe0XM4X+YLD
H/KHy59kyGwCaE5DvFMRJ7Ki8eQ88L1/qYkm+lUIJXJaBCEpEBGyladDxLM79JXDc8w1Vg8I0L9/
B7cUK6oNqUFdLOFAX3LyVZlRwGUN9HxsH4gtbvVeKvjXz6u5OATm+XFUTHoZHvkjfxjoAJ2Dx2UN
0hZ/rXtKIOCoSR9Ni5PpwdrwGJi40JUrYid1sxkm/JNg7W5WjehbeYkt6Yv7wni+ntYnzqEN3GXF
EuqxVchegxE86crHOD7q2Ky/o4Gu/gvkRi1EL8eYy5gqNkvXotHB0l02AV4oRc0DXYWcvpMKrOdf
/0vT40ZyjqpMzKpaqTSbt0P8Errn4xidwG0VJiAskIzP+AZijJYlLkr/NgJ8xaTCiz2/7Hpvn782
YnQjfywKOSGHlyikpPlClYdt157duUZf5C4cidbw/FB4HNI8KY0g1GYvErUNetROFBnUXALNigow
QdMd5B5LW+VryS0f+DF7uc2HRXI93jxW1zQrQhQOqixxlDRW53tRDrnNfQ8KWmB/JwOAWaRhWEXm
LoOVgTUp1wfAWx7N0xKVg4IrfRGKA7dZdJ7kiIwIYP1L6uBNrNByBPWI2qgHbUHv3sZhXkvby019
FcLozJ85yf235qncbSuMhB2alIO31Hp9NcKd62k7SojMAcKeBn3dc/SRWWTFl90BmIYItOMxqfNK
3yZLG8WXKsmEgZ0Q93IE0LCMgO+gxRRae7xOYCGnDRE3RQ2jrv7ZJpoalkXguvbgcE/0AxkDBCBl
NACFfa1IvwafGNVxjtoY0P3xABAgcDh5Gfa7+DdtCPgyw3eM5pm6ji95eto7cmCLjsxMBsxQDaum
G1p6hTge//2+W/KI62n+faND+9dLFRfF0QY/XoP0dkl2dtVJudiCLjT0tp/tpw6kWjDyD9pGsf3X
DRDW3g80fuvWN05iKYCjU9H9hH+F532B6wvCbv9DuKELxMNMjKpUAxP2DzCGL9F7TTFDLrzU6c5l
b02iQrp7lgu3Osjhu23xMO8jOs6RYV4l+jmKaB4aJlQrhfwss0ntDPoD07APMKVrlF2JcZNylVqc
zosZ7rEOfTazAO/5dDXr2Q8dauEUNlUtuuiFrwX5It72Hq0YHKmtnKAA1C+GU2DO3dHhDTTD24I7
Ku48ZiwJYkyr+ntS3c7L4wIWNm03ZVjBFpwcrCtZ3aP/iq37rQkBKm+VNLtr8zupXN8qRhYodgHn
rJ9vRuzDGOZDeqZ7pQpVPnUwT8DQrwhknFQKShXRB/kf1NvuXCabogXIkN+iyHk5BgSnx+vpM0vg
tOa/x3u8q2F3vMxd/bR8ZpcwUJyIcgKSLO/i0wwIuwWmh8HesKXkiEd7VDnNBe0LWU4XLekEFFKf
TwgbYcmfzGYMAv3Q+SVd5OicolLAXDXi2oVr0sUv6EDKQsPoBfQ9ScI4h+mv8l7eXA3rWQd0TAdj
T0u3djYcvMUGkpSTC1z5msv2ifCUPbIEO1esgq87kxqqoWPNWHxv3kpa7TpHjeKQoUK6k0LzqRBY
RqWcMD318dhq3JuV7VNMa+fRMJ67pwpsYw7gAmeDcvgFoDamo6vM4LM7szWLEekpQOA+VYsVHXLd
7IhobumDp9gKxrHxMT+GyT3ASAzB1Q5gnTE7euYYYTt4YNS5i/US+t+EFsqoKbPf4Yb5T7gbaR5P
X+0kKWPWfbwhAVmrLMebuFXbW8SheQlsKB0eao3ccsWfOAA9Okt0eQJBPhdzYGahKEJD8wWSc/r/
7eQdGONrf3kezGHq8RA9FNvCWLWzG/V69hrJ9J9kvdRBuX8mnJSqnaBDDJMadv/pcFJ84h4NnA0d
gHNdHam7UE2uitSvxDLtB+7bR5dGBlWV2hqQjxF4tNTvOuHSLajGPpsdLymzyMq3wuPZJKuXDGpn
F4duwh1CwFuLPfnuooxYKjxNuWugO3PCabqxVBl2TuDoaf9SrzE3oaTldVP+8D6ODAzAwkiayp8a
aua65y9ZM/nbdvJHtU72Qosot8btkf3ZpGM3MmB7nWpEZ3SKvGKAxgqXgBH/c5a3LBrf7Q5zXU/c
bnVXxL2HgxRatP1TKZYkmrTzY7A/Goknw8e0Tv6GLJEwIrgyn/LePu4hMLNcONMgIOzjAo+TRAL7
sC2nbOLw8W263QK3YmgpkChTUJ2K9pY2eMhL7YzUq4U86qpy9J7I95GkyYODG0prgnXIIs7Zg5U2
+oRs0FuP+zo5tnflXkbFgyQVuxfkF2LpXVj920BYpnE42OQzg0KYZHXKlwyexzWlxAcQk49gOPK/
62LnleLew9QkgSi0Vs82JOHW87xbtS77DrJGmOf9yu8TtmR7FAhSDi5E0fpxzWjjc3XKiLa/4j7r
XMvvH8dbcebflDPQ3cxUy9l2W5+jimUN98QBZ/PatI+mBrmnsGjW3R89FQfXXlZSD1kwqG9+ixk4
mQbqGSz5wY+8QtKHiHxzrDWIMTQpmIf7Kx2NRF7phoOPCRGq7Bklw2aSxzSs7DytZ/9s4vnwJcdq
jRv8E0c+GWy5xQFlGwEVfsJl430fD4mjis0GCrVdqUXE/E0fY11E/kuaomBATSCpOu43sN8oHoEN
lSDJzNljORCqG1bwdtqEa2CCMEwUzrF1WmzgrzLhlgDJIwdlo/WZ3QIEj6v38rGA40Ob+KKKmMPI
zLy640OZST/7kdZpF9EvxwgPhs4FswtaUWmsn3y8cH1mrCvCr5oLK51n+OdwUaaQZSoFdx3UrohZ
5IapW/cOSUkQdnL+7xKHnvwwurLpsknrxh7FS+6il7O4JPj4ZPW5dlkW5ogUpIjQMrftiVnesCfm
50TTIrVBOrzYKyW3A6aYWjmxFSwSbtJB6IwFxPWQdsu+cOGpMfB58GCwALQ9bc3qETQwo+p8qY/U
YV+Tz7Ulb+OFXoGkpwxEbsDKUCzgto7SLXMNmXI5x5FYgz6WkEsygbb4GPKt9CJrGpGfXlzmMZSp
Sm4pE3CrJhGZpeE1caJV1ESc+lD1rOoDBVEMBy1Lmm9dWA9j5XfFjyf8I7OjFcVN2NEaMJzdCtzX
0pU+TWmXGy/bX5jIl+cpFB76zKMa3byQA+oazpxc3W/PGpf2zueGcr6pCVC3iIxqBRRHzIxRuUjc
RKE64edQChKfaKMRhkWC8awAZv550+vArmWP8lfj+grwa+8NuGgUapI5BrtU7PAEPOGXQ7TIEoFE
E/g+zidWNPoGzVQeYgJS4b+ZBvW+a4eafVryZ6YbBTOR0RIOQmPMpvGyvW9sqPyGiRHMLBTw+310
faLl0AHpDTw0xoB3RtLp+zrZNjoU8Zm+YPdIvYr5GNs790AQdrmB7RM4ErsOAO3ePhSU2cmVnHOd
Q2a7aFZVZ/7vjSJyw/w+jyb4itDGke+fvMgbQvCIWvI+etrmQ1xqttxPpP/jdtmF9XMxSBNNhWrM
2HnVdIIX3kVk09VQSTkB1tPVrNDCS4Ffl1tcMgrvaaQl01Cc7utROBHVtfqtEKfIKlBjddsvR3Jo
1or9XWUcfCD5hYMDN6GdT0f4tt1ivqoae94tRMo+/oNweC/0UycFtRifdGajN+sOu46naq+oSiC2
lFnIZVOpJhESt/lREMj2T1AEeW6BpPgNxudUeziAgrPhihMbWlbnvx+47ImYQDgRtipYR/z6IkpM
4FXXntaDvlU3RJZmzH0W5KgKYj7H4GfXT4cBVqwOm/Mdjb95oFwTSeAxkgwL6AEY81S4jYOI5rsD
4EO7gADOFXxw/5blwO97csalNgqNoEEiiYSvX4PfgejcXgl/hkWeUfQVDYKxzX1zDjbAofx3AMMU
2uwE5y1R3Y4X5NcRa/cqaauGh/3yshy/vR1SkNerz1NQSWBuzkGfZPN7HCrsl0lM7RcA4GUT1p76
lkRLlR4CDkPV5fxbXMiCX5pvsenorfXaMQvEfbH1zSg/IJ186+OWvYon8NPIrGjiAQ+ffcy2I+ag
H0YAxr0eZXOM3npCEXnCs4ELp6WG1TUMAOKYXIEqN1vxzJSCPaF1oZGpEAMonMLw/e0D40gIwnfq
Ab3aVBGaA8oBnsgk6A33YOCJCRYS1LQPphoDe3cLGR/3KK5ChDe88+u1M56CCOdA2biuUDoHNLUG
zOSWx1PURRDO7eP7ZY1WCyH/0BAyrJ5XYi4lS/mtS2wyF6fHPjRQE1G/82uTz3Ek/dL6BuP1SzOS
ocaQKXfKMGUYLkwZuo8RclMWIVkKN1suYNWGg7DfYjBx8TcJampGtTQe/F97VY+ioGuRew462EWQ
9x7PP/EGxMe3DYLaObYZMNRj0+7LuizM2TYJYZNVZdxeXrEcP4KByDsnZK8wVXViRhG40mv130w+
QlApu2MlvzHqVQtULlj0W7az2HFPdXP7RX6/AadR/pkWdzb8ZDiYK3HGU9eFMWNyxOfgrUW+f8XX
+IpSWN1zqmS5l9wCT8BQo69YgLRQy0YwWoKr8126yVqwDVwqM1vZlQaoU4xAwubovadT+3WxhbaE
fTwAr/fBX0Ili26oOmoDn0ZVmQjS2t1XrlZdAxRO8/gkCrz1mQwUHTpankABTBb8//yUdMbGgMZN
FiC/4HvtCq/gVnKrEWtwIgvUitBrAKicVExcE5Ox20r9CzdXw265hXTM+GI//5woBTYr6AQjdc2w
bZUsiu4avtX/XkpH3zuKlYAvXgKuvnusc8rzklNIIM/FP8YCrq33kJfzUC4s9edsUSy7BY06O0FX
jQ0zN1lCj0N1Oh8iFuSzREJoC7Gb7kl3aUIThTWRgvyzGuwhjP8BkBQjWO3MpI8ggfas6uVj7S2c
t9FES5pB80BkHcZz4hcuuvS8BgbVd9E14LYWEUQeVGq7dTMyyD4A2W9dGjdfy9NtCUpbK643KM6B
TeCSF4fVQbFk0I27J7XJTzGibqWDr3uxLeitpQUJ/Y/3iVgcN0UXisYEWRyed7auUYGdrcDMSIfk
1Jchk3mEbb/xnlpkcEaUeErGklUVuDGVbCTpdm8zl6vqsDbJN71QK8hkBJms4zsM5GWdQUxLXT3o
xTpr3k2T+FhOTt6KKojXblJSnDXTxWNGaj4c9JeBYJwjhhSztrgaJlbKyHoUddJcy33fbc1JzGNO
lER8jY6n1bC5gv8Pv3ZECYIGFqPOSKpNsSILmqWTWdV4l0OHv7B/bD4iVq/cihQ5C0VTagViXkpT
i78P0m7H7a9ylvW0t28jdbMGcydnBSMZep9n2kbBV/oMOX2Eu3RFv4MIAUtdLoKIQILkSVSLYhPs
pczji3267MfBbIBjLKMW8xhPAbrJvvQ4xb3++skxxleoI4ZLuRjZwE+JT/skDGapZR6lT+t7ks36
pt+1l7qxOjmfcC+DpOPVL+cveTB3TjNokrTku6n1UjTx+lw8azgSXB7WUyTMbFbpC5yFOe7aBQlC
JYQhDjmfo7yJO4OtDbBTDp4QpcqqNZT1R8Wl0vJfc6CLsBtqLO5dWImGGCtPRTTHce4qDTHbHBj0
f4rv0cbobQkKqBNqPTfzAbIyH5NBws8ipf5JEedoBI6O732BzmY3Uvdvoeiq3Hzuk2mNSva7OCU9
3jRl6pabqMOgKsqxjo4w4yc35m+xzX0Okrjr2rB8s4tT68Fh836lfhK99XFJuFlghAn/R1uheys/
QA2qv0O1JDTafDkIiEUdyp1znAZERI0R1+DSZxhZ+IblDMnIppvH2cTXLchemfJtmSBPmgEliFog
9z0GJrBnB1UxTv/UwhfcXL8nURqhk+KR3vWPbvamoFg1mfrR8CCaZ+6I9E9xEambhte087Mxrbzs
Rfh3244gSNc713nxu+7cuxHPyxakerPLlu8NXb1DIBNZPgBt+yGVCXNnPBvwUWh0Ts7UO8Bn3kpI
YuwIjsyzkSrqzV9SzK6Kd5sYZRZUljrY8FTuMCXwzUFi3RVKK5Uywh0QMmpvgUuD9NpBsL8SpEQp
Ir0HDK+kawwJnYeL+y4QW7AQAPHdaLzpa7SsFtXn5qucP17ytQlaqm4P+rrQUXGtiekkU9altW0w
PfoCo86nhwnvv0gKcuVW2nwSzrckUuLLKw0ctzx9lFbCoqQFpQCgZwujJa+yD2mfn7X540h7ruBf
xJLNB5pcgXI7NRWcwGnw+IgsfiaYzcQrQGD3ptgUotZ+c/AoEBxob8H/szqZLYAYwZI+hg4a7Dwf
eICN/J5eTosRnaykRfsJv0Rof89EBPlEVkcRMQmOqvPiihiPszVZTa+oXVAyIRSyjMW0jQRfGlzF
CdF1l+ALXVlAwfhTHnC77rdfkHkVv21pRCuFOoRlTkN+zz/UU7iezAIg83/QvWsvAy+flO3ekv1r
FlykilRSk1XgkrdSwiTaaqAc3f0RTQitvHYxCz4BlkCLg12zTB7nXEutt94RNWJ2wyUvK4x4KdkX
hv5s+vD6Bi4KdG9p6qWMHzw30acPna4j178I+8SeuicuXan5tibFOjS1AYTosj7FaBWJQ3CS8oFS
w7kski2MZUrxtWIlifjMmVCOsVQKlIcAzsGluh9CGVGIHkpo3TaYPJ3BDBbBUNTMjWmMmsa31M3E
P873JZwPqBAC3I5Yd91FoXuZ+WoWyGZJJO+BtQiSRJtkdqAeFWFQRIZkUNFZ8qYk+90FqNt20J0V
FZjhG1smT23EJTOzZDlLu2mAE9+PZJMHUxljXdgzwbpdU0RiB+O097mDeacPk7G5tOAdmNbiPZ2o
CC1WE/38F32i+vY9LxVGfHUaGI8TZYdqkTkqET74j6kAL95ZRQOY38anZ6t5R6I7cPtjpncl+fXn
X4tMaQPKo0N41ba2Gjrd0xsEHbf3u9H70NIZ1NsOSACe9we7bmO7F2kRQlDagEsgpC7sBwVaL9dT
svr/4v379rkmW4p53bUVeWa9GZBF8TBWUcvzO8zE4kOJMg2gZ0jCXppEMM60CCqNmy5jLx/KxWs3
qPi0nfq3TTB3PdADOFBGZTLCBgyukTj0Q/R1LTML9Mok1W8bSerhZNoP93QRwo4P0DCgjgKX3oJ9
vcNvjx4gN5Z2IDkI2DUhpm1TX8/Xu+RCnWNReb2cziCDxnUlmHbSZBKnXW0wqUQYIiw90skhY+0M
EO0hfXb6tCkUwsj4x23nilO7fUJ1aeBQbdJmM3x9JqFn2e6n50vWPteLUQoV+kjsq3hbudnmLlL1
I3Elv9bjfe+bIQV7Om5q2Vo3Z420V5X8qKHS0tvf/GtAwCjkPQ3hGQW/DU3pULD8/cNTeqPNAd4C
JmQpBoupwqErp38Ys+5UO1wm7ZVjarhfA70J4drNN5D9dDdjwBS+vxaoU/4oOJxxSL6oolfBfnMH
Ch7mYodAungnj19vKBpBTyoQlVQtA2KVsl6ovCckxasO6mI5nf3J0ATCdP5eYICtiQJxeQsTMNuZ
Gvf6oUoQSsGvG2YmyxjTlgbP5Os7CPs9rLHiBJNQYS+N/WXtpO14M+Vl6D4DcE1qI2P9eaOtbdI8
144oNjyM7pK0XT8xY2atabZDiH+U2NgCfVJCshVC+fLYTyxFCoxG9RyRf6CCPQM9zHdzpOeQNgFJ
CvP0PCxnIbi0P7ppIVZJ+vbVKHB5uRixlsE9x5/HViILbIhv/XyG8xsKtlNtSobUT6gQZaZtypQn
fjp/4Zlq6CsFAE3HK2JhrqB5zsp3oXFiFzC/9puRKw3PtTXtmR01zPVgQbxPG5+NGEUDorRjx+f9
wuGhO5/dBH/Mzy2rQdxUDhlGXBM2o6U1izQhmGiyVqV2qaSrZGDmX+uDsWpgVaRyOjCAq1d8nkv7
B+6voEkHf1nZd0Zc7Ea3tH45B9Kh1dMfHST+5+397gfsYiAhSwY8XhoxqkuhdaIQnw98KYqXOKuf
0nvOwleBsZ69VftaL4wdsgfLfX0qIrAKk4cj7GH3dE5fCG4OBBwAT2LdJ4GHV6hbg/2F3+B4nWVv
dZIC5hGZpHyuNDilwkrGhu1ClycS4ZUUEoQ6KzaJUBMdScfqIgHpvYWxpDyJrtUgKYgG0MynqXgE
TaXolaa+35Ojz7E6zq8saq6bDZ2JNfS/r48Qp4pGPau42vQSFy0ImfdqyC5PyIGcLutJK/Yp4kFp
64c9Y+gBScOlamld04mIQqSEHbIIbCiAB9ilXIS+JxChx43loMm0n546y9NPtugX7FevHjmfKKdX
mmQrKszmxCs3iRDC3Ujxmm1tSI9KDsvbfb6pLanzE595ghfJ2oSn8dNQHsz5QLxuhySYHFy0CvFd
IC7kJr9GHVdogA9f3scTzcILUa8+zyB2J7wMdTsTYX0JDGrxdobJtyNA4dXfX5CTEBZQTU9llNzI
OGvkmSquvC94WOGL1k1bsaxoNOmFWgoGCN09QpH2aYPhw92lJLdydc2HGL66mvIOJuwn4RzcnDZ0
z5PTmJAzOTl6NTrhFKqoFnKyUK6C1yRihPvZWmTwbhQr79aX9754bpYDQ+QmKHjzc0jt5NY86yvj
0JuW8S7/hkPVjaRt6Cu2h4YoX2/dQAVQyp8lTtok47OCHFTzcQLGoXArc4QuI77/rogkT4mpS/Kh
2WcnZRf2OQOWfWcMEaTnsS2Hevhe9wCMrzTVYp7pBuVEW7mR94poHmJJsDXEcuvajYbOJrUbz+gN
+kWb7UwaBMGOpewePbOpkw9captcf4cC6AlQns/cnWyLj2cZb1AyWt9GxZXprSwRBt4QvBiA3hoJ
l8M2IsI7fC0m6/RGlxtp9xAkSiwOz9xGYHdDeoBaYkAuXR6DX4cJN/UBWnU+F49Rn/ao+gHua+q3
Gzxp1FpBSfm0K0ZlcxItIpOfq0m1Z1h20uRz3meDsgZV1dHC2Y+165FfkO1FXsISgHt/1ea8otLd
XAAcwCzNgKyAXpTh6+gIV0a666zzhWIiOdQDjcMFz9sLt1bOAxZggQjWgrtkMfCL5ttwh7tno1Dt
B7QOTcDvLO6pQ7x769uOvdOpVXTy7WCk8PMbol4M7s431jpr1Tv2S/MhcZJci3IbGhEEwF3iJibd
RVqjG73BH5H9XLve6CST/IRTdcQdHyX2kCETH76yKvM+tVWZikRqADQr8VKmktXapDACFQZ1u/Ny
bLpUr+Dj9d+O78UIiuSCb9YcpEjpbvpXE3O7YhLDqdRJeMolzUGBDGI61Vdi6kAbQuI2gLmbmo7Y
aOFpJvuo1icmNL37Sh1DIIsC3CjzRv8k+EjbQDAXX3cwSUARz+NWTxU8acBlnh6dCTSHICZq8jdO
hvffMswgKjEF+fW0fKLKrzSrhRD8DOEtf6N5FTMaqorMzFbZZg0/Dif+sKFsdNSolwzUv2vv1BZT
+kB7XkGzQYe+2629e8zOZ6yxKwhqx7M34aevoZOq0MDVrwDLQ4hEBpPfF618gCNg8N1Gzzf8fAo5
WX1PcbwzfzvtqABRe7ZbD0vXV2zJskGeLaogE/UYNXjpTFxmiW1ADaO3h4cpIMUfm+jn70/M5D1q
ZhC+AA09/4N82d9vH/WpLL0IWG0EVkRTAbL9zep8DDvikSbAgeR6qoeFg8P0VQxpXJHmo7NvHHyQ
tZbVa52/vQU027OeiawiYNYvjqFyTPU1Tpq9b0IIowGqxsxjSgnzj6pG6jsjZbjA1vQ7S0pxi8/Z
+IqPjXHwuPN2odaf74/ge/7ILivPXqF8pegkBhNyDTT6NnoAynpJkSp5vppNQc49aorGiwTZ1wf0
mYLuC+vhYioS4Cdg7EYImZYbgxN86KvwaO6TTqFKxYtGgUJmTaEJ+xh99KNGILCpjhdlktv0r4Bp
fhVuc4I8GcquihB1cHyaU4yDwcLhxwcM1d1hAY0oa4UAfJvyGyn9AWUZqThA4IyNSy7dvsmdiSc1
hMc3lKHxzXYphBlI//iY4JfNLirbfAks5oxXPmjkQlRxodY7WWBsaPvmXK+1/RBHX/cGdTodlCXp
ynH0Pg1ga1fz94GwV/GO9ek3Hi+RK4DVFKxUA34mVsrY21p2mGCs4LtmTCfXvCt8nxlh+48uzdxV
FJTxq0dBQ98nYMvGz7noTXQNDoMGKqAZk/i8GZyQzoWX+LkxF5tD8kT+RHfnorYuuMnRSIizERNg
I1xX50HTshzz9G7Q88AgwGCPa3wBZz0XRKC7DiEw0/HAFVZArYOmp+UtC/9ip0sywmIQIyn33FFl
3ScxSGoy+fxdbCVgrKVK0azdUIqEB5hEusf0MAW0jbgosbAMQi69kW3Gj8YYuIqPC6YLf41vOjsK
4IQguUHh87+Rd7mc7agw+4XNE8wpQqzcRcu9yFnyPDHFC1QzQaK5dar8dkJ5NOmYFq3TVCIMnT1J
KlTI3UHhWIOqXQRhdaPkuL0W/WoXMFnsW3BfBJLNHPvXUXQ3vPN7MUsPRkPZn/G5z21iz9Sff/gp
1eGqbL8iccC7nRrTihjcnlAJZYAgwRL5mlEIRi6jurbcxF/goZ8SLqSw2IOVNNsD4tY5QLIobl6C
rtTfxW4sBVCn+gN/xNr4j35HaYHqCedUePtircTCGUH3sbolDXJ14VJ0DWmr094mbJfGLORQDQSN
YfFI8/9ANXQA1t2Gt7K30kvbdUul+TDRH6sioa90mkTVmaecBV4ztu5aLUt+5BkRA76hnDPCxZhz
E2UQMZbte9vTN0US/oHNztddxTetIQYdilFTqYKYc28WaxLnSfjHB5oOJpW6ntZtxV2hbQWgzQ3/
QhJBwMGZWperoibCy60xbPxfgP0jJ78b8nfmiiaS+sPPdWehKRg9HSXr0ygkZY94HlelcChCGhZw
2Ya2ATw5dC+QDj/1q26+kMztTqM7KBsOni2CF1l8eXpbX8Lvl4wZBMYy/NRChLUAXvLNGntMhQHw
aCHbab6JN3qvJMhVMNpliHNnaDyq/ArSMqlF4ku53uInKi9ud2DWjM64rjs+DRPemZbknL77s3Zq
+W672kvIdxclAl38oKng4Wko//gFbYBm6TazsuAfCmOEDnXcrCStqt8bvu4XQXDGpdw7tvCkEURd
TV+/GDxdRwvZqNS+D5IKPDA+2McuO1qoLwMs7W7DhE+pqt1Hw9+GFhwW5dW1ISmK1OsIqIE/QOwR
IXn6MvvAGv56q8xeJ5InmsDDFQPwxVcKz0AueuQwdGOMPovdX1BZZ4aGpvw1QGLJlzM2iwWwB0TG
u0huXnmBFCh3Q2qUF63ZxjhLqsvI1MdNB0hShEeroDjS3gU/y/HAi17AQA4Fx+ZdKD6mtyKdI05p
gMryd+9mQHS2ZLMyADUvy/KXBz+o4DQkqm9diIE20ihOT+X64Z0K1knzL8cSjcsqnvd21Rd3yGcr
+iAxmS0jEZiu6KYh4j/kA7/Ca+RILLJ8EVUacj5frXBu02DgP3DLtwRmL6+C3daDsBeyi3whYAXN
FAkrSAQinka4kvGFMa3baKyRtyj6x/HEGO8RoWEKHQLBjQMVgLHfQ57CvCAjwPVyolhS6OuO0oNQ
vWh5F03+b1JEhj1fZsAsuiJLgDDCW4dLqMxcUDYP25p9Ifbbq7Gyffw6e4Py2pnB2AsFlrXGaq2m
gAR0y87nFglTIZVXoTJ9Z7DYJQKtKLO9kyK6Gnin1ihFyfHZU122vRh/in2hI2olbJo67h4jr+Ql
zdJvcvmbKuW2K3iKB5wSeW4NhC15FlLj+NIMWqNaYlC3JzWMorUP6HhieOHeuzl1/+FkwK0uBoFy
doPQakqjrojfb3HIk8VO3YHtPabaMUGETlcn2flZp6mUuUjLNCtTxNvFrypVMNgdEtw1fBBQtF2c
BUcsDPKnCLCEOQbJQ+7nYT69liPfrtodYqfpMOqZ84L1Z5m0/kVU1wBZrpThFhuMiqTV2uSPZqy9
3ht9Zex3uzx9sidiYFyOkpEWTfNTkIlpHMdVAeonX1rEV7OIw0EnY+vrDePXOJQJ5uClohnmcIc/
LmIC9PLcyt3zSoavwmZsRHTwbDLmb7jR+qjM0hOiawG4Yn3YMPCAZ/M6DC9k6BUBT5+iwzZiNyNr
1Sf1i+pCuudgZI7AfJ4ZDzTFPl9R8Ae/F9otOt6NfuJjSXKGfC2LvOW1u1E2TcdDt731eaWsN1oL
L3KgC+FHn+67iZQmIqFvGJgmA+5cr/Q/cMPEbcqpnjsMB4C+uxGxdGT4uyvRdfXtC+7onGbktCvk
XJuJq1OmJP5z6XyszF7b15VyDDpt46sL0fr5ZAzKUMZBKuUYoElKcldN+K/4YutZJi950g16fiI+
eriJunyXld2lDjl4H/ZaFbrBJix/WK2LjargFEI3T1Wff05peB7sTS0RNIi3r4152uo68JzL5HZY
4CP0Tt0hwgCJH4W8DL6W/XhdjW6Zm5lIuxTnN78nP5jKuN/LcEAWpiLpRyN9sSAbO4H/bkrdNIfS
GNmm2ZXkkYpHBOY96lsmgfqSS0I2hhiBtcKyLQoSyaba6QqPVX8sPRmNhx+xPc36ZYgNSjVl70hV
AsTHciy/7FPvlUDcKCK9c/m1u/tw4sHbrSaJ1pt2U7/wUDoaa6OjLuDzyDKoJzH6lRVbhr6qYvwC
KEil+5bJzK5f1iEU5PHLegelLIrlNPQknelp3YdFClbnDOb5gDWp9oXR4F8K3nsA1DY51w2TUHPy
SsM7gxAXNpVaFrVfvJXoA26xACCObuJoAEAVCBXJxDv9TZWbYrlNSro5v7TK0zf0GoZZxlEfc2iY
xWoMEpAEfG77AcBdWxbKPiXnwse7dX6WoRdRdt/xQhyIsj2qmEmZre4QCfeYfNy6L6WnTCGAw3Xe
DelMVqmsfOoscam0zIUEaIe5qgT/CFSF3SlppubvMCUBJvK80ZtD+nySMx0GNz+TG7FK1WxMCYT6
3e3WOfdqp2lFGbUswK7vR2W8Yg3vP/72FB600HHBtYK2T1ZRyupeqU6dYFSLFZ9fKUvTCKO7zIG/
+0Q/aZJUJyTfyGlsmQ2UDCeRK/7c7OeKPMg8RT/2E/gZmjA61JDfuynfzPpJuaGrMu2ec72pgzsA
MVzOHRTvnryVc/gyGD1OIRBNmYjXNdW6MTyEPdF5947BW1B4pKzkmOqPA9Syx5EeT2fOeRLosFT3
d14OH3d5/CWQ4eTM1J22jw3XLpyUmOw0xpDxOSdTjVhwSvLFlvXrruTiJrihis7O/UjnLIF8RRHy
P+3o1HlVxbv9h5YcuxsRXyYItnsmb72UisMzQNcAsK+xP+EWD4ksxRCPiHiGvmOHVce9owFy/x4B
NvZiA315of5+kknuPiReXKBJSN00LU3fgCxfTvfZzCSEWxlAKuPjMIE+eYK4zyl7fR18geWqPXEM
FwhNa6g8o+e7TJydi3/lv5sYz/8OgTfJQraJLAnMGyRzM4Y51ivoNpYlSEhMP53X8RN4yMdKGi3R
/tV5cyxSDSKJn0ym22XkxLJv4wO/oaCIrQjZxKRrzJ1fFp/cCbq+ALf9w6efd3ySBcc4GoZqW0Ao
+bn/Zj8cqIcAHkaSFlqczTz5tfpUXLMDbcEczmLFXI5H1iPmjWAxSjFT9w3kCl6u162j51UfMeeE
corw0SyKH3qp/ahHaegSvHslxGpvbxRQbTUBSuJbfgtMMELeHQpLQ8aMl6QONDybRKY1nCvY5268
Q/KGxBztZVe7qe/yEB9dUow0KH2JXTO8VWWX+ci7s7z77gsXVX1iqUTZ870gO/LYArB0hpjJWJZH
Mu+9Du7rbDZvm3jHCtMXNicl4U+38cQPtRkmt4GqWlxcUp1tObJi+N0kovagq80Ug+t1POKW+3sA
uRCNBEp/ntxPQ6p3jkna0EXgrgkz5q9F6EoNkHP6zplajeHZ2hY7CZH7D95Ebz963HMI8dB8JHrl
jXsMZq5Zf92eWG/Dfa9pEFAtMn1Wt8HJTB8PFCRs2Zlq0/o5yfPo/dWynwhaBAS+ZLsVJZUc58wj
V8srEjR6RfLbpC/IZ6hSo2eYLiPkW1g27CmW6w0EWJeUHk9ZOWN/4vvqdhydOmreu1FLDDy77OjQ
Wb3hejonosnIrXlcg4Ob5OplK739IkrFwWxlABbtQMZQKjqjfDos/gDe/8MBpBxSn/TaEmuhEqhf
E8CvH201uLF4e3hW2/JctDtXNKK/LjvT06YcCbQMEIR6++CimId8KoRlhUN3qjAq34pA8QLcVn7g
gtx8ydounUafauCbI9FdrCGiZwTvmRxWRTNfL4O0tQJKN+kZ8rP+R2tYwURR5sqyb8vGUYxQqdIg
zG7XwVlk6WeSkI9QdzPIf8QbXuarIbf+pO+lYfAFtJIjoyCqV9pykDvOEZYVDPqDQnNJeBGjEZ3f
sBm2Qhf+DFa6OVlneRcfpVJKvRlu1FjuxzNxfFamAB7dBu4pKcORJqTN+cWmjX7cNM7Vfa1y+kME
28iZXDSzbUvkPPJRwU7JpkFNYnxINDuNzy5UyJAAxYz5XxSJ35/3cYOFPV/oE3pOISayakNRU17A
f0Y9+yY45cXFE0QUgcw1ihXPlbY67vUlMFiVvGHL8MGK8j8TRTGPUhmph8k033HDjrM6PjNqNlkA
c1ghZQBJEJhX2S8G7a1tyj+qnDUMBIqlhSvaginV6dVSqmFYk8bwdLwwRKCr3GTxPvOSkkf9HNAZ
6mOtNxSiFxLt19RHVP/cMRKp7Mago5lu8SNR+7di0pcWa9AMbvwtdeeGGIQBDgEGTutx7+toOW1j
wHfv4ec4I73PRPAWYF+TmtMbBKAVJUPRVe3H0+zUdeVngJfx00e0bX39rOtoOPtAYayCH7hYzbK+
ApyPg0AJQANKA5mJ1msYMJsefxjI+HmFS3Mm7/c/Kwo5Lh3GeX5KizkxRSdvFXZ5RPk+t6cDtouQ
+q7hCvLmccJskDEseaFdRDo9yxfPZJuXFu1p/rqPVuT6TfHN9gYaIPUDC8LI/jRWz9ieN+Fxnehe
wn8dcMQ6zJpPEePbF7edPDvWUvE0uzzIxdpOv0yi9FOlXrfpWL6WWky2TUzP4VPB+nJmHUfdtbFj
9u8Un13Qg/148LQ7zjwGPnPsApT5CpU+6zguo4oO2ag24mIidH3/FkvBxRPvLZzVmZ6NzM0LXQ5Z
SMvh1fak0cui2e3cm4+sPf3YmotmRTxSCV9Qp4Z4rcc2WY+V2BDTRdHWZeIY/ck59jaginvCdvYv
B0sjd+i3AOIGF0PD18Ckri1Zq2gO/TWrDi04dkqmD0vTEJi9gwMSgAPKip2faZsrNe2pkVXFMJ5A
inlXuVyuj34UpfUtsw+9DZDHxBt0GQWlCTwETACgUs2n1ELuK9B9zmn7Jimi1bh41bHuwIc+2QxL
16+wYlXq/C06cMo6Ta+xzqpKNZLqF+pjOY+VGIgpl7i0ezCut9O79IioNEj9TsPWApCjrMwCUgGq
798fan9QjjRdqHU6HjFUtbraxzlSoiIOCGLSq17OTtSZP8v6X2TkXmvHycb2OVv5tlnUDpUE7U4O
CfU1lfNOlT5LSFc1lbcBBYm7lOW2514t2WOlXL/okb1zc9lZnz0JmiNCo92LeVmVe6LVdDN+ar2x
0+PyVPDCAsTqMPH/pzH435+E6i5LtAxNHhuKSHq+FXFQahQMACOKvgrKDx+KRMP8qQHbw+UJt4co
SDY1dqGbPJCzGEFRigow3iT8uPthzBqB/iguZ326YYfHwGfO9/Ae5n1l/lMufnJRkZNGq6DAGM9z
8JYE+jf3x+JJoMZAlBGFwq0uhmdjIsuD5JwNOzeeSWAJ0TCACC0z3eK9fKjQHxTd9QxGWCV1dGpI
iD+6keCuE5zv6Xo0Z0ppZhP+kHUH3cLQ7NfWVwhbpws9vCSv6e7Xfe4nIRMp4NVgCsfRkD0py8ZU
PlZGFA30buG2yXa+Z1MyGyhmfAZWK49tdNPn1m+isTScFqjNuvLEowhdkhozfyIkvFSeHIaw5kVE
GWhg41NV8LwVvR5ehkLxuvsQqGOdrNg2sUIeHEf33xqYspCBApq/k/cRU//bD/6ZkDMgqucaIKgO
czyWTOxp7OSPVPlNTRSxPsrG2WoXdDkCLODccFl/rI3ncv92omZRLERUqDg9JKZiVZFia2l1aXBC
z0TOq1Uxfr8bAs9Jk0hZQitL25t0oTGbwzqS2UCGMq1ViBDjG9FXTSWoDprZXNlBHDYCQNA+gQOD
GpQCkSvjOcLMt4wFQfmhj1KypBx3GxLlPpzMgYjA06DxPd0Q+vqy+99+IGyR56TDuBA3KarUpee1
1Dgug+LtX7szQtllfPaj+efWcOjYBBj5HbUrqHl+y/o7r5JX09busoIhi4pgI1OyNoCWJuxmvft9
HCh/fo0g5gHuiBuE2GE9exO0vOJWqgh9v4ETvu39qouAKFXDhq9sRR1s2239jv3U8hYQ1h3uvdHq
hbbHS7StrXlw/EihPjDEU4rUpBmXlyRl+dBQffEZS24FK+isq/33dsOs7mF+iMBEJo2aUefTVubT
CD/XLLAM1cyKtPZQC/qUOkCJAklP+gSXI+ajLKHOLxoXm1KyC0f0acQpdGDPRXeAZMGqUFqcyxH1
ru2ml1bf2qfauyGZSaHI8tsUYKvhQ0kC4xtW8jAQGTyLmLZH7kDgyPXx8OIiVCWBFCWZucfZnqzS
DWChRuzdpA3H1e1jAsmgOxwHy4aPiiWXN1ji7QzueWZMuyWrw/IwvJR5i0A6D0veHb1KGRMYooN3
AriVeWoRRAFAMZKUHyL0+QxYDmmrLJWZPeopxS1OERjXI5AmhdZRptNjhmvBijGCkMTH9OmN8wmR
OFAu2Ozyoxn3mSMa2XYPtMdHTGg4yr/EVx7u8q54LecZkmEtJJEbDNg4qw1GvfKa08Njhk2Y2E9h
ZFw4FLAe7Hy81TaoRIQ8h2S4FuwJWYN03vJokG63PrKMSjFi3AGK1cwoGarExP5bFAIs3KZgl+O/
vhVE+xswJ5EQB/962/RiAGMVhnuahufSlmCl18KF682z8Smq3Kwzmmo4ncVH84L39JLb/FcEL6e7
9iYwcmExQ1NchJhSbsGmWvs7JuvSLH4sdR5STSbEoZeWbMZTlX0887oEogZPLvxbJtLqDCFDSOGm
gKpFVtO2TStwXWPm6DAYcyuq4vhu41f8eZw1omEzjol5XjWm0mhB+5pCfI49qBqB22PyFVemz/+b
BoyFa5bUpQW1BoQ4qkU2CqD/7OJr/tWk7r3gANcDB+l2lbTQFGhbeuyKPRzKAMlhjSCtfO0S0bfa
1HcSqxkBNYLbB60h2V/hUCnX23dN++MXgzrf/wGFNBkYxynBuYzTI/VzYn3yRIlk1CY93u3D82c0
tKhRG/bxeNm+DBoa/FbsLo1oSLgDJYWOSm6KMBBY7swJqmfrYwPuaz/Vr/G5O/3oDfvn1FM6KQOX
cwls1KZVolW7kLmeZZQdmnKavD///x6ZHx8j++qgc4VEfhOIn5EBBc9b53IkdNtj42OrVJq0vJbs
Q6oBaKFaHIe+mxHCvJdZr9jBkZOnXFcYbP2ZKCnlznfi1gsSoBbYoOr8JtGafTAfyEAK10J2/gM8
SF+VXQwEHQ6U9Vpe4jO7asEzDZFyiDsEtPxzyWUE25fUkscJcpB18BpMoQ+Gj6RjUlHqNMpa6/Oe
ZyC8kU1irMxR6hR3srOY+ZNfSQ0YaDNreZLRHi6FNJkPlicaXG0sCco5lSv2o8D+hPZaMyb8R7wp
Sj9Ti3qjvQRxuuGj8xuI2hoBbsNiKVtW5Coemoc6XAR2Qz7HQkxl6GIsbYlUETe2hQ2QxQz5OXwH
jL7SleR3lsPVYB/Am2cZXk2CyGv9wLsnVgK/dp0SRrebaGoSikAuFc4HV9x298BHbxouuvDvhEDf
CT8koghPTZj+JzodPzumJuhtgutY4H4WU+hJoo6fhTRSDFLTDhBRmZaIz8WH2z0Fok8unXVSzOnZ
xvQAAJy0bVP/9roYbQrGqXJU0bOYzLllfuCGOfM5GFrNhQUVI3JOkfxXj19Nlh/KyzXCLIBWXr1E
a+6hBBZSakb7TGo8oCdeS5WhwO5JzOsVHoBfIn52ypfmHyu5hiLlR4v5rln66dwdPiLNzjOSQSz6
P5rJ3/J+bjZZzsTSEvCvNjbHZNASvZR0R7gUVIa4Xr6BRsPQEFV+FPKaHg5YvKvO0RaCNCWCJp9H
39qbb+VoICmzvescICMfqstAllGXW15q7CZfP5xxEsaB4pZuZBzXvxkg1DHXZuhaWcUwjfBslvue
pq25mkz3rk2W2xY2MIvyDuHkDhqKBhWK0jI0zlia9txBIyIpEc/HM2Nl2iCr1+jVlYXAc0MVup8z
BbCKkCE6SvVASr/1HbqcoLIBhENYXmdTvnHL2s5yY7UtLvSEOsl4Y4UbNgquvL9PeANZUsSxIDR3
5nAEBAK8RbsGIWWWvLMqY4PYG1E1+i+W3qAla7Fmud3gPLArZ744d5+HHxk6xgL+3PkMvK3cb9Id
8iEWh7gtcYkYTB6BBg+unuzuVRP0XmUtenL8WrT9UOTD7m3lz0ySg0wWWtXSMpD4+PNTnM4XsAns
qXVyTkcQZ6jbQAO613QRgy+yhG1XFBdIHUycVfCjhE94i0FzCWRZwCbX3HsuK2io+9TR8AsA2XaZ
kfFqAvqyOJ0UFik35Aw+PJgUPx/5Z4IfiN0l/QrMhblogKkduMRJu6+58UyTV9uxFE7gyXus42e4
JibfgcAlQy4aWy9vBF+HeVsh1Uunz96Fwu7O8+CUSoiUTI50tXJ3rKPLEpQuK3AR4ZM0V3Rrv0sD
eHt5GT2sHY1dxWIYfi3XsP9NkdU+eYIoR8lExUwT1oFap0FTSP6pUVdGabeCoBQVDbds+pOSsZYI
LmvF6J4G8f/QNJ/ppnnWH87yN3TCvPjiF8lWmSegdA0JiYI7WOCV5OjRaGgSPoocO9f43amlm04f
TmRZ35Y/ewd8jtvb86vunCv0QMDwLL/3i9mvn+v3/Lb8X5Ku23+07wnLMqIAPk/yfOFpgCVjx4HP
w0l+HFQNErHIg1nZ1slTLs1huPvnpzu6EC+Avonynnyu3soQ86pGQsTttrySgQ/kgp7IGnSFAvOG
g4YqK2mewSu5EgjDrd03dxA4AWKQbbdsGKXL/PX7wqU8F+Rhbw6iHg8F8B9O072fB84RE9C4h9ax
/fmUZpw3vHoUSfB6aqPR5zhdnrd4o4SVsJqnfB3NCT1JXI9ytHwg17EwPuo4FAYgaeo5mtsqr+Jh
JJgcXdznztVgweWYU0xexnPi8I74p6B9qEv2FMOuqPLHEaITBSMYwZNYBomhqbEQXpPYSI0rhiPU
NxbSXvO8xWTJIZVF6laGnh0p/5TVoO+XAXk7Ju1VZlrZQYNyb8j/gOqrepj1+qCqdc3g8f3kYMvT
NSMKv45Sh4Il78lQcB1/PsvHI0Kn7aDHPgBYEFRIwWnKI9uKANCy/cg0ZderYM/53dtAGpmMNJB+
f8TVdtrcmy5KUaB9urk7FraW5kiBpAVJbeD2V1A6+5yKPJkJ4QPchWsxD/+s+N0kenfAkBAitXQV
njARcLd01cxdpzBzplH5XMvYHPLiCUwprjrD7NB+A2C/pbR2hDnRmR3MY9V3YPZQsVBDDpgvpKT+
lTXJHP65W2T+sRW3M8a+xFNS47AQy7wOdyxw1r0ZIp8RaGXnzfDoxvpHe5UQzZXMt49BG4Atp5Dd
WLZH0j/Dh0ozp0epHegCL+iRBGCJawh9CkWtrnrTczul+VGbvJT4DJH4xE1AnMB2FzYiKZp4VmOy
lDVHD3pP5+uaFVKAMEvD8tf0Jcmlz+Szj7RC1uasvFzcJ+etIMzFSUXPPZqg+8s3448gDutC42Xt
Ik3i7u2XbTFUKhtS03ZVIkZJxt+hWdciXZp3dr8KCv9wgz94cAkDBUSAUjDZKh+i9NKsvk/0oXhv
iIsG7HtaWp7LT/Ox8bPpg5AsYQMTAUSreGD5KKJ2Vdjnew0aK4UpjYjKYakp1fgiaTsxHH8xVnun
F9ahZvjxAMuwlYFAqGvOqHs3+2cVl+sR9VHbSVn4/cROfS+aW2LpsGQViYJfzHoFp2K02HNSEIP0
b2W5T8cGFUTcBvZS6M0gr9spj8eLPQS7zZt0FI+DWUZdZeF7+LlZJ8WQI96oglvzjghuku+QFhNn
5gE3nbWn1xvDTJBf8n2sJGgrPgSBNBjPY3xr7GdCviiaIaDYpYW4fBT/H8c29n2S8Q9xcSp9MfMM
8z76pD30nBXlndyahezwvsHeCaGSXAd1ujNiaK8XAvu1AvHMvuXcr2bzdKhMjc6zpzQa8HfCQDoy
SJv/j848nA8zmxGGzMPt4Qsf97od73a8ugO42V5YvX5aUdi+eIkVW3/ReYWOgQcGfWPUGNqm9QwE
ZMhT6Ig0GZdUCO2tabI6+gqeUoQ1mXaOUHmmwXZtA4z8m5Y1nwk/L3dIrVI+m3Msc+zzC/D+xl2q
SA6tej3TtW9dmuB8HjxPdvuN4wep1zWEteD8KLz5rGjKXUFZdHfTkt5XgXbz7X9bFvrpkR+7duy7
g5TpdZ4moa/OGcAQcLJnGhP/qYCrLeIwOiMxl5IbIuELVexzqnzZjRsNWtHq/xc07izV+YeAVJ8y
Gickw9YlPJkKSrlMxC4QMJTrRcA6C+YrJ/PV7ItE9/jBKuXEwYxX+vKWIKwiQQDznlcUP3GlZT1U
zRgo+oHW5+9863w13eUvOqjv0+ltOE+f8836KsFa/67c9QiVirHiQZD0fDvZyvekiRQJ8MbFCNCE
gJ3XHLQFClNc2BxJJ3iS8Z9Hr1KT0Xou37Aewq164QMy+0fC4d0yz5wWP2vJPndj3pG0bVpHFIuS
xwOqEmtlZM3wAdGCZzKVhwsSUPVgvc9vk6J/2FEGopDtMkLPnqgAO/YQeV7OvnZ2UHv7/KWrt0Oz
l1+egLlGQuJsRUxktwfYcby5RIb/SRR+ZuMyBYDgQHmjGnAwH/WlzEqNUgv6iHmDEATq7we/U4pm
aqdtsnsmPYUiEbwWin8QYrKzfc2kcJdXq7/2FYixa+c2iIWq47gDqwdCU61P5b3YNa0bAzDZ5Yq6
oEqxCCNRWixHiKQ/d6vUeocgHVTAXAK6WkwfiTKzstBjpx6iTWN53eraIomp3ZLJs4HJisB30kKv
xG3tiqAkpPJ22sYN3XuWqxXlM3go8Z91kl1nZbUUjONid1Gh5ca9RxIrmTwJ/CYyAXdaOTTxk86E
apFw+NwKn25DiTYAwPJoO32amY51eb/bxY7AItjl0BpNf38H1Nmf8XeqLwpB5SdTJ+qngsPkvGWy
ah56bMSrf0nC68YiIDgwgcG7S+60ri/BF1Ht6N/z3oCnK6OX/WH0GeWrOwT5iDFRSQYlwYS0e0k5
9KQrA8FZOxsis24TMZzksdqjajxQYBAVRvfA7xYQcEQYb8YdkT6TCI0YnNK6cuPAPDAaBin7OWea
7+hi+Z0zeRuK7sKr/VLTQsyN1N7Uq45O0wMIZvTB+KtJlQveZYRQVE0Ri+S87mcTp3eVBRSdWzTD
G20SdtvzaZ65hglxy9/oYUNX+ibv8OrMg116z4XhOGRqsNrqqcbLFFGFUvn1GWIjRohqeq6SUtkU
wbDD26AKzfy1bD/fo6aolVw/yS9HtPoC506E27R33MXsEpi4r2FVAHNoSdgNjENyKUOU6UcJUSc4
e8UlddA3reiDaJBeQGNQFSV7vYWpdVhndEjK80Pf6H1W+i7ltprx9aAB5VRsBmt41qVa8B3StY1y
/Y8k0R9jGGoRXl5++WpZTl612RQsDn5DNdzmz6zpIfal5vumDhzpVtVSV3iYzbyz6awaNVZlP8d8
y0k7uC1OyWL+8OoKCDknv3xHZqsA/eMi2nfRePot4cqRYsvXhCuOWvjl+EUeb1hFjSmkYF3GSp2F
jLfVRRnfk+I8azdYL0xDJ1Y1YEMEwjFcyIsveqZlEsB41StodBa08pnidjI7cuQ3qSysulOP+tVK
lRUIRGVzxNnkI9YeaaZdIqqsdu4qmQwc1yU87zkIpIfAe+4DDe+Qmu7RzTfZSMDTp4AFQr94SFtK
vdNdq3gwrh6BzKq0sqL+ir5nzDozbi4SqsGUCOoR4GS4Z6HFl5lX9kzGqGtgOsM5Hw4nszdEnUA4
RXsXJEov7tCDYVzPV4OvtjjizaP8ZO2170Q6MKAlBbdlpDibew9pS+ZTAivtkgij/xCMntK8Pg3v
EfKofYrpXHjDwnDxgXN6GNGEWpq6x3r3EDuwzLCrxkdVE50UIQl7oYYaD7ybSJxolGX8X0Elfn1Q
FjMAPzdLW1cKHr9N8ZgD25Lo3s4XECq2XFfspY6+Apy3e77/1JLfvPc6amVy1hXx8KyM1OlwM74M
CWrMJ8WduAsJRFWeAPg02GLEHoMRlx0OTleGmZySSOnfuw183Kt+GTlJTQOOzO+NOXeAWXK8zfYi
d0A5MWfy+QU9H2Q5lI+krOrjT6cR8LSMD6yByrtIYfC9/Qt8BfmPznBrNr/M6oiQicKuuOGRQJFg
57RGJ+hU48H85DjNgwmRTWWSZu/sCO7/Mu8AGVpVlhiibZDpgsj1+TReRM7dCuMG812YSSxpKGYo
QCirAq6AEXaTWH8SUzZdTRGR3tYJ4cQwynJRxdQz6j7e0yYVf125OihAqJQbfCDneBou5sBamI2e
JnxtGJq7PnV+vMNj02soQatANykHx+M/Km3xOmWjsU1YLAOwZiWySFR4qkXi5Zn7oGWQKea9Y0n6
0LXJPnjUjx0z5GcH4+OGeYT8TCPxS9C6KoWy7Bxhihu1A0WUzasm498YF/pOhN7rmaD+soNdrwyX
LSE90JwGcyt0OQSAnYlDArBdrzQhb9ioXkc9DVPNjcmBfh07LtlnQhqZiezX8gJBydXiJ2Ct+Snf
Q9vVrfRfIoW6P4GoF7U5j0YFWx7xWdyUae0L4b2OcKNnrJjdN0UhLa3XXK+zSZCmSMfd5XpoSPE5
nkiBEtCgJF3vRNlwAMGai/u45jcpQVwtbXD+U9JdTBd2T+4rslPt/2plxwyyD70nhLv0gRUYTekX
xHUmlbE1ZkOC6GabF+K/g0CyFQCvp9mXTY6SNFtTz5VPZLCEqK7YCEarBBM8pSuGkbXyj1oreCXI
hsm8+n2pnH60mDfTtyGoLUSLHHnxVQ59sR/9kQkD9maA6YGwasrHHMCdF93a8APKtJc20mTf0rbZ
eSEzse5myY4GUqbQ79l79zg7XER5YCPE2vGupXVhKUqe3zIJxQ23KtuU+2DXFRmfLvqkKDmBqlGh
ri5VT+j4AXB5PYIAnFjhXhDAAbCJ2FmSao0ZPgxnfArgsl7kbZXSLqYrTNT+dZxHnqr5z2ORaDr4
aQFsSJi3b5Y/Vr7/o+I5YGqxX//a0EW5rq24Z1PRFcP7+M3MNbumlviAWhYoS+b8qnSwbHnnvMUY
XYwB17JsJuxkatDDPY+HZBnyCyOPUBepLGAlh9El4yPpjxaCgXHo56tC2iOmbGVeVO3FSgXlEPU7
NWDyb/BHoXkzBr4uTvt1qF5G1iblMpw9/d3tLS8G//jcv+ucQsk6QcqPNVHSD6HoAeX+ivQe3d5O
+Jbvscti3i41abRkEfYaviPHdFOonboLu08MQ44vbM5dKqfZWKT5hd/nRWfK2msF3DUHd8xvo1VT
guG0hl8CYZi6F9iqY4xUYY71wIzsLFoXQrasRWB/NsPK8DghPZVco5q6LQSo4Lcm/ujZV33OmM+6
lOuxno5Q7crLT45U2s4mT/RrZmo6H5JEauWuG/HAlEkmTTYes4KWPMS1V3mahlPl9KheF1lWnTn1
xn9SZr+x0isxlLyShoXUE9S11btI0OaqdSoYn9U1XFsEZbY195UY3iYigL1BmHwHEnOLIE90mQJd
jy9xpf8kqmpnOojlrbS8We6UXt7xp1Kce3N8rVmQApRnsApAh+WKNokzLyJEG15p1GI4tSo3zAlO
I45IcwJk06SoRrpJ8POVwPr/BxNqr1bGjTNwSyz2Zq8qezdGydWmpjcjeXCRm2oLdelgN4cRxqqF
Ihw9tex8JzuqJmphsPNTMEEnkuu4huwP46Se/kPcJSX5gwp1RWrX8yDhjIcgaaUeIzJgabGQcrI0
4fr0VJyY5Nm2FLGgdwBkQPikxZW/+UQZKXfJGV/XAkXYiB5CXoRouTYXUMN7U84V0yp7gLFvV2HO
2ZPfIY6JZ4vl3/uyXhZGCyejGZklgOfrLv0VInyPDs7Z0FI9bPwI+CxwPsB33fYPaGX/WPtmvN3u
4QQeZOfmR6JNGrG0gxoabvd9ULui5jovCgwnclST7BXN/tFXMVspLPdv/Aqf3bLwAwPLbwRbaZT4
v5wmk6RQnNZ87TZhUTc1m0zlHdgk3Yvkl6xnD/GqkinkMEs7y9/K8DFDLpgm462txOEQz7lxU8NM
N42TSiLFiJ1p0XR3sa0y8Fk0zrOtuso/gqia73l5fmaJgeog+3sRLcRUoDSGsGQXc/io8c+30/GO
ulU9cCTI6EB/ITxMH17yG/d0LaeeQ6UayKU8NNFIsQgO0MiWCAGHVzO/IWqBFRCWjx1H99o1nmxp
XOnIBFQKOw/TXgcONV0EFbfYIZcriKAp8Iz8qyODdetnvxyElMQzaT6oRrdBzNE4vOhNee+d/qqP
Bk4PUsU6vrWRvod64at4H6yls1FUv3tXBUW8ht7gU2HGSjbSgOLYA3Ltk1ShqQkm8aNHHdmeqwLi
rYymPAKoSe8avFZJKUOaZDECEnpOp1szGytmsQibBgEgZp6a4fPpu2J9iRewZ77Z5hqPX8EINB/L
rIEerkdExd+Jp/b2jQAf0Bsmz5Sj7LhnlMpYRWK9LS59jb91z+GMZ+TMDGYrKDqKs6dzY9JoRPY5
crVCPrCGWDHLJYQpIGEj19vG0W4MOz21x3WGr5pCuA8k+axEgu+XmJKLb6cBOH81Qlv3VGYh1P1U
Q20vGpeHsu3PH+F+ZbDTSDwTSzX/rGdJa0hCS6aAPAVvs2iGVAhPpoDW/EHjI0m/JScJPgagIcx4
NaxF/ibV1ZLVKLpHAg/QlXUnz32szFpfBUjfieaLLp4ZMh8ucpDF5zJ+hX4gZfuvf8DqeJ+2rcyZ
h3+OmU1/Pm0ZumOtZBssdPGMrjNn1bheIzxH1huh4JykRHk/qMEj7P2nOFOXsMRYhCzXSrX1mZTS
PDHg2yCv4EIeL+3x/ah/uiBvNo2eAlReC5rTlAD5xIbh9ciXE7JTOKv5xz2uufRhnYa6eZMByHcT
n4EQV9Yb0ZSVjNFT0CQGDJBwMKLP06f4PSBldpMh/GWtnajMXCuhw2DsyesV1poqd+y1QEUYFXsp
4p6QU6CCbRxLS7of0RvrrYFQcjz54hUbBVJEgnoYNnvD6KsBlTxKY3uFxLSLC6KSKp3Dtg7RyyDV
62BFRzr3iPeD2lILeNej3s5TonLHKRqYDmQmU7mNDECku6EX/yf0H5xoTfCASpRu6/2tN3nawyAj
f3JYZW5xffXIEtychsQtRvSIn5QYuKrJ8Our8XeR7rZeIKxkqi4r5X+n3PSJCDvdq9RwPEVBBZdL
rYzJYSn9smV0um60XLvlJE1Bjk53Jfs+8CBleS2qUouoqxtD2lwilEssB6qjJgs7OBMOVC9SfGYH
NZecxLY8mG0050OlXG7Ua7hSHM0XBiuvfra7I8cv9ZzWd48yYjluk7u1Wa4805HOOqJ5PoM6aI7G
I7O1+uSEeE46ToYjoxexiegqXoXUiyXniax4BWoaT9q3efr0ksdJQNm80bV91qadHHnURqs2Woua
juU9oXCqQWcuvI64zhfeecnVbYkkfx+a7RR5EOu3ld46yCdYkRSn0r6+gzgz//L0Ju8x36CDb5bI
eecBH4/QLREC/zyTvdyGmaEJ/BHnzMZnS417N8kqfq8WO+mmeXWKwKv+8bB+bD9saKXRKY2Lpe1P
1NE1XD6eji8kVuhO5Vi/+HVzu3KyN7lH1XeXqWHXIF0qqqsRQS08TPwgSZK0dqqZHQAq/vKAZLwU
X8yRIrDGFA7LMmi8J/+hgYs/HPEUmU7DwRikMD3CJlHOSfAwb/66/9EtTrXskeivrH9jLV03c/XQ
3BXUmZVMIysS1x63KOoAev5HOIpnvbCiNTJSREk1YTgLgmq3nBFi7lKloKlc3oTj3cMT8XH6hr7v
/PyOfILJE2B8Fw6Ohr7+6jeA7sE0WLsLv4NNPaDLY+PZlPZxrHQzTQ/ED2SNDfEIeiaRTEEKneq6
eeD3BaSB+LRn3IrhR6wv19QjbQTbtZ9C8Jhx+2oBjykJAxJNt3YHs5i+8Gt/nOX29TEqy//hEJc9
3LB24KCFsn5fBChPVg/jb/0w4nfIxlboiJXX1tIWlLVFRPFXjnr4AAyTSftBlPs7Tk04T4uu8kJX
9YxRi4q2CtIbzXG0qjbOiw35tlgbsUx5K/1KIdZ0+KCwoPL4Pk5nPDvMcREUOmgkXZagGnrDtSet
SiL59uxkiO2d5XSeN0XCaG0wDiknk/errUklsYFWMSugOJpcf9snVh57q3y2qG2/BROLZ8EV1t+A
8hQcJ8gaBqXb+qHwkOLlOIkLDFbbPB2fF6WvVx3fFf38TVwpDD0laRl/3a5dfR9NNeiaecSD/PQM
1EL87mmhP+7J43BWnvjigItRps1DrgF39XccNJssVuvl4gwCQ5+SpS9GH23e9mVCLoZfr/2nu5mp
IUWcJi2jt7WBuymc6dNW1a26TCEqEZdFPk65qhwO1fTHWsUoHbo3SJiLWW354RvUeSYNvgwvIsG+
5ydhOVlwZ4jpel0PxSQAXYCBVMIGbNjkU1aTlum7l7eMfjxvD7G5DybdIfavN8WOjBr7kQMxN46a
Mg+DJ2adKUqlNPLwxbh0f8bxXO7Brg0j/vzQHEzWWt6ShMMDCQYuu840Ltglk9sX13hwDVfqYlfP
hunKxEnSohHIbpuvtQMbdiIIgkCKpxcPe6JssUIPNnLJoT0sGztEbdGRNmVLrYbCG35Y562hp5J8
/moXsVhx4uBepaiKcmwsmVt6UbrCl2vtOyRm7dgtEtGNdtN92kQXLvO/B9GW5Yq8t0fEhDbDfnyb
wXD2PhaFQP1mEzvt1YqAGIZoYQ23NHPO0jI51dsLwNm5K9GVngtfIX/WzQ8Hp0ornTGoJAODn94K
GM4lwGW0zp9oM5srhy1aoMBgqwAVtrEu4dt7jGIkpVszyXM9Vzr0CM0zTM8IAi0zkFd6mPBETLwg
bYDJELD4GGq9v1LU7owDv595EpZgHcJw28iu7p6+eBAAOH/AEXBDeg8Mlpkg7vGJt6qn7egP0v0p
UC/LS/TArHGymOsiP9dq8rSFPxonFCUkV7T0U6SBz2OQB6N9pgmxf8q4h9H6H0kHQpO60gKP99E+
Zim8C060jZ9bp8rGMkgjXnr9GsDQq4BoBIM0RnD8rgkUPz5QnpxGrChbs3k41iZ76CYG4rVB+TNO
dV1aza0K4QXiimy9PSwaf1dyoEWNy9YPhjsXjsyx8pwphDoTA56BRPCP38HSqdqcZ/bJ7j8q62aM
CmHE4IS5n+3FY59+N+IubHlGHCJXn/m3Cz7i/3Vuw2tlKHP3Ph3RpXAMVSRI5o0MKQtudSxQk6kb
dupXhsbydeP3qOc8/Pb/bY1BjfFKuFrZqmafHYlUcVgiMomgThNDMIJxRwdKZ04tUPEkqsGXDM+E
0QzP0/KfErtbo4lw+FJpr0RMcGDfJh4NnvYFZJH6gUCyQIxeIYsk9bsRdn/H8ZNcrYYWWZN1zs30
MtTZR1zd8fxP8CLnreWDD1nNRuzRLoGTv69BZ2cvnSwQT6Jphr/uphbi5jeISx0OOCDVM48wz12L
z8uw55vVooeEefyQTzqA8XG3hPwj1i4a+xyA8c1sx3oiz0EfWaBMVs7zt2iibl6m1yJ2RhvJB0QX
WNz8FSonaSaTbnELei1UtvT1Ch6AIWYNYCKJne2855m9x7BQgH4vAwMoUKAN8ccsaUGLHj3cnx2O
XvZrHXpp44I4XZTrI8OXgwdxWU76S650c7JPBCPF4v3bu2k4aD0oElPFJSsl1CNSeVo+iyZ0aAVz
Y8fXc/uIiplB2jKOhml7FCVRIQdwi9sg+KYYypV0r+kGQZhmxs2hipPlHdn78vSCQ+hjldMEcCEn
uvAHhzLrgZ5d7NXxNmW8mc9xGSAC89ARLCc4vAfhX5UU1Ol73zo8oqSDF/HFr6Ho1yDOQj0tIGJL
JYUzIvHDm7PXAQ+D5Xqp314x62RYdphup6LozjddKsq1QtYIGz5PPwkC24xLxdRbyOluXFqolk0S
RNz/Clp0RUbi1Jd+mFuWkGqhcAubQYRGGCbT3Q+/X/i8+2EqK7GyvOttAQk1ieXAgoHJu1ih1Yyx
kekBlgeUlzwP/qGz7LqT+1IShFydv+zpO/mXSvLs0HzQ5lJjnDQJZqWW4f+mFRs/Ze3+rdjHAOzn
OOVhO1/Ft86lkwj7+TzB2iZnkd+ZfhT/icxfA9a3UNowY44+X0nnrbQwFaic8vHXgsVZizjvEvBQ
hzR3ShFGjxHHm6l4khigi6JfSdFv48/FPaO4Xlq5xAEdohllrdmvkpeVVi4er1Iwv5Wwk+Lehfx2
sDnvjNJegBM34a2FkvkvVJDsg2APVhn5wGltHPnZIJyrtH/BY+mCcVv6gp7juDcSIS4ICM+PLsEd
oEk7+1oKcceJcP9sen4Q5cYBiNYmh4anjyh0L/JwWgtOz2s8yQBzQiVvvj0TsZ0ThhsKDrgx+jq8
7J7edC135Fl8pOl0WXa7u9QCXJF+2pFC0x3MOYup+2nMvsR1WBbu1iuhdjjh+L4NovtS5cUmaHTK
KTUZw5IFgpFP+KtpaWXXk9jOkpfosaV0lSs1PPZe+F0Z9kLOHPUhDlmnD2YDC5RFP/QBWY/TKiZw
6SU5O9Mje8gbpBAnksuHCJiGm//gTZKXcEBRSmF1HOqWUrz4PWwG2/+DjZJFaBJvOp3btb4+e55r
NgtEapjgkESi+/2S9Dhdc1UmpyAEz7RoM8VjKvlKuAp9KGL8rtHgB935UU0qx2Cwd11dNqoSjZv2
T6YNRVCbX21b2NMFWO0P094LwhvUE74oLGZalSr3Nssj7UXYDkUoP0aP6RvcaJvAq+w61V0FY7Zm
eho9qLfridPrfeug3kZjz0vtve54IDnZ1t0L0hC23orSADocY0v5xayEBBspJMay//y8T9lJcUtz
Wawjw42FmctCQSsnqwPngukuCHOz+LfHcgd7YfD0tBCuLIXgoi1pnhHA32JObLjtw8gA3eOkWmgf
2KVzrIuCcN01kYPyk06z6totj7NAPdu3dMelm4Y3tC288RDV+U4Vv3+G1YxMaReOpJL8G3zLHxs/
uM/2TNRogCBSetFbJRx/dOdd12+DYKIdCxIK6SmgdKHHS+U0NQa3980cmi2Toy6tu28QctkmG8JR
p3HKSK+o0eOK1igGDFzi05pHtJkWWVaPy6bfLmXuJFf0IhJiCI0f+o6rnA5zfXSiXT3QRfEa/WTl
h/Fjs+VaPrQieHCUN/SQ12/45XoJFWa0Q/FULG+HZUbBmjrNqgSAyCzZEei+n618LCPdzuW7bxDW
AMnddu28E7hA+Bpu6sRPvJE8V+wUhFFH9N2ErQqdplq1OcYnixk7U25kqs1wjRuA/98IasyhkQno
xQkXSY9GtLV9p7UIZ7g69wg2ccEHacHZW32YVzzTjFUnMkA0gyLl620CBvnk6MkNRS+WAwR0xJtZ
vAW4RUmAZVwTSqPetQqpnNNupMeb45LNOpKIR8lpmQktP5afH3z37u6+ZYMOGAVCbfMI9M/PqiSi
LVwpWgMs79+XGMn68hwI/PFFMbn2TgF4dNViWSB0+AMCBQarl30/BTJSqsiCbSri4LL5A+p/Vtq8
0C5oPgFC44qE20csFvuTmUvHbW7xAyaKbOtxfUOtKMxI7D2RPUbq8Isl44hfit+oqtZwJ2rGbGZP
DT/m4T5QNd1wM3wjHqLadorRYfn8W+4D/6rk85VGvHX2p6ezkROHXWq0uwRXBK/ulW+5q5riRd+I
UhEg7tN78VDOv3DeKEIssl5kpsS/h4RHVd2DjN5Nw4ccfWMXPNNWN2LzhQXyxtgCd4MX95Me4mjx
566WRqCBPnZ7F+eRAQ0LRsf+S3WYvfrWYk3z5x4diWr5WjLntLFW1yJHnXMqXlxpKiha0KBkIY5J
qEpXrJOLmB8Ye8fkwQs1m4jN/TwV1OXdGBNFSOxDCcai0bgPFRFPM+SMjz7VL30e/8mD8tFFmW8I
BzvzLqMbYcqHB9MEFTyjS/O7QzIl1PSdoXugR5E5R6/eUKn6hfeBG00cPpSRyZSv1jpyBFvLlURb
AVwjL8oqCzRwc8HkYbMpGfwGEjP4uGOYC4hhz95XmYfMzkqZ2bwsxlFvvdzGAz3oXlAq5GJ+XMyC
3ZYCeHo7CP0McB387dFzX0B/1FZBNgwzbtYQ8hqeGxnxQt2E0ZXBKqHKVVdFiAAx8krsm5QiBdoh
mM/qJ9hrY8XPA9n5dvXpq+04mr292JrCQf2mm8n4rzJV8PM2pin7lWhVLd5jv+Wka2kYfV9hjFpL
QYsacKXdd6A0K1Y7BVAhg+ySimnqMne2hlg3IJiuepEDsOivhqLDktLb3VcGaJXeQwRcTV4Ql8b+
ogs/VA0y6xPhE59EbdOf52OjBDkaNr8wIOqhaORJ7a45iRmh8Bs4zDLtjfuDVtfhdyeFDorZOaOp
nZLfnyQUUbqWUsBET9X9/NeB3PJBA3vv/5yCFktyC+gTAycqd3i0TgYPvLWNKhOL38JIi7/wgJr8
ZnP8ee6MRgoCDtIjvDzkRMwQoe9XExHtOZFCV8prmbHUM49t0p+dOWchWAPV11kqU2XYLDyDH5Bf
q3yQ+ui9S+e9H6bzqEh8cOcMVcQnw9lvxReqUPVZMARM7M2HumlHWKg8+HyhZv09gNamcmiNobxA
WuZLcAyITfAfqpe88/LnXqI0eLHr7oWtKVNY/l5D192wGOiM7ya1feWBHqXCqtwaS8FMUnuVwkml
itToll4ZAHHLmd0DPohRhscVZzaCAf6YPdXo4tMAUJq6ApK9EH6Jkm+2CTkdGyDuE9NRIcbbXIky
vG8YK4OPrRCqr/DfHGKBkQUD5vnpybx+NcS17Nl31Y6nFhjQ0X1bncsgoG55QtK1TWxQYKKt4Oj6
gPSUGNrXHT+RqQFU9oSTeBUvYRObFNymdncG0o5axaZ9704GdGyjoBDFb7INtCwqOtm+8wpD8tK5
7z9zwJ99jIwwRzrifDvp63hNbBP6+Te4M6rqMJSElxnLBLpW2gWwxYSmlb0srFEkqK8nwbRPPQhm
q459sORFuYF8qtScSkJPamLlhCJmpM5Q38r7j6m7m+fvARsQxnm5i3GYMMkGLQLKfkR2vVbKScHD
CmJCvkr/fZ12fLyQqlVSFRvd+TVpScsrEN6tNyVV2UgpeAU0Su3fjjbpM7PRuDmiSgp2Sx5KMuum
FJbY5cge8zgzwIQbrqnR/gxHXgyrbab7Q10cPlB/ZrBd9REoATdUwx3QRzIoGZXpv6tUgR5ecruH
AY7n8d4uFvo/q7xadFVNqRp/vICn3/6pni864lQKaBC/+fXYDrH4755nh26IW2JGDxjGEAYf0dJE
lSHwEOy+vnxFNrzwqVaXnfDT08pFAXnDlK8uYC/Qq71SYVNYK6K/ODJnyAgvVKiAFE8rtMvKRREy
8CjqlaPGRO6efHCXJr4NtkZbPjwGEfENFgNHbpmbt4imEjJFKB/oefScl6lxnEj8DzZ8NpjD2zPm
XrunJv3O53H2eFjIfw08C1mvyRtWhkB+tVgGkkwSUvu7GwETf5KYTw1V2LqSQhRp/641eJrvuRtw
SqB9xANP9dKKdunT6hB9uJulYvPUYEg/ww2wizSty5iJ8Sc7Llm/G0Al3o4j42C1w9p7Cj7qEBv0
ZZhLGrp5vXEgmMe+gu/iYgItSQ8bpfSl/AWOjNYzLDAqlPYMJZMCSfZEXc6RfOIPnDDjhT8zHQ5G
Jy1Vbm7wrexIiTO/ooKR1SNQXHZ9SMy6iLZFKgIer/yS9lYoNjDnzLQqUs7U4WsHSeJcApPHDjb/
FxIyyulBEoQCsci4xgi3Fl8fIY4hISohicA2vNhKmWZvDmGaFDpX6LZweGvx+wIp/S7sCeSW2pq1
wSHMIci2xkOPuhCHNs2o3EUivkmEMiWPNu6tDEHXOT53+ItLUEpCCnm1vhEA11xiqz+rUtaidC6o
iqTM1LhYCBmxV7TBqTrghbl5KV28x3I7IMJcs3JNPr/w8h8jH6EYltxrYctMtgQYyt5NP0uGQNT5
28L3zXdZ9t4OKfQ0CmrzG4zBB4SDywADeO30/C1UKf+D86aZo9oilqTQNfsBD8Y2X7lXaheB2ZVq
8aZuydRuFRjANLdygZRBbcD/hUMfJYx8sqZ365VLwCy0dtsWMTyPZCK8qV4zleJW+VpzTTN4LyBm
Hsfd3Kkk5ZLrsuv9S/fSLN65rejHWbWHPyEBtPq/SAn8Tds7dfeq6lrYWdyXGeKTIvl5IGxDiDzC
UGoI+buRAAnsCONl6pncL+CQ59MxiuOePDMzwvFXmZLe6d0/gdkU8Zp4KZtf2tlNQpfkDEn3oZ4i
FacHlcT6EQ7XU56jKE+ObzVYpne4AaicdHZT2Lw6XZ/7P9lSvYokhGApG/heiRryzOaQWxpExyxF
b4s/ISs6j4JdeQSUSu3u4KKX3Qg3HJENrl67w0VqaBm0GZlMfb24NI2MnE3ITsZKF49FMBB2DKw9
Zb0/bqtOy8xYLP1nZ6uU0gi57W++Lb8egwV6z46DkNudb7cUANx3SMdX4l26TwFNjvGNs9i8w01P
9yYdnjIHYevZTtJX5Ky9THYZD2rVxEgsFtRXZyxL/Mmt8eBPyP0PRFMYZUbS80IY4saTFY90lDj8
Ec5Pt0cZFvZLrymDobkQ0nzNSEH8y7us7joJmei9uepEtqiXwyZdBYq6joiLd4kk3NhtF82IBcxp
qltNMEKkaXQDwZ00lpLHdfIhga63F1oMpw/PP5t+OXRgvAHdyAL8YrJbwTfZ0VVWcE2NYvfoTy2j
LNI1g954EV/zFXvGGYupwQuXln2NFt2mb4Wc2nnnPVpED5SxMmqlV0MlxrwG2l/Ih51Sc7ydj2dy
pxRYm9c+r8NqSxFD49dmX+cSuyZdx1hL13UGV5UljsBVha68xcCQLil24hIF0QIBE0uo55QPHqs/
jUdBypUiR2LeQevB9Za6Te8jUrAOB9PmEqPOq90qNVGsVw2dTP7ibF5HOdPFFP6HFouk2ivIQNN+
mjGs88yEqbDx8sDt7q4RLDZqcWPwW1GKIwKucv2JwxpEdhfIzKsikYZnv2HwIKFj4dMxys7COZSh
b+9V18R8MKp5fgm43O47T3tytarxTb1Gp17OFCRVkgEnHrZ53orrUNBrJ0YpX32kwEO+s4DqXgfR
TIx7hutIEnHQ194x92JZY9+8e31E/PfLAtETjFZ8UJTNa7xuYhLHOJKBd1BpTxI276H0dTOdx3i6
fGPBlQlzcTcQXShUHf6eUHaP1tB3atOvQRnGGFLHi2F1rRmg7+hAfMf/VeKDaMOuN2kYa2Qbo+0i
g8BrAM5aXXtlkk6HfU1XLctQPCD7seW/1LPwQuOIAelgiTZ06SOaxDajvgNSqtSA9wRYOPQpLkCi
sPkGUgrS8y/JpNtBfS8SiilEVI/Ot7uP3WRVccyhXSCyJH1IDucEhXXKdmzJkHXDrJ0ZUraArtb0
IJjGFUz3h8UZYbfsdRIlwTtEIYDX23eWoHCpLAg0ucz96oTiaQCBFGptA1gSqpCELIPAXT6o4z2S
pIehVTGQch2V8nnHBsA+fTa88hhs2Svn1XT3W2mcRI2NN4JGTOFs//hwI2peI00OTyI+0fOSFTt2
EHgO7a0wsF8ecnjBV5bEfw5vmfen1fLgPRseod93U6RtxGSvZ+cGtlRbeVtrooNkrRYGy0E7b/4i
Futk93uiBqCz4D0R+OAL1i9KIV0lc+X6Ol9GTAfujp8+36NkqRoo38TgQGOCKEa7s/V0K22H5b+B
QaazK2WKCmgyuhIkqk5AdwjpjhMq0yJYiAc+MeV2v/KCP78BtXwJLbKv/MfHCniETpi5GgF4tr9a
ppTx3gj017jaQk3lPkTTG0laPfN/lfpseVRkS5nCJrZgb/i1w+e4qLuziOMOeQIgP5wMs1zbhw7Z
jmSB19ad6f+VvTMEG6AHKXesBIBpVPanQFdnm7G88/QSFqbrS2U8z1Z+4HLj5MOO3wwozmEAtuMd
Lv3h/bpQDRTChM1YLOdhyrHNl/sAI0R+AvUZ+EE6SOuGrfYaXkDW+BeOrPdkJX3+50p9n353ougU
riQpXptHmjrz0tZF81M7IWX3xXjosij888U32RF1RoNy8eMRtDZ07Qo/L2pBB+OwXacXjMoKU/3n
Rq4wj4HgVGpTbsNDbs/fB/gSGfkMTA11och+RmmCo1iQWph9fNs6LQbMeAFI1Ag+o3QEGRhWQ2lL
k1QcCoTJwpEDA7N8tRWQDyG0DKIr3sr05dIKudqEO6Tr9A4Ng2GgN4UbLYu38q3aMD1EBBustgN2
t7jYYm9WSr0fCGTLl7ObBGHofjNOgNUWOjUVSd6ifSoi6DAO+6HM+uW1P8sCLC52DkMwwlSbK45Z
kVIi5LJJU1dIVbjpD6cKlwBUEmceGXQu3T0svQfvgBG2kg6E8b06QKJBrrMbyJuoNsTa67+lEZdT
qoOI7B8n+Bg8KWsaLs0ePFPjyeh9N/SKZ0bcGYO4smzSTQBLFQ7/z8SyX7O/SQTMQO/WpTQjBz3c
S4D4acxZr9ooQ5gdjiibebLNJDhw8l8z6hx6yTKnHtZYSzWou6kIqMPTikEdp0qjTd2Vlw1jpPqY
+xHNwVfO4UWXYpL8R3g+ptjkvlFQJSF3Fc99RqzdWDSPOU4FKXUSWwxNHqtK7Rla/Ko6x7LlST4U
lsdZzyUSvFHLt9a8OxWTu/1S+vhrom5MndYAiPuwEaWnt7kvksnE5DGmadCJ7PZpfEF32caZhM21
ZmAUXnsll6L/ZfwAVvvvXM/YEKayhHDflBOQQPiMEtPgGTZMg83HBj6tYtv4Idn06IF2SBNwzghC
SXRgoYGfHjtgSuc6fC8PIw+Ph1h7xcZs9UZhmJw8RNgBR+8sfqqxnI9XUJ8aUi6LWIjgCBoXDjM1
O/rXQgD5j/6bb5eylfym4le4qq01zIc1tPzuwHIPXXbKyCynsZ8mSj47Kf7StxgeHfGZzSLi3bGg
ETmhAA7zqAtwoQ+dqtyecVp42PlDPDJfp4TPHitd5VSc7wp6CrgBuZkWHUgpNWDEZLoPODKs8RUk
4Y0YbtFhQbiLgEMgCEFEu/u1rZz0kx1Z5ziVgVrYTjd31wBViYPQoSZCJPN/o/MIH0q8bW+PQaZg
+3Cwz10PU1C4tjhvO3XdZNPEKFEtHrwHFoyli75KY46suLCzqgczB0bR3HPY8hfjmjL1JiAPG/u+
uz08P1kz+gsD+ISpBFFA72hp1vRFO9JUmxlXnFKX12oRf83+wC72Kh/4YVrr0QNyP/VIXvDz0Q8O
ujAqs/l05kiPv/rkw0GEEAC44xGt9fWiR7kYsZE3DPvggN8CwwZNXhuimBa7qrdq9v0FeRIkSEQx
IyIqfn/rFjilywlKF6UewPytor7Z9CO8o0Zdvp/4tnkOlySrq+FGnJc4N8mCmPGt2+4eKFWNtaoL
x5nYehESMonZpmJHvstvBfd16WCwaxR50fzoWqIqN1hCV7HsDkn/XNYln4eShxzE5lMOkjkyrOTS
zmesQByN6K0kM1FqBXKsE4Z2utNpzZArjpz0nFh7bVWq9eYNag1f7r1ZtBOSpvCsVuMdwPYkCuWx
0uXryBLBInycSoD03rpKo8svnb/hYNEAdugTi5JqPvCjVbrcTWXiwDRnXQPzShQzKkUwq4x1ZKSH
DoX6QpsAgmrvu/9MkYSOAoNpePRskCQhzjJuSTJN3oObiBlNyIalNlYjdSHyvMXLl2MAZWvywd0Q
le8FGpk7llTceSMN+wsiuyQYi97ZUcmaKxkNC9Ub0JKB5taODHCSS9HJrZEcM3wxai7z8sBRfQv3
z13jfeCR2jE1E9VRUfpgaxb7BON6WswFiCaOzhbhERqIUQbv1vU6X6EX2+x0783wV4L/rqBOY5tS
9f4MkVeeLHdsLE2JO6KUF2LzSy9OuE04NKUZS9wDfPNW8IKLzr0XA9ORFjetkoSfBixS6smPVylJ
Pb0sTSEhbYX+KAJBD0Ul8nvI/vyZFUWut7cuHn5MFN3U02jLIiFymtslMw5KGBCyp+REfFEwwFOZ
1nNtLCFEBv6t9/Gp0/R4gtlCwH8YlBHysboaM7q52PPsEcrMtF5TSGNIyYcSFEwf84M0gGvTwTgw
jiVz6yI4hYX40drWY0JjNfPEEUoCMHgBsUmVloA7ZF5EmQ3W4iJhCvby0BN6RgArgWzgz5NrVck1
bFQm4xdsawFM2gH3LXylYHd1qVddrH+7Vz2iH1XF9IQCVG+Fgbjxc1d5Mbp923WnqMk3duNFhTXk
oP0JoaW60/ZTwQ0Ne2tP/X11nnQFutD9AqtgRx0BbW8lw7vtmLuYBkUukuILPpck6kAuEodwfglJ
/gFxzF775tWcXgSR5RnbXVOdcv9jaM4WOrqaOAK5k8a3RG1Jcpsl1zXchsKz6pHs/++sxN0TwpXp
eCqA9BVNkmNXgm58N4hMOnOtnPMznmaI0l4kUkXQ7jn8WebiPZu8cBypIwRrbjMdos7jX/HTAIdy
M/YrHh9bPcujh+hYbn1+nAys8yIri6zUZwjBn29qDKzCXeH/X58MqRZCHbpjVOCe8jXffBYx2Bex
PyacQ5e63SkstzPAXcaeW0eRu5B0gbBFcaaqotaV3469UO2VK+1s8W2cJHJhtnvqXewM30mKU+s1
naGx934tz8mVN7PPd9pEJcg24nAOJzhPQI8mpK70BFmp0fV8dNw1fc+fTsrGQ8gFFHEMU+qR0xsJ
YtqUKY7UTWwjFCFJ4pCEvqJaGeSkudc6lRZOdrnn4iN7uVwDQvdWDTCnMNJftaJLdvxomp1W75gP
whtg0eGtR9XwAfoYamLqisgiMnqL4aKsVj1rZSrI1Nw7lTT0JzMr16un5MZ4sirS9l56INHvz1Cn
Es2CORr8GCU3h83DrV4kn3oNPdc7Hbj3tp+Arr0qm88z8cDLT5F4fG+lHFwDjUL8OVw9aRwYmn1h
tIdtbWWDeTa1POEIviJ3WtvUOzSyyBpUcIhvWHbYBhq5Co8gRSwoEr6GMnZ7Uq2vV2HPSlC4Yy0v
0LOZ3h3xNIkfVpGg07fpYkLSP3s5Nu+ECghAUkMJ5rPa9WOfocY2VyhxKD+8eRR4p5BVJhNUUbpZ
9R6ENxrjlqWbK9hXL5WFpuab985+V2s8rMwNxUqCLUrhMFHrq5QGSbwkJchcl4gvxNcNVfgHc8ox
3BTzfxPKdUxezIKbeXQyUbWY58J2lBmy06mQmS7PzjE7AUlk6+3nQFcNqsbrk4xbBZ5mpLCtPNgY
yQoaS5IjvrBUm/wO4425CPr8oYKSnP2E4HUnp/xN13EilgvTA4oQYRZcXKUE4feH3O7ODDePxTho
tL1u5pE+/MeL0luraCkPiqL56u8OVSsOJul08i2tSO0MtXcc5WZWezHnWE3Yf1+Rc8jR46cBYnLB
enI2RXbKPdN5qHEumFMfEdbS7rfV4cfJ1iiyY485cARgjKd5ReclYp0r6rcdQzWhBV14K/bpia4/
ykOVLIFZxewA5MFqdsli9qvhJvM0ysfcMDieCyW/eLeO5bKWan0NRqqPrm2XBA/ZXqVzXGNBIG9G
F9bG+ngaqvQMLkMtW9AAEmTq2LFcTGMh5h6QqDccfwZjp5DRp5+i7urr8YEhZnJ++0TFBvwjtljG
/tbWrv3XgLqgYcvSbO3pwdvofRvus5RJz9CoO3gU66r4sW1d2ojCAalehITWLQtrNA95VIOCSQkv
yAiZepDhdtazq/qdN4sDUyJN5vzz8HwPJWkvTQlhDIpfyZvWdIzOfQlHmZDLJdcOVV9U3i5OHQQp
S2HoTxjNIQhg9S1UXfj26DuK/HS1xEY+N/bU+D6MMQiKyDqY48yLo/Wuxwl21TKA+Piw2JeJtzMH
+V2zt5kS0Bq9r2aV6RtWzy2xHXgfCse5aJfBuVnWOSVo208aesqK36ByAaYqyuu0hkzHbKrrZ8Vn
lHarLE3f6PSI5RrWH97l7JMm2/6lWja8fc70VTwt9vPlik2PYueUZ9B5A82HP8jFbbWHUGylTWdk
z4QbaQ6YXOqt9HgzhLgT7GlNmvbDwNgO9Z7TWeFbsJcHXw1WC1d7JltUwIYJFZM1iK7OJOfq9L0B
yQXeQPD1I8CbT6VgQK9bDxmKayesCbND54BuVhhUDhrdIyNUc9LnHkjlZl5mIz5n3SWqppAM6xMc
xSi4vOtxEMmYYPLbja7pp3mDo2GS/2dkbd5fZOIxV7O3cwsq+iRkxn6dWYm9MQ4s6ODYYF8XHKoS
lUNc0yEeeRYUvVQUrZEyodv/xNm+KOfwLAz/CVXphqpztfYh19AF20zJOaFebfOni12ILTsLBn5S
fycCXyJOfLep6urnJ3tCirDqyU41zEWy/fWOhxw1xgQ1KvUkhb8WEuQHGOHI9i6T8wacAe3U4BTd
fHRAUWebhDiqcz0HWkI6Ks6GCrBu1DrBJPgjZxFREqHwRkno6nNKoZXurJvHWZ8WtH49wM1SoWDM
CLqRD9jpSBgPvjoTg65YkF/XaNKD0IMrFA3mGNX6FcSeFEo7wqPuMz0ph5dOvNJJmzkYWWvHIHpY
hjEizHsEHv+3eBKf63UO7M9xlPODk1lOCkvMOsor/+SYR93FQDhHOIYymVqf3INaF2sA+BgS+Ous
lZSXjuaWhaoIW3y1eeiLlL6BOsOnaaAv+miJDqqJeaDv460yDhIqRPLhj7R6pbuaes4aEF5DzNPw
3xVLpFGuRFkDCxvNWeCf5+83vAsp+uiozB8tj7VpAmGuNUh25Snqm1FI477Y8EFH8zZ2VBaJMS1l
PdMJ7m3o+J+faPYFTL0Cjm5ygO+S7NvyiYOcCPVv6ioi2fmfftQ/qn/pHT+nPo7YntDyROjIZdG9
G2Km30vblMxfx3Hbuu2QqY0esDa22tOo+2FJgU7+bqDwJTZFwpG0HrLkeTzSguXQlR88eegpq4Y6
kKOdi0EWyDArzgaTog4qWPal4eJQr8e8ZmwxCB22o8pdl9vBOMYlZNN9qNh66qgRh6+hgLJ8edqq
QMt6Wx9UXTpfmntHoiv/vnhkF3d+sHaucrD6kg2UAWkS2P6pUi+sAC5Ri0NK7OFdv9ko/YqvTjVV
pDSPy9GTiXAnseqRvM5+rFVjU0qHkvSHtWkrd8aDQlSCwM5itPYVDRzpoZo4hxzo6Bg3bbC7mhGc
dFB+u7WaTyIU0Cpa5wzgEReMISqGw9XWcr2dm664fC7+GJIumBmyy2nFH0pNz2+dZNs/N6k/5dhM
WEdZfkN0qT8if2FiX3rXu3wiMLd58j8dc/xGDd1KM+YlJ4ZH32gWTWZuEBJrvmf0A9bqulPxTgHv
NmlP/sLT2/Wx4AMfqx2ULRsuk3C5vOXMJ0oluDwYdt5vAyv4rlipUnTPBYjK7NzUufLyggl2MXge
UCt5wQYjfgTtGYASjLCgK0oAU4Gvhz1wV243qvcvHE81FxDV9lE3Luc+hndqmH9YeoACA1Nr/p0k
O6amxPViUJb5Q5Y0vq2wQwy2pMMhZF45tOqkBkGT5wA5eL0QSlchEFfXGH8+CvwPdet6zWAnrdp8
jdYUK3TE7SnVyTT88ggPt0brGLI2Oim/kzGGYbJozDgv1824sMobNl/Hp/PlAdi5V65RyacYGEQA
LXJwljYr3yCm39G5Rcw0y5sZoZayQLLxLKihaBgDCfuvLI8aCfgS9NXVtbKH3AIhB/r9Bkh3qAE0
DbwcLsEPSc8RsDThbpi7t7fYcexexsspewDGrrA27nUPpDiXU6JzgXdwjkbDNiAf4DCfQ+N2EzGl
UVqDsb7aJAUA9mNFzJq2nTOrUaNnihzjt91XfEalUjl7/NsgefhAApP1yuVIp7wWGyX6AKjsemi/
17lfY2qk2nm8sL6b0ZsNnC97srivUQX5/fmdN2V78Z8xivXZScvlKg+dsIpXQeGgd463p50P/BgP
dChGKCfmU5RLO1ewSV5XY/UEfmspdvW+dCxmoBr8xr+IiXzmq7+IEak0XBaPeyLqUKFXSkR0KOVm
L4Zq9cyT5vzQe6VHISnOnx6n47lAdR2jRynC6VXgVt0l8td7+mYhhkAPTiFtBezPun3DFE9XjoLR
uc9r3xQAVLoipNc561Lsa1zjKitX4IEOBR5ZN16uanAarepZSq1xCSO7rQ3JvSE0+i7og0X6adar
Krf9Jf3CHb0HyPvW8P3AnJEI5nuEiaWu2MfGzrf5N+ak3VkXtF4jpP2xpl7hhof9meBdfYoJ27rG
GZhOh9NkM6uc6pxKd5SuwL53jjRHN9PFJUKdw6RC8qMKmY3hl3pSPTmpxtNjCYHeZp3hKDuqLKAQ
+zBk7FJ6HjLfLueI1WarhzEqjbsGdDbuFD7eYkKTjcmfdElFiU84vvHsdAqMoSfz3XkiFZJwUiPD
DetBgrEfsgKFyQeOf/j4e1kgjGp2J8l88Bcf/AWpR1FoLMUocCJBMxPEVE7vykQubK8JRLC4tbP8
nXUGo+r6IMkOU41r2yEmRt6hU+QMKrSuvUES1BMvyRljNpL9pGK9ehuB7y/nuSbajystk5EAd4JY
zilbi5FYHRWtb6COI/czRZbAyN1vivxkoBA+cUacbd4jYOO6pCOyRwj+WctWnMClVkQUX+Rp3dLq
90vb1HfqFfFMR+hlBakYz6QkPHFmkNXqC3WRbbS4dHEAmR1i1qaJevO4p+t15cHcDTlonWNcbv8r
lsAqBy+T8xmsVDPLYAIux2bHMD6W00g2qYZjNy/SbbdhEQJgIA3sr/zdJHo6swx2ftu84ZyAKOFR
Tepg2lbBsM07Cffi1MsVuQVYeMPSClryxM3AFGPNKJcCtTbEK/Hv6pjm2/Xb/yki811sIEEcIYy5
QpF9vsrPnMonynPkwx/0fCDz9NDCDhHW8M+98p5gjVyGsIS3r/P3z49L76RpSzZjk6Peb+qt9hJe
qCwL0/rZHaRsgJLkbC5idwj4obxaQ2rBxYPKTLLDIrujuKz/Uc9G9IbK08/pAuPtbdSerbTYrh8Q
UU9t/Bze1q83aoQGK6ILK7sabtqTxfEaVrlYlS4yg9+9ulKjcb9KAX4nMdOTepzbErUkP0x8rp4o
eUS9qd4+dqTXsaKhIi5VQ1sTiE9yovOJ9V3+tYvvDEoxAsPn7y/pfAXInFVxSzKQxPLGeOgBT5j/
9HRfp+1APcIEn7igy3ovAk82LOjCo7Mmd/3hSO/sq7YG9PK1UR84srEdhA0tS8wQqU2g1Td0obus
RZc+kn9ubZAeHZVNW+Ki5cLBvAYgWzpzBfMwQwC9qaITu26gWyPefKdVyD+hRqZ+aE8vyjfs05PB
Jdzw+WsehbZalvN9Q1oFWYi0WKXU7S+TeIUjA1r1EfQ2+Q6YMFu59kAMms5po99VEOJ0/gEHewHK
tM9xIZpF3ZbVNYOIMbOheu2pq+JT/tqfES7xLZg3FA6UHgJLrEA6vyOwMT1BLzg/TdSv3LNJi154
0ILQuSoAjXyuAQWeAZMGZoFsDdWhvG7NE886lNWR3RAfrN27rV89N+9w4t+7nrQZ5F/Sv2YWXOf5
bw+omw1i+0DG2G5ipWFwQASkf15tAjNcMsZnLoC4bk3Z31cGjrfypmPWxDliIbHGgYoVJOpVjrpW
a+stJcT7vQMDWaBAxrGpsl6QkB8/jz+6IhKqVxmrYJ3JwqLc9agJ1u+1nYpJl0lDQwsLK2h5GxU2
ArEwtSpuLn5k0BB3DPHml4twTLvw9hKHwntQzVb/EidbXAcFzOlVaWfnCxY9J0ldr6d3EIkZ5D+r
kLc6FyzPlUKm+vj2vvVzAjJdHBxIoonugS+HY/h8iSvK/K2YAE1cbeC80+wKcupSsVsY0dkrzkZ/
K44jAotPc/VUuZdzN+GNF0Jq+cyM9YlgKPS2wM0f6gYNZu8SGhKt8EnjzSDbKr6NgEii92xGBeul
gEkXes/rMtaby6QWAW/sfEtVv/FJz6J8rC/+Exx+Hz+zHwO/79Fat+eugzOlGxCjP7MX3pOXyu9m
PhOla3zh56hOhhFtDTQ5Td2j3OtOXQoe40UHexHrItCw8nj7+jHQ0PjcGQsqdXopQno2/ydJvZ1U
snoZZVzznEZEXp9MXRe799x1YJwVYGFoqaGwY47qaxY9WT0Y7ill8DStIeeICf3FUSWDCFSCydFn
rtdPPzbrEur3RED5Cuf7GLV2/CLYukRdhMUohaRrz7IOTEBAd4iNNlcs0K4d61aT9V0J4+PlvGjd
kmjfRVteytQCspUsjo7lmnR0OZn4u7fzanm3G6NYCYr4Frcb+3PJSqDqC9iWGi+JxkTyqxCB69bp
trY1Gy8OqplwaeR3k8N/PTKNZfHsEfWMl+r6WnKbL6+znofsqj7Em33NAaw/h/HWLrgIWVhT4dRO
n8btK/Mr9ZfhxpAwtjg7nDKtMkz3X87ZB1tM2zeWAfYQLAaxgGkdIp7bHWfbs8dZWjUXpGtzfsSi
Klk1y10JTxrJoPzhaih6CaoUlo9u4QxlZGSoqj62Yh1iWSE2xK7urabqkFL55fknAc1734rVD+Ci
7S6Z64vZ5WiwYQA5mZX8swlgMdJzzSddhpLQ6hY857XPwrky2gB0MeXn2ShjwCbwUEcnq2KY2UYF
sFznlbT2Dgtcwa0SEmH4ZmNnBz0AHhdZ3JjSquz7fsKMSN3+eQl/D6n/G6ME8BPM0No+i2Cf4CRH
MOqzmtfRFgM++uFBXeBRI7TTVWrJgPnvmbBLbcaAGDS/2EeEwKfWXway/nZ7rdM0iO4cM9i8CFt8
kyTRF1Ubi0TjJGANbdFQb4VaHMYlDmXrRDEAicaG5zMSNLCFij6pB09rO6S1EqHjIljF9dESywqI
2oWnQUjL1mk8xx7WNodWsp1t/jLhCf/TAWs8KKZeXMgV6u0ZBOXwAr7q0I0Sv5irmk3uHu1v1WA1
2Jn0wloSlaCqAhMWoFYsRLB7N+L4moAyH/zM4XXcJUVk3/GROzRAE9u/8DCBQyN97OH7GOU3sFXS
CSqZDcj1x5kPA/+Y6OiJERqdxoFh6o9A8gkY63UrnYDbJaOF/CkF3yv6qlLC5VHel29NgKKOjoTQ
rWR69gcNnXy0IfJ8pSvZ+yF3xpvi54+9EJ/zqVXcHkewzXlthXQO4SDjoEM5IIDHbSfaoYRCTdrA
FGXoMtNyFnXzMA+ryGvb8AB3kcFh/3H3aC2/Pr7Xa3xctO6+5vxr0mJQDPfMSdON4k1njRIwcOCO
MUEu//G3J44254QJBKwelMSpKEwaobP63fvtrtHB9iE84N1v5n4vz67/Wf1WHjthvmufiYj06H7s
SJqSFPzSLTmnuF++VQgbKCk58/G/qdsoji55RTNNBFpRQm/gfvYS/L5ZsBHAoNYmfGzyjFvpZRLE
z9gF2BqRqq5zLhaHKD70SxswSaZ/dYoael+rWG1SYOzL04OS5x67P7w6rzz3pVRRsUlJnvJxNFO1
U6E/hZOB53EDwbc/pYvFEvEVveWgbVqs1T1INxa5ENz7wpYpo1ePhb36pyZzm2+8PyNj57atqcPv
yLti9bYpNWgWwv7lrso+Pc/rMuMGQBMXwjOctufTybj/eaao3WouLPRwdvdWuVzKDpfatIn9VFUH
eoAgVSRGo/BZ5l7YPLEB7ZpIUZZkzjPuK8PaEqed8QDBI+fvcTNnjUKbLdJ25AZmJivj/ddc6ZPT
8UL3R5ZqU6N0EafbBZGlu4Zo5xEqhGKoKRbsQU2MDY9OmgWN6mwfdcBurRd9Kn8P4yPpnVFrIKkx
ZfqEP7h51kYEytUmUiRqT/E3ZgNkAUmEmcEb+mNtZa4cVqFMMPJ9SCQ+UpHaEMasFX59yFu3Owdz
fhlApnRswwTGd/oCxRDXG/N3xtgfcZWZDLcAsgtCqi3WPPOYdquve7SWv6hGrI7vr5tbejP7mfa4
JtWlag1ohObcUgMFK4biRH52YS6Z0+CWMvZZCL2jZrELCOxkdwaqf3qa8+34fMKPYrS014tS7uK8
6p4Qdc6vKe6ujMy5FsnIw66Z+b4rGWtBy1dqCFwKvObF8+OKWUouLgdjSaOmA7xsYwqcnQx9Xt41
5Va/b2CUGRq+Zk6fd7V5dM+54iZGXm45xaD37p/pYWehiTOV8itw8mUOS03a1PGmjvM8NYZCNL67
nY9qGj+59eUVHZyfghy9KMOZi5YsLwyn+7di4kEGElq5bSoJFwsZSvJEhWB5IovJpmbKr7RzVPuL
ycppt4ZRchqjpmz+J/k3fCCl+PGbHwrNZkhdWPYyDh3H1mjyr7v6BQOW5N1OjMcWUbTcRUNz6IJV
oLh7J69cjYDeSUELiSlcikvFNMrvrdN54+7qBmVh7YN/M3fygbI+WRrlHkR6ZH19L3yUh8tdpOYl
cKTLm56Pp4P4Isp9b2cvbiXWbB4oxs2WfNcrEy9Rke3EeqlrRmcih0UcjHoHJotBJRAo5fi0pAG9
AIhAy62PpmlQ5jMs0FmOZLQsMlhIDUo+i45dx3Pszz+HLjsBVc7p5h7p8I5ARxcyUzvI651GswiM
qKA1PZgZxiUUcGXmbvXX1Om/CRfVHcFDFbu7IoSx4eN55zPRdWjIlwmH12DvDc8OYGZ66E0YQnjB
4hyMPYNev9E4H5gCQBYD6aEDsNVzgK6sFksyoBENo9omvC7kYW2jrAD0WoVT4zl4FJ7/YTQ5+q1S
tOEo7f7ZpqQvVVXsq0hW20iIE/2C0fu3j+MGGlHgclEltI2/7ncS6+6CDUaJag/MLpQAUFkheK2a
nFOEMhb5YXFqFoLmeV9QToqJ1fypdEMUFOfTpw7m2dBagbClBVu9qY2f2onojg4V+MvL4XKLeqHJ
9hZncRZlbJSA9WtaCVbFm4qOinp/k8UnbjoPmfedAXCFH0oxjpi+Iyps38odCePGpA/QQO+bgjFb
1pykPZEnH2iqsKvkLnruy9XzumiONK9wzmCZXWFqshLl1pEKaT3g/OFVtMbKKiccx1Tr197e3NAk
7v4FIwHqinIxbZM9A4GD82bLBvRKx93lJDXAREM5q6JRO0YFkgtMWQfVd/7kNOq2BrsMSqJYaEaN
JKVyh02H01wyJvgjAJLSjHUsjXiModgk44gdBnJ/SUs5VQ7IlN1z+PWEcp3FGpDKSyQCF4GfDi+K
BUtKJMsnBDE2/EkbmjMIDC/qiPcR9xL8HcJnIEPFImA08BFDJaW/NuM9PusUZnVIO104S1TpxI/E
F4DXgmeULb+Rla2kAv/6k69QmzzbVRMNdnOLo4q2cH/+mXOMMxIZpyHrV+1tugO0zys++NuJFXM5
4+uNxogkR1CcFRp5aC5wsNbOfmBf9EmhigKWGqWs21+wSSSI+YfV9cAQQQOI+0vO3heRqeINLSFr
PAhy6t5G7suUFYd3pgD0/zBtZ56oH/eY7OTTMEEvP9Stcz1qmwVeRp7i7TekEot3JuxdYoZZhlh8
tbnHVKoDGuIe1ySEiOlcUU3d5AhstdHfk30g7jFoP+X4Jv7gev3x969NTrDlkuHdBnjchlLf4Sn+
J3CKzvRqhwhuKS+n+Ah+Q64zm3v3GYv776NdPLtUWMslRy4g+1i2j2t+B24BFN8RNFtgVZEjr7SR
8vjaZuAnncwyMGVXIgfHtTDJtq8+NNZuuyAwKAndDuRXriuUEvUGEuuXUp2qtD4izZXlY0LzZYyl
xP/XVzGyY5ZN3LBuaUKwSaGf2Hj831a0hog2C5OcKPccfgqCtVverCmn8paw8U/D9TVsca/lIUbo
b99DOQgM7Bz5+jSvjEqkDtcxdzImn1BahaqqArlkfD0mtKQlAYQDU40hCo4UUbuU7+8DU0fcC5Uq
HZ43gbvdsR2ZBGIsiTtqroOZJ0DLZlq2DhZzWF7U0Cx6qNE65WeR3A/ZkqyVtj5XcqoBDNZIpBsV
cjtAcV9TNxuSGpXkF6TNuYHggKGtJ1c3sRkIvENy08iIo4/UhzTodX1Iwf65lHYeUpyaOK2IN1mJ
CyKHf3eM2dOjSRQVkkWPLwsaF38//pEEiq2zhijocq3ET88etSNAXC+Q+t7l/QOabZRKROjYdzl8
OSYnEyD+iOWUgOpZZ2cx51GVtqDLqwILTfPX0/GdBKHuzMEvzz4UQBR4iLuTUH3/prBdq+ImsHjN
qr5WmNtQ72veNarIeRORgO9IQA42f8zSgVjjR76BT+x9NHURVktw6zIdM599/gqjU3vuV7wH5zPG
gytBvMQBTSa3W2GttGgjAtxW4VN6knU9EiHTv9nJCwUE/cq2Uirbs6/RD2bQEFJXoNb/jNsL8FrG
uwOKQs4PBj2Wv4eerxPTzBXh0FdbS1/f5JUCMI6K3dEbB1catr5k4ApOO9ErFDE4+Fj+DxAgvf0G
5rinrWXPO4OHczW/x2b3LcWF+yXbG7WbpTroVR/ovkDzTAUmDhDpHTmVrcg+MOSzxfrrlg/g1iNv
lTULwfv36UgRrtGrE73bCmXEpuVLXT2q1fEbEI87QDPYTVHCPEOoBe4hYUn4K6xBl7dLvH6kWtH+
HY6fByMcpUJnukBbG5jDfnuepWsQZ7Benxt2IkQL8yPwb3iloFdlEW8wNE9H0BOn0EJ/686Hi5sW
oEedLnPJNQdDuXrhexUTvp4GhHniXAdFeHgnT35NIzl5TG9WdqeikqlQrag1HYctIRO2jXAF//wn
hEMqvXzrnDynPQtT3Y+x9+7Rkx4UXiMeqayCCaHhuYfnJc5qnZ2OpdjXwYuHq0K0J7cLzSCl1ezB
/b9qUceasQHEeBVs3B4zIvgAgD2D9X2YOInpvwyB8Bt0TCeSogdLLOQLsshqEPZP52t+86te3Nrq
7D3K2EFuka4s/rf4fWTvKbb2Y2hyRJwy3bkRGuUi+1yVndHyN4OJvn/owa6ZeB/gt5Aj14mciabc
ACFfeXeCwTN8F0y9id2pNl7wgl8e5ZEjhSlV0WrRP7NN9R2ujv91aFCuNmo9TDWptGS7QK87/ruI
FQK/17KhAyP/WdPFp73TNg2lEeECp7SWMSFfaZze2gk4tcJdmsgRw/7mFCEei0Ac8uxKrWG42u3P
t1ULdQzEL6fxOqeVNoyelCIIpjrRs8yTrpeeNmMnb9JDqOBDJzOvyuN3krxfk5tHfPcTSL4RmjLP
hV4Lum8FUkhGBUXYBeaq2LIDxhYnuIneiWvScEKzZaNrf6txvj9pHxt04m0NqRWG3sIG59KBcPhb
x6MQ9+KjG0Gi6lzlvwZfUlqk/du6iGQL2/DDCIQfPNGtv6nWUns4cq+/0dQ8WAnStizTo4wTnJje
P13iJgjWDpRrsMV9D4Qx10cxSG/sSRFJ4mkK9PYYrsbRnS4TXpBOiZpkN8CD/a3q2YmWHJlG35Nj
H+K90otgmPvRu29fOzB53dYAwGOg29DTWJv/wpZvji/HGvO7q07zD+4zoC6AplAg1jNgDOdXyS5x
HdpUoMyteZR7mQGQcc3VwpcYBGjMl0mbJwrPC/kDSXxOAcSDCNqydoMZa/AuFHojxCREu8pKY3CX
lW3f18hTMP77cAqqTQlWVl7Nu638BeFdZOgkvaSxo3wEufVX/+CPgywPVbUgQ7oJCSPx5km+FfrT
TI7SVcmXU0woqqhPhsBAQh+Jinjlq9lOtcZoElLzFKcn7afwqcTbmOYhDWQ8wNLoFR/7si0ewSkd
EOWiYCY5t6/wyfufiT5DnKShluW0MWpehR9nV4+F9F/llj8Lssqbl/Weri6s4z2oq9zab/xgPlvJ
CE1RAd2EiMJx/ul8gdEpuqtPH9kj4paLYns8wvNQqeOfDvrsemntoZLVTYPM2C3nxuO/RftcGet+
5ABQ7cShylIq/zZUbyRJupvJZzPyQHas0bl05J2A38LBgqJI5I7/xcX6wfsiKk9Zv4Ws1vrDhiCc
iboGNN6XYU45BAHqfBSYIOzASRXTaIXX7IOBT0GCIGMa50VC3aIIEw6Mmnrz/ec6ZFlHBtvIe5CM
4yldb407tS1gxyf6LxjXCntSigTSd7bPlsAGNZN0WBAce2hz10S4RR4daa//g7LXENM+8Od/D3fI
FGgpbeV1Lcub1b65YetMMFP4h8Z2Qn6/CWyd7K2aAxKPPtE0hRNQwFBcEF1Wx7mI+PMY6k7QuwCp
l7NAvporvRy1E9oZTeBJnuk6b7wx5rJiXECbUm/ZphQTVH5V5jI3LqMZL5KJ0ZRJtqYyVIFHvT1Y
NeRYHK0bZZEXppswJL+yMpQmSWtkkrPWZjp20E4vtwnOnkjD4s+cHxztvpYs9lPGoV6nyHbcsjeR
EnAOanf1IZQYhGc7vyGFqtd9X9OcbevnXmpqxs+UPEMO6n0pcaCKwR1FFBWe3HyZPV3zL2AycKau
GehWt6xAEWzwKpvFh9D9fz6n1WF6UFNQi1cSIsNRyZfjl2djdlp3gagRg7vitmf0NSyGUK+8IrzM
HHHXsUYUZrm0DVNsDYbi3NH4z+mYG0kj/X9oornvHgmXhl5xBlxfvoPerBZfl+KDcUNsluDfM05W
7348XA+ZH33vKKtrls0hpW8s8laTINTrsh6TDSzLlPiH5mlAu22aqib6ClYCydJRAloVgJjmU6J9
v6TArDBB1dFM1FgDy65rS46SZm/pMYRpiKfG957+RDfq5XdQKyMojIGSSHbbYQO44lpQAzCTVTHw
In5CNdwiavq73YxQBCM9uc18YCTuQ21KYL4EJkGWZ1++JyG/ztbmAlfaBarVGK4DX9Su3+4NbutS
nAV4wSlQApyb+CJIS+pkyiKuzYlSN3ld2qxQ6Mcqz/phmZy78RRI2Gve8+QuIY626PcPTt94ApkU
9XAEwR3uL/mayYHI5gNvg18kBdnSKGc/YOsbJOYEvbKdBbV8FRAHOwIrMB6Lz02qHrTJ8ma6h8PY
W5YgB0sQDDswJF5RO9yzgoHnjdaA5bYHSku9i1Ir7AvvfCat5cCKriYHXz6/tPzwX6HnYLYZpC/E
4BBqRgQbr96WU0PF7jzaAYuGJEt3tBI9B5/hc9hdY3xp5Z4eanwh1ng6uXWfpvkaR0C5Ei1bdGxF
gIjPmwab3Km3vGw81SWDwlOvwL64uVBiiw4sZIdE4hy00fdl8qOjJXixOF0p7D3hbRI3hulRw0hO
9J0TYP5DcrDl3JdCXhgiuL0hz8Xt4MxMczhrpsvYQPpT16cuPBzVRM3n4cY3LsMfa/uKX3Wjw3tk
bV5zGHBOjOiL1kiSiDnvMKgatkIyLncNBCiXfhGcPUEoPHWuv/6olfMc3cNnqZcCZvkG1TsrKgqJ
YD7ECu9pjDkiA7xkPcLGvS47mF4xWXM0MFEI9N3nYBB1wkRTvhmHltCsd8TrCRh72huXjefrupyP
xy1wCfh3XdENUdp4WUT4waFegZ0roZBiwaTICUIhcCONmlreqYRowEZ3ffbR2hv9rJdqQvT69fY4
gbsqRJJIaA1r9ytxzu2JZefXkEn5C0LIsKAYJoFV1y0nTBhOLAG36yXK6R7Fxsu384V3JRD7DBcS
Lh15EqLE7dKXGxfnBKIymv0Y9xVi/wlWHDKWy0MEAKpsMtmgRajioCwQv/A/qSo1pJ9ab8rU2M4m
G5uJ/qw8Xolh6/u4mtXV+X6bomnATI1kUkGKqo/W/DMCUCOarLBdaP3B99J+xmy0oU6dab1EvwDo
taUdX9qCz7O3g6H1fLZZEqNSYEx0CC4zN1adGqteie4P4peSqdLOx9/hGQrgN/0LIZ8D1ICWhYDO
coxsahBOn8Hy56yKZSEAm+4Vz5hsbHXBhOtJaj8qfCS9zhT1x3xby+he8g/LD7VZDAYOlvh7+hPZ
nvv1lKDuYn/skF5T4wVFJGnmv4qsRq654A0CeS/cu+1gRNaOjhTQBSaoXP//KmWaCEIYA+olKtuX
12zCHn6I67nqnaFbyA05YZW453SpXuvaHXdLepZlj6poNLbdL50ey2L3HZgoSs8FJnkAhxhwoi5y
lldHQacV0AgNT2Au6wsqIln5Q7PefF8OoVs10XB1/Uqq72xpmbEyEIyvFB73RWaAqMtJ+F17TEhc
mJ/MKVZNIGMasEwNIt9jVSyR6YgOhAA10ciuWJr0hcqPUGnmKAvOSqFCVzYTaKq18kyER8r8zu26
MHsiwB/WKgRlFV1aYWOgY8I1Xty68s3I48u5/CR8vXCXt6RwJeeiIdmB9Xk8N8upKDE9hqSpi784
BmuIx7he26vIdbuPpAFRs0VgUPoBkqvNGrs4r4foDmw2CTLK9XOeH7fcpjMrnSmiYl5bW/tXXYBb
bGr1Yp2ofdD3uqP9edPuAWJxl5Px6m6SSvBTU/8USLYdX+AishAPfLv3AltvIjkMCeJ1vf1+N8r+
33ehtHWXCywpp7Zq3sFXaeisAABIEmT+WGACfmGg/t4wpYtgDD94ZnC2B+mPWZ6gmdOff4zabbyh
n9LbF0Ij87O7zuAMUwDw7CI9Q1eYJzrjeicTYSMze04n8wUj43qs0sOoxrMDfWLj9OFMYcN/tyON
/aQ+NgDFId3/JlDnhBuR/HszolKqHHWMXMGLjyb8NLFkQiuLLGI6Q3dsxE+3c6Ur5IQzw5zeGf3U
15yYemxELhCrKrYlK/E/YUin+3ibS2YOpfznSesf8vhhXrfydHDOaTYvyVg6+sLXEEVXTfBpMSS6
u0ikmQsFFXz7uFXJcnx0BZlulUXpBAVr9+rq+rk+yBUWM2WZt9EGdN//XYO1j/d9rkGCw2rsbGOA
yXv5js/Inc2+jP0Su6P7PGthSIPPpPfN9P2cuQ0xIh4yG3fjfHCv+BpuVQZ7V+4tg6fcHIwLz21z
5lg2jcREE5MuKNOJGbxvUG3M/luJIvYKzljB9reaLKE9Qm1jthBYlb8lOKLYgxqat212ZxZ6C0W7
Be7G4fwpuZ+oS6kDUwcvt3w3uhK8GO1a5BkDguWvFLTAhNoEJwk97lzbRLJ2V6MTmQiziJ4UNqlh
47HrhBsN6y79oeIbmCA/2ddN4QrV93JK3LNL7ltuc2G6+hmfuEA2C9X+LydQs9XswLJgZHQAqEnV
8zYKvpjCDDpdx8ckRe1s0jJ9SYY7hHnQhYVZCrXjomhWxaMgKhxkV/tHbQDkMkx/wEEnK1lzTilq
Ia3ibhGcimnqu4lslE2bPIWZpDwcrkvkjEqCtYYII3neWNZwPopm/Sr7H+FKE8+KZxyghkfgj2Q+
ERGphM67aVRT1ONUrTUP/Kmvz9VwAk3KUw3n9YPIQBuNQcQ0dkSVzvqFPgkn7G1OwAuWkkmi4woQ
IadBU6W+lxhTOr6WsSpbtF4qYmsebw8BP/Z3McbvjVBykjHqxMuek8juufPo/bnOPA0vZRCD0KC6
lCGCfsDNWz9+DpCBH+swJ3rs4E35Q3NU1Aq4mva23A27akD4ZpYoBUtQcCw45GAq4seVAhIWIrIE
dSYc9twfkV62md9a3dnnxKCF8eSs3pPaocaBMsY0epwaYOOzNUGQNM9gFF+0yfg93WY1k3z5TJfE
s3kZ+3mYZ9N88q6jKUo/9BRQCiBy7phgL/STVR5l1FQxxsSUrjgqj2ArmwMvQq4Ve8ajaImFVbSt
+82SmKxMKcRpubmDWIYW5h7fGziT2mr5W51VynwejWvo2oKHJsGcMGtCzY+tw8sVTfGliX7U6f6W
5wMD3pYGHcPTAT5ZnxFt3sXFEmdmXPso4QtudoEa1ieA74F4wwb6Fr3tsTL2/CaF0En4txpy73Dg
rudnomaK5TzzPabPDo/Rgtn3EojuSGUXUjmsoDJp8b5dZUtOmBxyIrxJ1J7SsGOerqFzwjzx5HZk
VdmTEtbwH4hrk25bRF5FFNOzdyBRYtR000f0VK5NgLC+LWRskrSv0twRcm4OvF/7iY5EtmweNzI3
iVWhIuaFIr7L3VXsLgAzOr5jrnYVxe2AaTlwB9oe3rz4MG6tab5bi6a2Wjw6/oiM9VMe5AyB0Rmj
44P2VAg2gm6J9cQ895YA5CZ90xJsLq8e3FvzK7+THZQTWVbNqmHQ9UJhnDnwh8IfX3Nz7YJiViZb
hoRUR9LuN+sXWJ8gg0YtI9rkY/tnSRk/UAXzv7yD2Fw8WyC6w3C9KzfyIDytwIbFxHG2E0Zsxmr/
iX04mc3LYiCbIS7UHrLwFsdr38wmgQaQf6vTidKjG3R++eviSF2MhpS+of2xKnD1oFPamFA/FERP
hyJMtDJQnJuXaJDcYnB65JNCIVJ7OdfM88GOKMJ2r+tr+xcgzcMBFtNhvi8TKNUdBFvZHD15YyV9
v+NgBmaP955wcewz2X1RSpHBet1550rCZ2iS6tt8wR4cNnVlu6M9xdteXuou1pklklPaAS2lrm5Q
BioekjkBHYrlXb30A0C8EEAfRAIU/mZPBAfKjc5vTvPh5ESCXLl4PiPcBKFKKS4l5U3YuUCA+NfG
MwshLntQYB+7HvEWza2qptaCpY2pwNYnyWcG9mpCglUSJE02/ldZS/xSFZuU6LexWikuYoazhbrz
+hXBOGRPLjE6eIK2qRQbiVHtvF3c/X0nshl4fcQoa9ovWnrLJY+elRkaaqKSI6UheMRS9CQdiIn3
Cd4ziUrA/Qd0cXtDm7fcnRhhooAXKXdcMghUqU/JL4/Ih/VhuwGxN7yHTRpbboS+6sGLxLADq6F7
eDKmpZamLaBkS+3jlTLvxi4E5Y7p3sJ49uZ3D1NOErgxoyyDGsv+0aM8jWMaC5NSXVQPSiUnDuEC
UnMIJjuNnXb2TfmFbqEkfc76pqvZVdBPIjcHBhJwZ8Q/mD7m7/KIHMHkvXn0Ly0WwOkW6RGNP+aq
eSKrRaozzoCu3QwVh1Y3Qe5UeJN9v13CYC6CGd+kFO9sIjE2VFFhcEwz8E7QNth5wLWhBjqpj1s8
8fFaJhUKKoSfCrGrLWfWI0HcxPdLbI+dAGLYtYMYBtn4vHf6dvnhbFNbubg/g09rtSfeQpm2zuMK
M5LumrRsy9afIqjKYLChgqlUK7jC7GhsB5gEJ3kbPC/8Zq2E43ZTj9rhwkH5/StGfN9p4x69vOy1
4GxSLQukF95InGWIu0nmLX5512omgjVs8IRy60C3XOFwp1WnXIjsHF0GdFfGbNNQy7g4BH8gpirp
nH+kaN3aS0vqiJZl1pnGLgwvIIJgcgjcsKb4uDxSMUBNca0cEoq/ZT9RpkpQ2p0I3MbKPGqUFMiH
IfBHUhg4WPniFXHnHJ6xyu60lYudfPeChuVyuIt4AxyuJ+lC0sG8fFHvv4FQFMZIEnFXBgxYDycj
/jq8k1YHTcg+iK6hSMxRXrqPGwt0F4mtBIL6qcPoGpBgR0EuN1U0ASjZrBkgcMR/pWR6ugh1GRsW
zef9ujzHhxvXbNcJBJZvDW6ZtHSCs/aqcR9NgmQ7okFBPXhjc6A9fNX+Fi+iPRrWgajKKhDZpF3U
PCyNKyk/pQBuawRQzKD65lcgMSJjj6mM21W4vh79381ZJJhox/7y9xLTXPA7ZZV95rACnR7qDVs8
ymxx5Scur4yHlHd9/sWu2+nKoi/yRhhOk7RCcYmNyqBQ5jaz1k+6ATDTV82M7Z30d4FlENZLoSdS
i71opYmFE09aZ14ceGIxEbpMdmS5SMpK05GLdPSiUZIRn7v5aszDySXKDCpI+iKD9/29CNguPPCg
jwY8WEyCsD4/s2KMBwQiLUZk6mB6yhZSjqEd7PryTO3WnBajFZtiTIpRLmZ+K7OuI3/yX/B20KRg
F/8D0OIbXaYUiX65G81VlA8hmHiA9EbTmgLV9ohc0S1kXLXPDV1utHnEhsQgyslmy36CWuf2BcmR
uuyKuiuyuNNN+MPKMrTExQyoDNOPiHKnZ5rVLnh9bSnk+6HuTAYrgOJbVhsE+tVUqVhVFVgBzbH8
sAv6GUEoNPcpGA29gs9TI1oeJXi4u1FN/D5Zd7afmnL1ux6vFmzwRgl9Vhjuu7jTFoq8Z1Mu5F/U
FYeYNw0b76hRzxXwfVj7rcb9ibLkEUMMESLRfOieVzn07ABjhWVpXqZ4qI0kM1t48TydhOxQEuYB
GyZgVVv+FZV1BlYNS3xlXVmKenN8q9cImWqiGyCeoxrl5X/S6jpJq8Q0+aF5Zrr8WXDUeZzMgOmZ
ZvokIDigJ84TgzKmKUpfV/xtWRMvlYo9nCZDZPC1UHtZ2Nloc9yqx1gc77I/0e/QbHRf3KKiqwVR
qxdS6hWsha+ngZRUCodAE4wuN7+CweX2R+3SQyN8W74tcNipAXx0oJDyGaJzK+Pqe7Jn3m9rq6EC
w/EIWogSYKOXLfPfXyDUOPMw2eof6AN0eBhDtDt09SiMeGFPHdHeE813QcT1SmtQuEO0RMTd3gBL
GeN9QYt5wZbfBJGPzmJ1smQFqutIXAJBOZtZh6m2tOqWoXYbdZIkFs9SwGrhXFv9piVNM+Fm/92k
so/sysUh7JTiOF/YzLQAH9MBb4OFc0kCSQyFEc2apeM0eFaoxeM0yLbcwQRAX3aUlga6vZarUrvc
8MFxbq2eNgmKJuyuc2yJOg9HvxrevF429ZvdCT/H42Q94QPDSg4vM6e9f1dlB3EmIr0Wik+JelWX
mXRO0oIfABEOpa6pzabj8Pvl3wE/DlUr+4shGB+iQOdmiGD5TJYhEac7rv8VgghLY0eIUu/l5sNH
KHnb/FKOHm5AebMfh+CfsjYTnoRpVPr7/L5W25/GkyQmHJCoNxnklvav8o8bl4XO4dG8jrfR8hFI
GxrTq9/1/8xtcu8QDKtb3IqDfzmznCCFabze+svRxPiENyWxHf/U4RZpMAMC/Q3JpFu6aZ7jIdhg
ZFXQeQUxQVR+aJA080kO7jB1tPbCaS8NBcPi4XHT1zsXL9BQGroLStnx87/gTd1CmgzzaDgiujdr
Cfil7nAcnT2G2ZWqT1wDDAZIVL5Nz8ThJBDEh4eSTcjKyU+olD8mUaVkGULTf1ftUkhuLjsbt6A7
Vx3o8kY6HWiL3+C6ccwIR3Y5vxN6edbF9SEfVzm1FAogO5HUllAnFU3jBw01NgLW1E+JXQRL6oYY
1iyTZQWXhqdmAKlVBqaiLjEJBMllPPq7a0/wen1Esm5paRBkfnJlHW8I7E4ZBenfjH5IGuQ/G+B6
u/GYYh/aTxA/2s11Y3o4qXK3LnABBqOk6jgCly00oyJk8oba7uCKIXhXwsgsxozmpMfaQGj/zD0S
tHhy4pdmwyrspjCnPFUzZTKGDjj/te82D7pTZJ4vtFRzDIlsS52GN+6gphlF8IcCS+vvvIVVbNrF
yBHLVqDi77xXoMH3L1MED96S+S+QlK/ut+tIDlUzC6aomr4sZhRxvLsX/JIOztrUYw+95gjSc8wn
d+um9Czv2wCpHF3Ft6QjobCfdwe27TTbG+YeibIaGeeZs7ouc4x1Qe8216sVBdkJr1MoO20cE0UN
7Wy8biwst2aaf9k3I91qGQUge9ZGjoEcXqLiGE8mmXzg4SioERLIcSrVhayzqcJLnDMDto9nuSGO
U46rPkUNvMonyGPfT1uk3S7xuSjOWgTIvo4oid3ixmM1FKWSvewwtuA7GTdxWczOIVdtcu+7YCzl
JzyqJA3XMRPDdAEvyTB6GhUfUBXP/O/9T5fzESXmRwJbA/xuPtApZJvGvjvyx4Adm1Wmr44wwxog
Sp8+DsfPsQeQQgYY0+oPty0wRhsasMM/sUwQL156JYvD+wrdhylqnGN8Nw5W2BFHR6K5wYWhJZpx
vufMNsCpThJi6yGMVnTUMGv5Raj481Cp5hvXDgUv+T/FI0batsioCFS3Cb6u6YTcKaBFFSlDQzEf
yh84H8Nq1hIONHf12kvYxH4o1EoGRTaeDa0iIQOqBB3x+yzAz0MPQo0OlOY7hqGoNptoiEDl9nJz
iYmCIzUUkCGJTTLlK5TlEbgtJ4ip3lWOP/mN7eB5FPVqq+4PDtNPrjFpIsCC2+Mf8i0ntsQa0ozo
q6ZTI6f2egcked8YabjxG2NS6ZWYUgl6Cx7w+i4M/j17bcMNEbWPTJGGIlchSa3v1mueeVZdwolc
imt9FpkEZulB7dguSmzPuTAt7XW8KrnYujeqHxCIciniJ8bQEGb8SLZwOV7hg6i+YLv4jve9XJOs
ueGN/WsUrQfL41ehkFeCwHYUlxsSnmhyt0cwW2kpuMioj3DNqQrLDfAOzUtYGFgHPfa/E6SRjxAN
dXsApOK4lZEKRX6Q8L40xwiqcjuiuNdOHehbKwkvg1cL4n3UWSuNCdA9kT9h0UWklEQS1IxVImF+
AnPYHRpnMOWRmV9q23CYlxw6UbEIYYdypVW2JGweiNC5D9WEDMZNMRx5CiAWOxbVfmT9/jSmge1Q
GHZu7BHeAFq63IUCY4TurIQHpYjiOHOKH0U+0ZbPqkggTKq6HkiGFhcRn/k24Cln3PzzBT2r8j0E
uLrIvYAJH9GGgBy6Bi0IJxqTSi1hIe0muxZ12DpYc8MOCBjwirCOOCfhYJ8kZar4w0UODoJ1Fw6b
RSLH9O8LkxfqH3YSRHX4KLE9RvE27WrRKYGUsqS900Le/2AmVA7N2P6BxCTqWSGWAzXhygHT33Aj
gKuJ7rBm58VUdBQATDGHxaIG+VjfsUf75iPtPxy8/+5sAxHIyy0t6toddau1OpPm4Dv7Sfvtz4+y
AAQWlsvcX3IZJEQ+i9DDQmIWWxVGcHi/xVjcjdwVPp+Jhiouw175Wk5kgIYhYyKT6qo6fL0/GLHu
swgQAPCa2T3XMS2PN/xswGQbh0pBfd9qqtwWIjkG3YHb8POPhmkYt/g7+i4YNOF143xvum9CgL78
LqH2A0TrF7NvVAnGAGIwmJ9PX9pUglJCOmBymmMcFY7gnshInK17JCZ4hV+8u7ZcLSo/pEvJuR7m
XmvAz2NLqcTZDroIrX6eWYH8X5FRE36etcsXeSXdUKtleKB7QusDLELvLAUxIgrBIRmSTPhw3ge7
fGroCubj6Td2PwkNV7tSN2/0uM4S7aYAYybS8zRE7XKFjI3psTgPfLFe8xmJ6+GJLz6ZenArFVOU
rmyx2hIWOGKNdZdjYixt5UxCe0PbdSPULUSxKlor3HkdFbXp9rVj0FRtd/wLDGYS5TSaxxoXSH1T
WMjgILTUZ833tGdopBknLMorNNG5ZpV6l2VYLWUAA6XyBrWAW6hxcQFTA/elEKgtNzvXvxqRIJ+d
hKPBmLR5c2gK6yJX9qmDLeP/o3UdEdBle/BOCQe92w6y2Qnj4dGKvIeyxqiNKZ2agcSRV1rPgI0D
W83Gf9Lj9K4A5VX+itt6KUZCC1p4/bBmzdbg12ifGZs5M7qd+rJhXbQf/ugHyr5uHPw946Om0p2k
UwlQDf+Bdn1JZbUd90bolSdn020L5cojOCn1jGDTJuzxTvoKJJJt6rZrM8kBlRBZRptdiKFI6nAj
PFYlR6szc7zAz3Mzfc4/UXJyKJmoA2+CWZalw5gABjUZFHGcNrmmCJiLtZvb+i3qDMSF2rJ4NrK2
yTCJ2jiE/VBlWRuu2bcubH9lG6Ucivn6V19w2lOAok4hTnhXNW3jNoQ7+TRrMnoxtDwQT3G7N7wt
pRB6Mk2A9DX1LqluThUwnfWSzOxgtVnkdHcDl+ICrikLVGQk1YrWSdsxTgWacgtz2pjY9NmPocV4
aj9lKWGJ0j+woBC5ebQ5olCx87Us0J8F21oG0EbSnitqYwp6usT6oHE/LU3ZF5CQUflPjkiZvuqr
XNh/vbGrv5IxgQsUhj3lpU195xaqzXGlkG2bGiFRMs03i4Eqtho+PstwnqEwUe+D8N/MkdIpoPI6
2Rk0CQO3/0xb60aSTQbgR10riErYRFjfKwUe0+beAhqQVRDHpVYxdr2fnC6I0qUJIiRnQC7J5c3l
4ZlqDg1rSvsmwzLCB9AkJD2qTaJn5jSC59udiHRJ8pm5fhHaP3hOyr5UGlsj8NRFUpf9YsYdHQqc
BbVRvMAjCGnFl77cGa4haBt2N2eyjLo6YdDqQdZ9Ba9nvERVbykvM2lZmMc9zgLNHvnPzrp7ev45
nt4LeDX06CCRvt0JbvwUOqpPZW2s0ARgjbhmllQjMHYHYvZn+Hn6I4bubq7VgbM0L8KCndsBT4Jl
b6bpUjPlGlhgtAJVzvZWH8sGXizUiu8p5gQ+VPyOPhiPOmnK2tsvJLvwQAeggIFLfhYdydTKS5zv
SIFfjyeIaLt/D7snSIT2MyaRK18m1/8c+IAH5cjKIQ7gUVo/OzqqN9zyKZBr3Fryq7RtPoBEgxuK
Dh1M9+L5tqDJA9xS3XBe5Ws4vayrdofUnF4Ss5t7WZCdeAxyespY2eYnenkDtNeK1BL0UFV2zdvd
ToSre91eU6ds3M3Mkz2oLXBxtzYV+4UsXraGcNMtmXdT7cDGOacIrh2O50vYqqrlU+h/ljAr0lcC
mesPXem0OleS3W4BDy8TAYh10kHc/afhPyphCaG7E5efYcwdLBCJmPSGeoZcYDsuOQvKKcrqLzsN
/CLSUus1Zv0PtJ4D34zVJZXjWpy+c8xtViS+FRJwjrmJQ09PX68py3LATWf99dI9La8BMmJl3Cdp
qBL9YPF+0Cw31YuQ9rOuGDWo32LmU1/SrWCaevm1iQJH5N1R4u1tyC3sQb0GAvjS7lnxfT0AausV
u+hEEf3qiKYyKs1nBUS3kg8zB3VkInyozNebgNLqKYYoF7HKATLazTZsvLyyfphwpijgD3lxEyHN
xS0zCyeVdV+8MUbYIdZQk9EjB+QiLpwLPIkmxO/Y+qVPiNW0HmFdltW3DcSuBQ0DvinnVgquCdYE
yxoyqVOs9Fkcv67mQucUm1VFGfkT9clC758mhU7MB3fUPkxbzzkmcmLBBY5yfiWZyG6+rkav58dR
ldYGYOak0V7ldCevLZByz9+LUIrrKKho7JHzSDvFdEMeOziAqUzs/9tAnYY6jNRNZUw1rULPzwgV
k46SQb3DUBJU8+xUnawpfq69zBW37AhL8uSwBeVwOqcU8XH407rXBErY/ERjH8tFJzxoPBFpJwxL
t+Br83Z66LSMxZ7P4OPR+nIzpMvEslUnZWv9Me0if35BzLY32KX49LomWXDcENkeMOWiVgQrzc1T
nMSwYLk6YcWzBpjRg2pnqetAz5AMNtWOrQSoN2yJbbYL1BMGYfDWeidzamDbkNol+jS/9OjPhcI8
tcyzkV7iTDHSCa+srA9McX8DHQOs5OZz903gqHKoH8oxyhYAb+1kDBGR/JQ9irpbN6eCW3ObqYFS
X8JvKL/ysylaQEMhpe+5Zb2fJUT+ZnjxYbQfJlGR02LqwblfvGRx0OjHRhn6ZjXAj0KG0S96xatu
k5ebljKa3KhmWgsS7QYMzikXb8TW/DmdyeBdXaSbOdKh/noxd959ucFmL9UuWLQHDIPr3lZ4fjk3
g3tcld3KfxQhs3r3t8QWxL/9BJPPkFOkPmFKCpR4j0y2fhKbU6GRkCEm3c1xefd5lsrYStmyut/L
QEoFPtlHvD9gL3DE09o0wkCdzKRBpJmiA0UxXWcWLuzsqNTgSC+vN89+GYq5X1jCJ8SULeKgt0bQ
Q/CrBnVVfb+nKL4pdI5u7W07lItRGNJalLC/XHyZOGw/+nAGEsfYcQ7wj2BDzIwguIRpAX7520Fm
oT3HrIshm+jYxD7L7KDSCgfhCZirHMK40oBEg5LYzfGlD+d33cwdUxQJ9vq3IPjzYe9WzvOJ8uRH
wFCeVTm8TJnogiYBryNTbxSSs4i4bSzySYYj1sR20yMa+k5UtbMOpViKYvOIwSRgcOpsTtMITzLE
+AoX80x0E8iEVDvzwoqp9qUQQqQVa3AGS+ReyaVTkAvla3oEgI+pNRlqK/yfysvXsKvUTyfl/eEc
SfKB+BHbsuchOrqrcs/eU6UeUytYInSL/vtjWgsjLMac6uL70ie/WiBYKwwZLzYkIldnGNeR7Xbm
EYnCNIOrTzFFBHowS0hstYfMeOxaMiyZT7ifhVax8Kp8PXAgEpiEKXHaaNdK4yosGMBSj7eFXKsN
h5k9fVZ+u03nCMXlr6Uyiz6XRgMPoJgprCA/WyTvYSwRNE5ZuISxVvHbo9GhsEgptEMDTG5DRDQB
k/uolDKkEdMVxKESbvNAT7RVOP70fP8UgPvg75R+QH8MVSMn+P017b9gNxwqPZCv68kysdL475jG
B3kSPgijlBgW4divxgu4Q6J79SpgRs7Wr06KIcWjlOakJGxmzJvDt/nrqAAeu4UK8CYyAO+2yAVl
254AhD0MiRPI4bwoZUIoSvzN8tAJq4CJjyYHBSgCJOG6XZCzN0iZlhZWk1q+hmcyRpTVfbLcrBH/
fvV3FMRFtNOWnPMkpwrCZc6+0JkpOcisX8S4P9ZognkOhWkIkH9BdFTzTVHz1b02RJdECC7vWe4n
2Mfy6pNlvS3PyQeOfIyRzFPlwh+cuFnwNUh0WGFXIwgP3fBu+Zq+U1YVu9mia8FAFsgTq4YUzbd0
ov+7qLLahpLDSMDRTtszL/+hJWMWngTZxPj/EcKh8O0aVcuIMzXXNmru8sUs9SP+FStx6xYbq8ie
RjG2D7FfvEnkCfzrZkaxe1obnbu28EqMKNVlqiyPi06MDuMXNqz3Q0R1CPnLhqqqKaM3mCfYk86A
B8/tEY4p4mzU2vT3EgZtBDOOC8aXTdY4BF/ZAZtik/j8cpbnZzG4FpP49RSH14CiyW8lYox6QL+1
Hp0+IeiTu1V7HCEF4aq3TxCmyLq6EECYRX4RM9rZvzRYDduimQFfF14n4OL140VsiqQqBViVP2aD
t6HqnZyFteIfZZylf3sw9GejaFXz7OpKYqinWAeXtnXMlmQ6fTYkg8zzGyHtXBA7x3eudRqdLMWh
LELSR9lB++HcRyPYYRC76H3gjtaN9mNm5Onu+cZKvdJNgC3lknlAGzpxFC1jZqjzU7dy9re8kWL+
V4a7uV/u4C3w4Dx0n43vxZxtrMjjilm3TRV5Y49M+8q+WGfDgYC122PAc7z6/+Vqg60QxM/x4+5N
jwS5RrE6YaT7alE9MeY9vDmuUD01NmcSXxAwEQ5bVP4rDTHL4yRTc7DVLu/FVYUD3bo2l+tHKYFo
126GzbbSFirlEubP/aKpxf5KQaLiUsVslPE47i35qWi3ufkrvA304jmGHyJh+4aelhZvrMGmdZw5
aT1vIDb0Yu43K2MJwI5c9k8OLX7cHVFO52Ziw90nt0znw690uV/NdNtRbmTG1IPe4Bab9LvXkQre
HJlkvmm/bIj+QvZ+CIcvwk9/XTf50uqcE/d6R1nguOEvEG91+FHxML6EjMnmBjAthzuF/MztTwBD
L3D0E/o7Gg8lFUwCS8gIVB6V2eeBM4+Nl3qJ7Nk3WhWaGMaMCQuRvgh4qMgoxfaRgofF2TT5SdZF
l1HT7WPjJaYS+3TF+YK4ItcALo6mn1y2SA92aSRkajf+RbeGtQw1pZHggPoUSukasRveJDLohclY
RoqTBN3tPGL0abANP/nueAPQljollzHfa3gqtL/ILcHBYOJkGbMvcHXg/zO2Au7xGrGCUAHdwxoq
5iw7+AcBKHi8RSxsU+5ExhSWm0MU3ZuQz1LQXhtnKbWSn0J8xyFSVkMBq+MTZAFo2zot6SCxFfVI
0K28veRyPLRrWmz3WxXyTGPnx226FnPEIRjgH1CZW7A4rmgBex+Vku0TJGN5FeqRYVEuk8xQzJDf
tNcO+XBxASYGNes0pv5sJJZmO/CP2JdtGang0FhHzYxglJ+9C6g++1VUxD3ZLU6AoYLCHXzqJcjr
+Wvy0tCKNfjage+P/+NzQZevEtXbLCrVJ8HIOReoqgUr2TEmBurazAeqFGisUGvn6KxB3POSkJ+P
saX8X1KADy30nsSN3hKBlJIPD63j2yaxljBkw+EPcdgo2U+8DXHH/u4THiUzIg02lovpegoMdhOC
WcxvImDn/sbjLwuH+xn7zk15mCMKQpfrbq86sO6oX9wXGVbm1LPzJ+rIRNkxDbw5DcdTkL66Sf8T
AAJnyY4NsyQ5I7s0Wosp0ij9CylesuvAanOt8xcOrfbBok5q1wp50gD29eUaalX4wyESN1X+FCb0
Cjlj++PE+GJg4wmiBKnq7rY7VRmjRpJapjlwlHqAYfcIIxviXkcGkofAyFuFwdggHsCOL2zfYbxG
148u1EseNZ9mzAqFYEzbAfEwZt6Vr+Kx22TsfKfmzZhwlk+ngeFLC1TPHrnlpCGkewWkt2T0Rmvm
YWABrSh5oLtbWT5XripXANIv5Wvd8bZINsyzsVxD4LHc9RaaUhctzpXrFnjQXZhUlfj22GB0MWPS
15qas3Bjpqru6mSwTa8gHKJCgq4EeMx8txgb0sOxgvvFallVIWIqe8dYImXYCi2VFigpHaT+L//I
lFK5H3/LU6MYWWlfVpbuIxGcJlX7jop4CpahtqkHmhetVu27E+3wvttlNGnVJlC4UwxjBUjx6GuZ
f2S1pCNyl+klqiOrofwR+M1hNqnOrZ69s/B5RqAOez92yzRc9vnnO4iUcxQdQGmbKEMYI6bNDJQ+
7xxcgRbqngb+sn0F+ccOnI66NlJfQ6BX2zKKNT2CzwfyF3UUndRc7xtSAKwrO2Q214B5i46hti7s
wruo00L3yENXnByfWAsAhU5LeokBgkho9b6EnaSOH7fMTB+CBFxDXhGTMgR0FY7dsqdbpV7S2b4Y
sHm2joC0e8PTOpV0LCyaOnGb8Z9JK2f1JxYvhW4i+1ZQxYWdtc/KP+I0LrgG9sOdHU+qmlLsyIHH
hbsvJRfjdNR562EMp5UDRdCvtP+Ktt9wHgGV4QMPPD/WrwBbWbj0VKjsgGpc6wuTXt75Ru3WE+PT
ZdsrVNfK0FtFOPwcAzTvP9AyJas7T3FdQIU4NSa7iamPVqMMPXRLyNnlfQ/flFNZbTmO3w0I+7wv
uAOUiX9nD5ieklW19EirskhQbtfzlSp6RII+OTLCbGnh4UeDIGoyiRDM6YhXBUdTxjV9mC1694or
YfYBFdaFVGTlhhas2Z6aE93eoy1RSMV25PtubU/nwIcj/pEgJ45QVRQRV6+iDb4OTROxwWQIE5Jq
lT1sX6mxz2CvBxE+U6b7ce7DoZHLs1rslGTM+0RpiyQhTkaREiQ3DEP+IiF3YWm7k9QlIo8GIL0n
3FM+lKos1m4XqsvzdVkox3JyEmwDT2XVl0vtXhZH5xmPAsPQoyi03tuqjq6xr0Tryym4jaQc2ihV
jQFWsOrTgk17+IXNFsGLILLLirjV6GK0qQ10FiRLFu3Rp/JT+2cfAhX006CT0ba41v/NQ8LRuMC/
KYPH7DCiVGUWOnwIDTi6RromVrA+4Tx79QyZdamtCeYRxK6iLUIvWPMbIyUPQ/zDNj6JOFpdLnDM
UrN7OzfgZSpAFQhorGTIvMuik1yxR7cr7CGfdv65MT0zwzKce7eHaZXsSmDWJKu+0d0Gsd7mPsdV
sIrmJDIuqUAdtTeEUvQSaH5SOfF3QrwRoiZTAy6Z91Ih6KZUZ+F1UCwRDu9XVzyuSTux6IN56Tk4
c80+hZcsnKH4+D+O7HVK6om1R5oxnVdYm163oaQj0/YQe6dp+tQhRqAfBYdpJYh9ej2qpJEL8bLa
0F2qL4oIGCKtk8f2rJM6ZAfX/kw/Z+ri1aeQPn7JL027jy3n6tpWFs1zgrD0HdnQqzpA7F2vaZh4
MlHJ9d+p9o5K38QBSgjOovUVzdJRpx+pxrj+HMrLh38deVhJl50rcNFXTk6/AcAM2dxUAUWIj5va
GOVhPp9lj1qEmnyLnLWOn+++Z5oJwpw9NhdnqG+fBzZOycCax1OTbGdMv5vweptgq8HMFYLWjXEP
zs30o294M0Qk0GlW5Y4HyMSgkCKax8XhG3HeniQZd19GmBrF35c/4T46V8XXGlGGntJ5bkb/gRRr
pVC7qX9PfVKHZgwnNICiFbwnP9doJnYPW3jKDmCkUkyW7aGH/upVlmch0gXaSc8Us2L7zf0syvKR
8hwGuHOEr/bRmDmcXAmuk7qXaLxTKtiT3IY0wIczMOw4Au46YABB2RFfZV5S5Zkx/oD9xgPQRuk/
Dnr2lCNumysjUZvg9A9rv96PeRLLbEFce8E4f5vPoVrO0iOJopxU9m3TOM67RtAByXLbZI937fic
+tJGVdlvjnRjbVTnCSuCeG3IdkaN2e7CfKc1m8NaA9S8SNPBKz2Sw8Mu4cLPGG79crSfgdCVrj93
3xN3WivTwUBCGHK6HoiM+cDvlJTzIG9LljtowXO9YP8ZRfjnvYOzkurJZUris+Ge8fSM9+qo7W+W
4cmhZTtMFr079hGIPRdNQFgwZauiAS9AmdZr/E/AVjJptmj9dfDtwNtqs/RVp3Ay13ILW5uAU+Oq
btyeN+CXcWKncAoui2OwoPVwgp3KIQlIZzp0D/c2YRB1a4JUE+hc1FY0c8GjVg55A2EGaS05g+AI
G9RcUd6EzzJKeOr1bY2kZWneQGO0NsfcAphmfXVU4yH93w4iYHqtDHzhQPpP/X2Yahdn/UICxKG6
AUIeo/yQuUwNH9wNakN3t/jFrTFi1kfTJOOy8Z8PX7lD4WdFqaJAOVaSpVPX0DtTpmmwykaK04Y3
nUAcgOLKqhE6cJIqFq7krSldKbeQnESwKMKWDjsOZjuKKvXYDJ2bkGHcAUqGGJMA384aNy74617/
2SEBNNWaACMscXYAa10/UDJHC6u0vT8HFqeoTowBkdo6uQqJ2eQPKCwrWwfSxUdDTD9dwOCiNk/y
dh353cdV2UfuoW4T8O7e3tfhmZFi+IThWNlj8Yrnp2U1rqpqpO81uj2JOQXBdTm8N5IquCx9+wYn
Af8PUxFJrr5gzMM+OlOj6WUPj7ig2WvVauksfMm4ZVt9DM85Xmvnscj5z2NIRuzqj3Kx7yPXyDLT
pWM6WP4/jEbk3QyYYygL9ikkF2mVVWoALUWrUN0pIM8QfNgCoWFoqxX3xheKt/rVygCM9NK5bZmT
UNUmGirYJWam8CVXYE6FQ4mxBH2B86/WLZh3b6x/Xmx1xabgc/pc2/GB8m9kkZ3KmZ/ZLhDHnu1w
GYP4f73Ht27FRNlCY+9llY7UlQcasM82mI+gbq2NEy3G/J80KsYNcSw5b0eEZVGqSoqpo01FODqx
OioqiLiB9y8Ccr/wIoGYYY8llP2LEHoJldnZ3shE9vsdUpwsnappZADqXrZ0+Z2lfIDkgcHB2OZ5
2wvyqcy57rSzQhWaoY7mDDKHCKzkxMgXohHFMEneP6A88wIOsNlVuZhOaPdm8n+h+jlfylgzZj7X
ODzgLc/etsCUeAgIl11p6NhhCE+ev86FfP19HCjXx0Z/WTdU2EKLINYwvVC88c/kXGu8zX+A3faU
xnt6XER9nU1DAosOgmXT3AFgPRKie4IKkc6k2LsxivALtRRq81sfNQiB4Npb0DKT4F+61LbQh156
gunPgJolh5L7ajtRkcogVcrzbbPUx14jdJdLcJw/gOlGPtbVzUpA1Ipp/MmOACzl+hPOnaZc+B/v
uN2u/WgFrGVhhRr2FiM1/UIqaw46TjMfdcQ0skq/NTYh3buW+TbuglYXqJ0l7cn/BlrkGNShN7Em
UHEMnE8TfudDp0nhAZ+z7KK2TcNJSNbbOCHQw8Z290IXk4YemPzVjz2Sx9GjUmCd7V5unlmR4w5k
5QjIT8/8bR7vD4LojBPXSMB2suCUTFxg6D/blP4FeXS+6S+sXFNWMQyJRhKdpd5XIQiWEXpdrzVZ
Zuq/dNL4G4cXZNjGUZdsOI594ohYazf+qfiVqc21y9HE0Gt9ouc1E2QUKxkAWM4lM2YV040xwqoc
ESUFrM4f2Ec6sd+HGeRLYd5an/fVwZrb80H7R79IDBZmHOYJzESCdJq1hPgTqxlRLfCVIk7uCbCy
ivTr2Gn3AZcp5L/NT4tPuSdAmLXTosPw9laHnMjZhsGdkxaDQN3Pr8np2rDSvLxvIlBwbY2InV+K
wYKd3BGs1y7/xuiq/PoQdj55Kbh37pgwClmsBZpiOWwPrpfnM49jKjNjGxJHqAMwEa1gvql0TvRJ
4Eu6rOcO2kzg7cuXZ0rYOHHC1qfUqZpMUwEX+TiqJq/kM2z/TD9PAeLp9QdrWEZ7nBDc77MjHq9N
76c3gHzB7/Xhc1paRiNT4w2XAV2iAalHMe+aBY+4fUb9O29PG3+tlXkusiK3T1m0zSv1kHIS7TbO
9TIYKtGS5mIdxrF4drMWaHGFWwDZajDVpGI2Jtwgp2x8x80B80nPbgUTZ7fg/KP7s4w2RNgojOy/
CuIMkSvFYqPz4F6EDQta2FABF2Bmn2Bbrol2M3b+qImmWI7qV6Pg3G6FEdwE1sDu7OFjYeMY9C9+
krrm6L4W7zgrCM+15HaXLd7mzQ+5tulOj0/VyekjvLEX/JUsJXu7zxZGqaPmRi2f/zbK/Fk+1ct6
0PzPDnLtTmDnYGX5drcD4K9WIIzM11MLCkTlGtE74hiqGQLFXHWrpx6flzlof3xt6OnlN+SS1Mb1
F7y7UmJVKgVFV9pCAiKoTXEJaZczsl7J5NJ9ZAPG98bmSkrfsyMNh6G1CD50GT5rhgAGKlYy1lmI
w5lt0T7MKCZ2t0oqbrel5gMAp1pdJq/E577358kNJc4X2ZJW6TaeoY81EgsPP1aryKdD0fUwp2Eo
V2NXE+hov2CLfVtg7ERGpNKD9rhneK+u3OtOf2L3SPipYTmrZuuv7j01kYTvwETqn/GI7fMRQTDS
zeWC0C415U9n+Mx4sNl1uEIqqbyenmx12yC4jvWrZBYhpTpLCig5uyoxJjl+0U3B/Wtu53c+9s5y
pp36Ds7U9yOt71UU4U7ZuWoOwUkk+j2fYfRO0vp7AYchoGzDhi3VvM/j13nR6Li30JeAlFeIPodl
X743u2sbgPA47hy3dp5uk6Eh+/ngcVfq2BzBi/K6LIoI5u0iA2lhVPLFu4dxQP4Enz9nUAA7ypJK
LXKcE74QOVsxvhti+j3PIY5JELE92N6A8kDADxWGypKTcXrZsZ5zuzyf/lVD29l1YPW0ILvuoAC8
8UOdmGsRs8KOGVNkKG4FLqhTCPY7zjJYaTyYXRxTleV6VItM72qzKvi/s7pjMr0zG1D239MYUgnv
+3dDnCvE6aAJlviGWoF8SXmIOCe6PPx2M/jnUEtHHqgU1DMkrlcz9viMrw2nUNaUVg0Xe/nnE8XS
8heuJq2OLHVk2yqvZ3T7QxslmtTAmxmYVjRnBXXWj0ExpOEwUYt7yjyfhptCZC3Z4QeoEcQsJ5cF
og196t/rLCb+1JK8dbYinBjtSafLKlLxflUYE3HX7UXFQTsiVMjMcVH2fOnfptwXMhqmRmnFgunc
Ifbf9Ali7K5uAOEOvvodCoRmoO0Y4vXDqIJOP8LqynmJyTXjtEacsXe9iwc+Swz1jFIz3xYlEWsn
0ZFVTo+xccA/p5YMA7r8gloj/w15zl2u0kt+8h6MQL5mMVOQ0jJNfS40C9aeMwtUtG6jY9Rpum+R
OO3zmAW+QtiiPKfHWgipu1BSVqcfXr5s0vvOBnJdJSXsuPHAfNxPMyLBdnIOaN2FUTm8yEIMD+Cm
BjkzljWy+18THiVH871ubXPwXFBiD7xaR5cfvEQ5bKPQto8fiPTb+nVHFCR3zRN6HYp57+lR5V+g
E+Q784uWminnG+q9i0D7rZbJZo4lfMNyxP9u6vEQAaaiZ3wQuyERZB17OJ9J8PiS2BPnebx8PN0d
GWn8IGSMUYV3w32bxXtu9TqP5lPAGKR25Fb7NDyNX5Ek0QlQS8SJdPPjNQVLZQlb+skQkAWAJOoR
Z9mk7LVMo7b0khv1GaBVamRhLHxgAKDwYitFG7iqBQsffydGRPWpKxi6irAFPYuoIceYrICGDCfZ
JhvWu9i2K6F+w6fWvdnCnWb2Zg6bOG6WJiG2AMCkskLjYx1yX+j5GFSzcSHDdsttJUESH0tze7v1
k9QHchaMirLt+VFLZuYUgIJG8Lv8zjgqDOl0tGIYpcK/Pr/SlvwfhOBULHOzuNVbUyw1lM6HBvkn
KWlRVLF6kSYwoxwfFIufmHCiWFj5Vs5QazBFIGFAYs8TbNvyQ1noixyM/SaLN1lthSPdI9NoG+0X
KVsrlJzNP/Rgge4y7H3U2YNyE2dAiJOT5STsxR4JWDA7eN51Tx3K1Jh1Sc+X6jndwYVsSFBkOCuu
5ElYyncmf108u2sDzbSYp8lSDGYHLZvosDVPp/pkGqEeo9vSsXENKawfgnnW1HbVl0mfAPqBk72X
sGIEUpVvGOA4mVUQAe8A1fmKJvuN+9Z2eSSGsOI8KcwHltlhjSGi4QM98xlbQkM8qJJZMS1wjF3M
tXfRmXyuvElLSoVD0gV5hk5GydYFGof6y3eVUbGkSliRV5tnAADUyRsL6iEV40kRGO8nSljCn56a
ovnLBzPfiX3N45qD+lDRVY0EnmwcMtky1mLHlA1w9wzbvFChR1QmUi8ZyIicV0gtmBmENtKfLr4G
1yfff152vjNqJjULD2DJbfb+9JU7yG43Nm607wJL9KiDcQ11IPkU+7eoSNw7kgIORpT7pyrojDy5
Vrly+g0PywzhqHo6YNf3Q1zYp4eDNJA31gHwji2dRN0EqUmQqum6pzkv4RSyaQ83pyEChO6SE7Xq
4XI7IYcvEVmP2RHyFRCtZv/0F6GP0BBnFt//5XFV+Ph9xtyZfFmBy9xmrXWcATV7GH74c+MbUovk
VZkRHd5WRsUw5pXXnE9BMK20j9yjLw0pg0Rh55zehc9DQOHiH5dXlVA2ImSGdbkf4oRJY2ioaBBL
4UXV6ofPfhmAcpmyRyodC6uMtGWCDie3V9cPWOcttQPCz0bC3DUlQLTKXaxRBs1QcqF/Z6ntdh1A
eIRzQiODx0tmmMJNnjkM5Uz/owPhDVSQM/3x8L5D8lK52M1tLK1Naz5e9qTsGBfOpf9Rtvvp0g7t
lhK4wCRek0P943s0mh6Ac7cIwniIVkygQMk8jRsivXPMBmQh9/ITwWQP9W+OwECJHbRTwJYxLWF3
HpnyisCRif5qYBNAn9H54PimkdmykPPv9PU317iX55XJ+ZFDR+XAW2uGDa/AlSjAuYwiHAWXy9jg
xBha5BLDcXavS/F86G5mrEFox5WGoUTkZ0yzyVykgcXNeQfACrp1YMH71E8tniULFmnT6XfbePL3
TMwEo+rNO6et6odgj8hfEwQMA7ma79C3k9iNZfRNjCbFACncSwtNtLt1tWJqL2KA1t5kt5isjP+U
FsS9SvDnL2NM+mNiO+wJ2DJunUZx/YcZ1HWd0giyz1fxOHvJlmH+58u41f+m+NK5txSK5QP0Imee
iEQXIqDAx4+p9YGuwagd0iuShKbFag/AuhhtaVkR2wAy0vgTfagqV+BMUaf3H9kSQTo/ndW7o4ZS
Y4ncqw8n/KXQLFxAXgQ0oVHFC1zevMSC61zusx7cvkOgg2GNdTSj4BlgbEa7lXepc8d6MhxOuXrA
MgvSFHEpViSTD1S3Atr2ppyzdkO1z6GLimaXNp4hsQd9jVm10zL+A9nKIVx76viixu8ZeZM+QBvB
CDLbD4gnRFxuTvKSkmnbMIvNSl81oeOCMi+z2tTHFCah0IE42w2h6ohbkWgzK2wCQkHRlvqPDxC0
rBSYz92j0OXyzC4NaUe70W8rrK6IZJpBOvsanOeZY7+U548xiz0N0HuMRq1P4/HfMLi03OrpOx+6
6+qtIfmJbbOH7uje+RJGBdmljZslUMnfwYiDZwhhqRND7xOMCTxta43D7w4jFTSRtbCKD25pWvuV
38ExcIU1vqaR/fjdmMgds4uMDb9zis5hPbZp1cqqs6AvG1fVWgPQDA6DYQnttYQsBMHOaU+6HL7Z
c9gWuENrTmYLIuJnDW1ORSq2fgyR9Nqs3yPeisTdfUpf3RrW0825wmxgXu0Nrc2azPaf/8SKSm4C
I8MgyFds2Y9QpE2n9e6EqXtpCcgo1KdIhGqIcJO9j8orHcO9RSrZM5xpRhHC8yPYwiXnznnW6Siz
DLnJbthQWNldmtwhD4PlP/egiufMBdUIHCNCg7mGJgNWaUArEPdtp2+Vtf5u6/krDm9UTUc79q+m
jcA2MPV56IcE2SJBItyac9BcTL42KxDWzrvxSJZqW9j46G7UNwzlkRkG3bSISjcDZabJQw9MZzk3
1v9Zyvl4WdHEUezJd8lP82dYe4P/Lrnd8lPS5+RhukPFEWOae39YZgmPOtWPBlcUTkPOFf33huNb
l7d7480RXVESH4+mudxicQxM97Fp+Ta3xfxtWTVDvrQ2iNo8qUxEVwtLIaYd8+eLSPq3jPSyNrsr
Gpw+5gfdo+xgiYEs02xek9cPGbWd+xooPo2rCYH+lIPMCo5xCRg3Jr/1IfxKNaTgWkC549Rgzj8F
0Yi3rK79wWB2cgeHkRBx/fqeRTSUnBnRTmmdw1XOU2SmGgSBNf3twVDzNin5rvAqBmJoklKHnyS8
A7uu18t2lg1f3PYBgZ8gK+oaa2jRJjadtcIhVj5gU77aYMzYHUJek9EUdPcW/qxmx9FqEZaaOxwo
etxeAiQ3crTdc8qjU7rLdvHIwsoTT0kF6+vlD6YRqhlaDfe/WvGGdmNQvZDnmYEzYeYQNQ21qFKY
TVu8yrTUJFLxOYOT7Duhk8Ohopdp7SAkQelDZEWtjO865LAC1ceN0tqQYn8f4Q/EW5KXxngv/FkM
PQbpHJ6w+L86Z3E4ccs2zB4UPtmRfpyNT2+KCUFTShWI07gj1yTvEZLNilP4BoEes+OWsab34HDU
J+GOR64J3/vwtKDsg/f6bfJ30ee1QmXASDM4VSlppjQKXNQWRqAz0fsHjsVvtSfPnmxgG9hcKNsi
cw3fwmQG+9PazcKKP/OYXRi/OAUwmk1j1YBgKB2IohY5iwgWwU8ZsrWTHJIR1GE451gpT0xp/Mnd
3FBb0yFpchEWtO99CVurE91hhrn/x71L24kc+9yDPYPjgPHT+n5l0HxuHI8xYiV42Hi5seEvf+LE
Uk65soJxYf79/T+h+VMnKpd70QZN9vYTiockZEBqZ0Ou6TDeXJifEb7d0PzsbdQO3c1RGUYHoKlP
65oBkmmX7xgYEio6Mc6E+nQ81WUmWHP4IsCZlWrmX5w5fJMCnZ7tf70jmUTee2XV+hHYo6foy8xw
gz2O0NGGU6A6FCb+1M6nmoDpFDLQXtnBbK4T3pSzuBBy0PxQYoQ7nJGBaFhHNNq6D/1FBetAtU4l
IUQVhUW0jCqxa1Xnrb5uCXGqSAiO5xFL0U9yw9SyDrwSGUmz5zrsRLJYph1uNuBYtvD6rqkHyj1S
OQ5vKn+dsx536dgSgrw3PJL2Api+PI6g4xoUcnYn/vYEbUBAXiHhUMkC7YmPc/Ij/K3YV2gl+F46
wlFp5unR8ihSb+NOIy06GuXmpA2EKY6L4dW2OvbpQg2WbtkElFuHF5MoLMLueoVipHmczwM+cEzR
Xh6thr+4pJbsDwooHKngykdjeOBTEuUHaGAkaZRT8ArSLekgW/R8ZhOTVlgTw+8TkF0dKcrdEqUX
Xt14M+Mt6/LaAfUZQD2JAEz8g40SHO87x4BXFg+AQXP6fJ6IcGgW5Ju8t76adfrCFSlcWMyBwpBR
QqfQcEF24ekWdDvEccqp/asp6dgUzYI7Wo420LP+51DmF9YjPOD95NeKeE22hUjwjagooEam77RB
gSf1hincec5mAEahiwEvcI1YMpcNboEbI/T3aDghrDCdo7uxIG/bd+hXdVwg6hWqc+VHD/eoKvht
zL8RtRUmLfrh2Mb2tAsLrdJg+xA6zkDphHbXK4l18tU7opevghWN4H6GNlPLTkg4yM5o4X1RMLBF
r6xsrS6nnWbTTRtwrIfZb9Xr0IO+0WXqSlBAeZ6DhiKrio+R+BslbWqDy8T95Qo8yqjt6uoKj42+
ngL0YNlpox9l36TBwA+wF/4JsrZNpWTfphRzmnJ2fHWcTRAp1oLKrE6VvDUjpCtqma87sXaYhQxW
4lpzMSC2dox9f4iFj3YyuOB8l6rtMmVT2WcJeW2zRDmziJmmn8za51cZdWtvi4KHxiBRVXsVjcLS
GUb6iy/aBZJyBQgohQq0+BUJnDjsLx0ie3+8du2ufbWbd9bdpManJxfj4aVeC+m2RTicwqVu2LQs
bgoGVC4xHfhA194tJNn2O/M8U0l4zCuWaUToJjFRuaTnVz/lZrV+eNQ4k5QHODAaRYudLB6DsO4C
z7uXhFH+skWRE6SGDtbIjsRRzunRwIZeEblNk4YezROovIYSBFwGdTEAIMU8kmIq2DXfdDU3RrDj
GPvNxfe2+OL0JAVU3gHbTHL/IB3OCIq9fTO6EnUx8LnjmppreV/XX/nIhaSs+1dp2OY4Uj1RVN3k
uPAMUy7hddgndrOkhUjPiOrRncfNZ6zGXaWNKsjWeoSIBXQpCqPitK39M7QzxpW5ELRk5+1/t1do
y9h0As/da/z9I2x87CvHMjZKJwMFUw0dGKKJWn4HRmHZC52LKBQR2ST1JNo5K39L8FWyBMez3ZHT
nzI14TNiqhr9wJ1tPPdON34FtWU4SGt5879Dq4SCB6S7vpu32i6C/AFfWa02UlSIwmjI0aSP80P2
3qhl6dh67I1haBNonMxqYclSc0Acd9mZaLwyMbvbWYWiBFf8WysZhCQ6d5tE9esYbom2uAf57pSe
yu7Go79vV3xzpYsiQrMxquME1f7h1kkB4W7GZwxbIH50zcUkYL/lyVHDcFd/ZXrTtIBsyVCHeOTH
nY91RSgVBPSQSR3ek5tbB/Zk9mVzwIy4TQeit/iFitOTrvyyDKPrx2msocvj/MAVcr+9ZXizKrCn
z2an0nWH1ScPiOLQEZUdfyx4rD2niSSUpCWZ0OvwP4YP2VfJKZCvM1yQSkg6waOsJGTIOUYG7ClX
TQp0eCXZYkIqk/r8ahs6QCXXZGz6hQMUkiPZcoX2VT7tWr07dESPG29SkV/d5NOdqgVGpRA+HOp0
cMuYXMZpcl/5Rfqkq+KGHp5A6osTrbXAhhPE8bNBOH9HPDAtY+KYa4K0U2pKXbS4/DxpzDcj7eDU
tNL0X/sabg7injvg2ge9Z1N7SW7t0jAZfEh2OdgNyGV8qLAe5u7WahmZRlUTCX2nLZeJuS9EL09z
6fVOwiklEb4xfeNZ5ik/QJP2fh6wdyW5CwzYnMHTi1MNTd0t8MiNdC7ZXxLgKUuFOLgyyo9NgyFo
PmtycEfJvmYUFr351S84PsJb61s/VZdow0zn5VnsDcuYKvDISmyJDmmhnIcqH7vT7oTL+ozjIESm
w68NKByRuBXPgx/47xp7UzpTsEAGgbAU6u58+MnuzwJB/fzOyn/w+CAVm0Cht9DE4eKUp0dhAjQb
X4qvy3xtSLTJWpO0GjDKs+pARCxv0Adwp0AgmHlOpz2kD3TPloahex1P3MkI86yhGYePd0NRj+TC
/YPUfsOC16OTTMAQMe+sEfTHTFVSngsmAFw0tJO4RR35C120ijmUFQx/riBmGaLcfAoFzIpiGOVd
BBTANWVto3fW5gOSoDyeSvAp1Ks+k3FchOBMA9kol1wLeh6H1rGh0GPFQ0KUrBwQXTLIN9hVpRkS
fHnlhveOyI++MejCBibrQGo0Ln4hju903u4TQih8p7dvAMhH2osUc0EBOXbH/bJDuwbNg+tmJx1d
8+idqxR9T73CT9VpsKaN+ngeqxo8LRygkO+fbJsKtYsXCl16YQoveiGdxYiwwSafG8XSvh/2+FZJ
12pLWHekks2RPzkgM6gUxWFYZXkJm/lVu3pbbir6TJ+jf6CsblcqaTANwMwAsQl3B29wArqWQfQm
ZoYfn0Ee6/nxZ8bXvNICnCmWCuOdVQp3k/qH6h6oVcko6Op+khwQniLGFpqdkaCXFkLsuWJlqp8B
LPNTeLX1mAVKroMb8GxRwp1LBe3PP7EvEqe0NVcYkXJHKEPfQKzTSArlteBx3z/UOHK8lV2v+xPB
hVzyG1WaoqOdCti4YZ03IHeoVWe6ZhoGygxmh8STBowLoycizwx8OxLfikbZvpm/0Yrr2THUVRBY
G0L3Q2C3AWKXLNqwml5cuj9WTJdyZfKdgAzmYTI7r6+ZIp1X6ROTBIdPoPqgel7+JrektbWHcWKW
HviuOsv0ODsnjaqoHABZesqpPT/U298jhwVXEnNHz/AahQF9ip2JYr9B9M+C2CRvA2HJg6dtnZcI
Qs+LpMppzQR2D77DU8BRJdVCnTcVXoBka7qaA45g6bIomlAC2RObYYe5wvtKwXcOgnty9IWfD42w
xbYw3+N0+l+SDJbZNjck7riC9w+HdeXUzFZhwlVJKR/kN9Tv///kVUBxK9QyCFsZdr/EacxHc/y1
S2Uc9dlVv1jsFgfv7Kdr8XoQRGcx4Dh/Oam48NrqBmI6brcKMCz84OgXvXxALtpd0Yrxo2yg/tCU
38tXcAqagMygt334K9L7fPzeCotzxO+qkTYnY6ONLFkN4razDRuzTpIthe2agTxbzaHCv22oXMxB
RaADBU6Mn+hcc4cb56qsnbVMSDGjHKXGh3NsP8R9OR8wpyFSk/n2VYuopCx40Pf+Blom5bDw9ImX
HIZiw7UBS/gcMkikGr+oJ+/vEKBfEKeAhmsomjtsrtnkaEArDPOez59H/vApiPe2ScsBRiKD/iJk
XRqdAX+W1tvh61U5Xz7O/Cp1tnG0aiao7BOpHtvasO+E3SQtGlV/oWCXCw3NQaFDPCiKcbH38VBQ
4wwf3xUL17tyK/a1V/1yaCBkaS1VK2pTlK372n/gppAyc9nBKslI8smbt0CJHEGOb9EMvbf40pTR
RsKdJj2phPmjDIr6hLLaR1Td1IC/iMhw5D5p61Rx/+ggs+Yv1u6Aa3vOZalDTFp7/CFOZlNpoOKp
nzrVN1XzXMiNLqZiw1ngTubtMUnebvREfX9YKLBzQvSB42uwmdnyEjIrrehwBm+XTtwmdoLzjGHj
JDKKWdx8ST6gUot4q8Nf50Y68MmE6DAgMk7jJbZn5AsAXRaOsvkEStAaxBqjEo4B5KgMkDa/OIJi
kA1OUcLD847tP15U3KTOOufowhSnsreAdBNn0GBThjb5f0xBqMms5poD9EN76ptilNw01Pe7IUxQ
b2bFJS9I6uWh9ot+WsVt8H0kG+YLdo3zk9gs5caGCdKPKm4oxNpsZudq1Sh19D82x4PGcpw78eQ0
l6Lw4nb3gkKV55SVNtmtbVbdTJRY7HrJnxX/9OgoCLmQwYIEMWD1U54PqofauVWrtnnTloe9DB7+
WGevLQJQcWd87UUdXDSMZJdJs7SL0cIytK+EFQOVrGS5DQELSCl0SACt8N6AMEfrtTvUu+zKah2h
WQU4O8c3wEz3IO20n1wkZ1m3XfKZersXfSyYb2vpwPVZPQdv5O3H0seMjR5U4JMz0zbZ+gKveBhf
FeiVaHUjUNXp9wbMsZ7T6FBydIfLtNMPKxtLUkRBY2Qe672M1MW1tYHYzCPXT2AlepXP/b2Gik9u
5MDoiMyEKBx8SypIdqvEX5Oa/T+vbTKr9BxyJKG7cywUtVihwNRO4/H/AedL77U/+JDnRjM9Aoi0
JKPnoARbaZQu3s5pYwh2dbbH+XELvk1Vvs6FllryMv2cecqY2g/NjVgn+030YTQcef7FzO4Tu7Sv
Z+e36eqmcKlniJP6gVjwjRdWF/gvqCmkoW0HSb5diToWkBtySt0pnjvISWspRy/3udjjgOLTaaNT
NC9suw9tjnntr11jJJZQ2YEXI76D0EopO25fvVUFGo2oygRDH8vra35YVsVCyiNsQ0lk7OIxeg3f
6kOMshjx3/I/odahs5kZvLN5gEI5m27Eq0najKyXr7PEcQgUTEn1rK6R1iOIkzGXzy7pgW1H3kqW
5CYfYdIKBd1Gma/ZzCdgjGtoixEIrlhNcTF0p5VLmviWahuLyNJNJE5TgpwXuO/vU/V4UzZz+YwH
YwYzy43te93EsWoDwZfSlh7O6uLe2nxCVnj/HSF/Mlc2tpomUImqbC9RKP7JruMVCSq022b5P5+l
z/GpSNc3bLJ3t82mRuqUjoh4+iLccsAmo3WXWKpiAtNM0Sj3DryBBv3Q/B0rqUu5ExbpjiEupACK
wr13xGcMaA6peQFMTaZgiuj35046d+aMXcsrbrHAdZJwqQKnDmas6KtcFfDD6DwYXELDtPGp7LSI
WIB+HdtJtTR3VNdqM8Zmhuiz3/jw30MWgLmKTixXawWNy5QU0PqpFbCR58pjbkud5gIL55MTGju/
6gkANwGeZ9WZrPa/hzdr2bLdeIugruTTIVNbhL/n06DJ2nNBCvODYlJPtPJGlL0Deu53W58xL6pY
Xd5TGB4BUTv1HHXh6HOH50/TLIWQ+Nglf4Hua1A36gqshlIJaAmfOU3DuQI/F5KaL24EpVsoaz7r
wJ1iLdSGjHEBo4Fu3lsX5reUsC0IDGm3kNlD/Sxwd1TLwaGXoelmRsgFPU+GoKrYiCoAy/HOBd7M
D53RWlGYLdy65r5biT3KcaTQy6kqZwMwOxuMU4ET5bT0AfCG2zGuZgvT7D67C3u3RXyEjVa+pkRU
xuNO9bjqKm6LAc33bgxuEK+pHCkgR2NlLu0H729ki134afIu48WezDQFqwLE+KTkMz4Jhoiacgen
hw2HpHD2CRpr6LPHfv+u9oIkIfjTUVQ2PZv6lZyf0YzEGFl51gy9mzjnCggBZunFMqs+ncj6C3fY
0Apu06JW+/t5HRKGf+PMzttt+2QojBe818wXPma0xn5+h+Dt4xw7dpmVGLNlukYyYpRztWwSbdqL
dCvnpkzFefFxsV8OS6CIHkZ4qU5Ku1z6gPMaKleib3gy0upub7ykJzYsOXSMPtsZHuhwMzatLSur
2NCtu9pZOMuseqws6Y8Vs0BVAA+14Ekf6SQwOhiwiAEEVuJWw8mevPtgi5wMKFPv79OQwg93HDO2
5ujEmBXYpAS0sSMCuAcbryMv+IyWvO/qNaBePuVBzXwF0Kj65A4xT3Wu//2QSG9K97JHaA5hGSkf
VL7hWl4EaidVLPvrozS4ndMyikvtzd9qk1G6FsDylJ0lk1dcMiOpt9ucmQyUU7pxTBq9tMUjadpu
qzTadfLWEJM6pU93wN1cBwLBEhHxReuG+pVdPgF6ymRm32riak9r2M9bjmCxe7AVL1XEuuILzKM3
He/SVIy1J7YhiYUeBNWhiT5L2B6vTJp1/MlmXkpkr/+jPtdnUIZlrrkEePWzR+IW4Z7h4pSZSdwD
iiVqsEe/xmh+O2ZMThLlp274gIWEfLqfqQ9Lb1C5FD2j5UPBEHb0a4qi0cVwEhCg/dEILxXqZ0HF
6EhgFPyXGZ3Z9gSKmTvpJiTKwYzssBThpEFNxGkL4XIC+pnbcFciuDr+PU1VHznk5JVx4dWSN9Ph
hvkop0ewqgqewLOEI188gd8JSNxcGjLXLwpkPwUMs5Om77OzENVrWrDKoa/YO15G5wGf8Mf9RF3S
4QCELyXjfi2ekd3+YGCU//CtThmMW5Nk7moru/2Em70G23gT2QkD5cHy+VqNCjUo1YcX1W3ybr03
HZfxxqOnP3q8fVoReq77BUjrQ6uJQFAHnHDZQ+xBwx29qw9O7YHchUCwjwdIb9FiGCXp9ESdwWFi
r60alpS+0GIikKBGzaaso9k0LsUgc4Beh7dELk0PiN5X0T56qp3RYoIMCNc12xz+1p5xAwgc9Ijd
ji1q+I9vr5uj3eemdlFA3sciGPWky9wN6EkUvE1UQdwE7dYAILzRfJ0nHMBfldwnr4B3gM7ZUSrm
gp1xVbe3L32+bKJREixDxZ5aEIRni7wsZOW34T06esREQ2JHeM69y8u4509KS7z/EsEogpm6bsOO
noHF8aUZLPeVkQYvi8w/ruT484U3TZ6UcCtbHjk30f+jUaigdvWTkbv93XZ+3Ye4dd2rQVQRdXyA
1a/+pUdWUQ32J6b47M5tZoAkFoZMis7R4E0yTu1eheXvu2CAzUwT6rmfzvo8cKmYXMNOHHwQzEl9
3M+q3YKTdM0mzTczmzHtmE0HFbPDpLxgSmqS8ihvFbeXUKffrZ6fI/EAEoPBCLcxOuQS/TlZn3zD
5E2a4kr5f48A9iL8Q23EyXb8Xm5H5yiCdQy+9wGQafXO4/XPCalrUGlgi2lvKUFqINo5RwH6Jl1c
byMdSj7Ey+cHycbaRW2n0h3Vji7K1iVx04u7LXq3+VkoTHgExeqkclk+COGYto47d7hNjAFaqZuc
J2QTCCIjNVmmbwETARy9UDHywh/A7R7LiYMq07D09NvauQ9mertK5oyDEqVuNMpcdNqZGe5Ebq2g
VtK2galgkdRyk+Jj9v0TNW99fir8TcZ3BgSAJDLmXfcOjFoS9eJvUwngWLVekmzbcNhZPXyTVo+0
pVFn0zs1lingsFzMvOJXJO4TBP5sH99Kgv/E8QnejKJIQ/6OK0OFQVLVqltF76l7Jyk3tG3iFPCx
H07qL4CWYiRzyagKQzejifW4sMEsfziuYpMUWwFDf5QOyna4nowQ52HcctPi9zOvOVF0Hm5oK4NP
Gxe850D8XWExKSpPPvVzHPMb7t8SgtBuhAkKopI1llst6g/HQz3FitL4jvJi8Q+XDHrgTBRfFxSd
5QBete9zvUO2U79JelLXFZ/0ccQ36u+LbECfQDm3OFBhXj+xro2Ah0ko/rQJXN8m3t7QxE5FqGaq
77FvkNDRr33THB0K0X9MM4TkCkPRmU0XBNx9MQgJS81cpywAULCXwlRgqsVka+j1gE95Gfuspst8
oskHlJ6lpM2o7XJOFU8VvEzmvDMH+PeA2V5TMosz4u3Cw4svvcfXIt8+eyoOy1g74UTWjkFtTbUf
U3fE4QiQae6N5doCmtq6LD2U+0uN0nP0XCQGHIM/ogv/TjyMx8U6SckL6vlLTK8MTIwGM20l4K5Z
nzDHNqI32yFE/QPX9NUrUMI2OGKn3REMM75UhFJv3ZNh0koXO+PzPoC/g2o4FsJNwB0T7Kot6lGE
9GgVUSrxPICJjTD4gtOTznSL/98mxNLP65ZivDxsPWXBu5ep8VQh1rOR6QuhdzEvrYh+DE82drJ1
kVzKvKU1jsdcxy+uAGKdUElqqdmWnUbGSnwdgJahlPrawh/HLdAEbQwV6XOhSdtLkN1yiPhm4ane
zo/ExUdoRMril9BoSLIaErT/okWVy0OwGVTledsYLjN8H9aBnnnh8DYnprPv0ReED5a/+dA/3OMo
HOQmBtg8UaRPsxk6ijxGx+PXwpYZJlMz0hShVB7IO75QIQUuaoTuO61HjJz4sQeABvqhqeOwrDgq
+nMiCnSzNPYTR7F5EzXYiV53MeQ9wBc26VU4d2k6p0/v5lrGB98Luyxfx5kt3q4yS4YRW7kJV0N2
RvlVKEIQ6Yf6690ytNpj4HQEreLiIE8tkwkAL+J8OganaV0NH9FKCaPyhRVAL/dlKAGGVdNi/MT2
GS5tRRez5qCOjz+mVsj9vZlvc1sY8OdEn+b1B9GhbByq6aYJleyikUDjD5b0FHAL/ogEIEyPtnn1
1VcGadYNiuIfqDyORv/f7zM/DgjZUu+osJXJPk5XOg2vrgcXl8sj4n9CtPK66EjY9WkRtZ+1tnEC
+UizE5yrf62cVE4TEK0wsrarLPc5UzZIDL+E834Cl1eulnNZLtS4r6LUFZI3Ne8Dtko3WnAMd9UQ
3ztBYmxYWxOY4Bc/qKhEJ+WE1KXcP9+dpha0NzJldM04wsL+LkV8jkT3OxL5NHf/VMPOfU9p2U9s
y5qtHK8uuqAGT6+3kVVLBklo7wCWvma1wviWpnWmkmtTZVQpLD6YQw+7PFGnSSqBUjnYMCRYb0c5
eLDcNFQt4g6F5cNNqecdoT/DK4LcZMWy1736NsZeNiax41rXMaoTR7VW/34hoDNnL607HDRZqMlv
dIZdgiH5wpQD+C70weLxt+1ybqoVpNybz4q5rfyMH8bCmgI8JsPeiNQD26lvTF++KlOnh+8CHfBT
3pG7E0cKqqSMfO3pA9m0xjkXLPgeqDMmaNWmqCHNimQ6cxMEvTWCq42fIFtoIPDp/xnwb0YJiuRA
6fG0Bz6YDZDlR+JOZFKDcEmhPrV4oW5GE3x3UKX5I3yZjsCHdDalaGkAda15mpyFfpfdk3fh8ue2
rs0IgchpZ55lwSyzjjnO6zYG4LefkPb8dG0ZHgiYmXKstB52JgrSth3obnjdwQua1YJKZIaltepM
qvnyLnjgfOaXrsIItIxHXkHDupm6V/69g7iDiAm9iTZfVs7eH2Hn5goerXIMfnJ/+Y4llbjl9BAP
3ez7Irrn84BgcB7lX4OfM9lPhPOLYRrs6Xu+4mBU8heVgrcKC1flfGV1skAgQNm2KK/XrEhkVok/
jKI/Ql/bvkZY8LA7yngypEVSUb1OV9vcEPx1ffDQ4yVSb/sOjBTaIJIKkOB2EecqSHpKxRpawbYm
fm1u0RV0a9aH4WXCpZ94a7tYJlYNlSTrVX1awwCKV0PHac0so/1IFNtiD87JX8e8y7C4t0BGAEpq
M1rp8ShaEQTmpBmCtOrLE1BxM+jTT5fi/KrSF2BB3hITPMv8e1YobAbwyjAxKKCjfPNgs+0ZpSH+
ZNxmeSaiJ8lnV1hFmBiXBd2ZUamcK2DM56SXHgPY/Dulka7ANfiIla3+r3o/J9Xfby1Tg+h1Z4Vy
bMBDx6tC3qFoYVHeUOLX5MBrAXEIdO5py0LXKQM9boBSrMDhRoeGDYIkjNZFcls+OR7Qs7O9RfPk
pRmvBs8b/hLtDTOr5h9BQwb4+GULsOrzzgUtbIzaoqQwjF2K87GqnSejwyI9CyFRjX2w37h3/5nj
CqUoTKnCjVaJlOMAvGxpeRfZlBjcgWRkCABj9Dkxi6o6qJPBujIc8/GJ54rtYhF+CRZ82M4p9MYI
Ovl14dvM8GqZ82umovolqpnWd2R77/YUVYXs3teELDESWxKg//Kaus55BkP3bjCTMgoFvhjFOG3S
iDjxF5Xcz31GW6LvkLNQfh8kRbZ34IFr84WTUOQPeopp4/leemZBIeKsG3FIQEpkFXtd78AYY6+k
UVr7DO3LBJqtGoq7ZoeetWuZsWwRwmdBFex1NQ53leXvbsFZnRGzttXQ0hY6b5UZRumHsEBhF+Qw
bxhT9hBYEojPi2tB6Oe/as8P6fciaK/Y+iY1xDBkeJ3sUH44Q1O+zeLXarzXow/wDZ06c/MK4xmm
1E0bgvcHfjNA9jpvlwWKImt4LbyXLe/iE3M4J9YNl0dtmT18nJG72Cp9KzfvXM7tk0b+WUfyeWMi
cA7X4mGIdzd8BOU7Zgyc7joLV+C3sljHP49vLK2LyPsIfnb+ty6FnySzGJzobv/4wyNL9eV1LZmi
gxxm/TOrX4DBJmCONEW9hOr4dPac3zLky706cfobzuRn/qyZ9wqRTgXwUX7Hk+uIinlF+S4QqqLa
HAvmj4RNXr01VPJymGrl6G6ib3WsKiBUGsyBMe0QHWJ8QY0w9qV79Pse5BPU6JTtCnUsstFHVLA9
thuOSk3msVoX3GygXfVptjRZ4P5XlIsb+OUXIcnVJnUXXLUm3yooJm3EDreXaBeyXwkf4vVzC1ml
94ufxjpEK4CMCpOSeVHuOPy8zYdxSSmj8LB3aoO2pTF3ldyktRy53V0CogFaxyYBFq2HpK8pnW55
eotfqF7k5IHAVjcJ7dGuYk8JqADGWdxLdHkttS6NuUjtnbwl+CJBAYVN0qj2ubGP15FClDX5L9ET
qCUCNtnox97Vb8yUC6DPA8LEF6vqfsh71eKNtC8jX9St9AS+uZnx2hx1oJ1t021Kthkl+P8FA1af
4FR3dP1Ez/4694tRcHT8jDNZciinXk3vB5q7K2KhndM/O6QQshnhRLEDGhGNhH05kSusoJIBjKZ/
zNHsy+lws/dA9GFaJ8b8jlYHi68MdEkAVXc8IxtKPnDU7DAqlGoKXbbjwHRQ/1uYis8gLDsCO29f
u0pIPlrr/KcxJyYdgUquyqw2q0DrizU4SUAQIUl3HdWRB+RKbgfxNsat3ef3b8rdWB4UQDZhPHJF
hsLQdk7elP1KO4vP1JEgVjHsV2IokxzQoAtaIRIfxo3DmzfDBi+PMJqvD7V/TDyUg9le1Jppo94m
x7VC9avvAMmKXTIxAz6JzADDCTq/7P0fSkXizkmvqGHWjCEj2FrwCFJ/bceSQ+cuIg47qk8qq7+f
oO5gV8/v5D8HTI5kqFPwK7Cb6WUTprCI/R4CPxKq6iYVJyNCofkmBGINC7myIcgiHUqoKlXusGt7
r/t7PSnyR7CxUHdlqK8U71ljTS3mJrNzNsq7MRTqiX7tF4CTju9eMbVtEfigg2C2cW9YRM3oxjU+
GwOxnVpDLNDhV0Uk7Vcet4Ec5MLqUdRMUV2ljhI+htvstTijL1k0kC/SLuO3lZkiGi/m45L8oq4h
TFO2F+tW8okX5db9xu6Mt63EPHO1tAAFFcddE3imJiPywwsLL5j6aiC1j7OOhdawAr+uzUEIQBys
B5xWJgJ44OhfME2VG9wSarCnkB5PSsd1o1TaoqCMRgbssqBc+sfXNEQAwlk22JsO9vAd61QJ5H9y
zn2wRp3GKE+ZBgDwQ6CAhuqVGTkuAu0vCS89bMzc/HdvrcXkWDnZUx5I60hnIVeY3u63kQ6E3UyP
TdAQ1UKYwjLKwnBjWO/ZSaxLoyYqx/qQ4aeYQ2NwQHqKjjOQzs0iX1bv+H8PYZpsFa6QOPOu/NK/
D49ptQnLRynMx58FXQZYHY1dsEgWo7YgfqHtBMsqvxacU8EqcuJ7f5UFgegn4fUwOK7/3TByFJp8
ZA+yqHDcmaghpFqS4QecDKUPBZwOgQpfWRR2RpyIDkBMGAnHrJ08AqRN/prRmh1qlhc/9bPTI7QR
f4YQHN6PjcshUhq8RnKrJv7BpXbvf7ByBrV0ph9PZtLBuKfzV29fvFKLov/Ohzk59XMSlRaryVKS
C2HhmG3q3bexutdEpFk+cXk9BFkca5LZ9h6OgqECuIlsGYJ7/bUZZE1A2VgcSgi+4eWCkyRaMtrN
LNHRcF0MrRHfqCUBLV+224TsE8CPWQlC6UvJ9hjPAXhIJg73yqMU5vRxVe4z9v4+QFP7u0lTlSGq
uECZj0PQ5avl67dp2wqdh+7BmXsNz4fEriU4CtwQ+bbYJMdknhyg2OR7HnA8A4h9FwnxmI87qi9o
wfqnlOFW/3+EByAm3EEju/1CDWarq1HbjTAWnjFCqCxI23SyaPaq79XPNRt5vpuTUPQG9TIZYnVn
0RLhhUSAWcXX9WKsJCXqzfWmbh/fvj1OtJ07VDFxUZ1JEayXMT+U/RlvhFmZzKrWSqOZE68I2qzv
zcrSs8gvfgF0JdzQTbpCYtztIlPz6R0sniqa1AlEulkUE92wnm4uYxQDM+MKkLneY4yGcSYQv745
QRUgVwVJkpvvYNLZfPuxhIb1yXyynGjbT37l9XCQkFj1Wc6x5u2EyfXRwkuoQzZwf4bOgzBv3FRo
qbBZF+l6gsXc6+1mS7gw3Fmd3T94yvQ8yYLNRxAAwOzx5kYhg4OezJ8DIb5EhAqSS0esy0hHe56S
NHt2R81yQZ3Q1IYhuBXT0vZd5l9lBsd1a4UDALjj8GEcRNUv9/fRCSzfUwGwkvqKskXjgnSxYc3u
51PFkESsS3/YLPWvfzy72kQWMJxDqp2SsOSbUxtCBK5vD3MDfBaHl6qvoQEI/4TlMyGM7bzaugq4
wBqZZ7AMtMqsU+NxJ3+9/twdfXLYoO9Mga/Oionh/kdVxw3h3DWpwkdxfJr6J921Vz1JhpnA0Msk
UMdx0oco7u5mNsYDQxQw4e1uZWR/Ak8mO5QFFWf0uUBAMwgQ9I11YKSJaSNRO/KR5aupXHl+uAms
pTVdAF1+YASQLJr72INTjm9PStNRKI42Mbl0rwk7g1CBTt56Mpr12PY7jW9gRomdemU0kngImLN9
uM5wbT+U++7tbGk+NMvv53NuQ2fPIqcQau0nh7XBg8Lq4MlmTFiAdPnE+/rkC8PCCv9OI2n2VHpB
8BW7jOsniVQ+RMSm96iW3J7zQAx/GsGvOE30ReGrQBzGjwmufwiq2jidNJ7DS3nTPUW1xvAEyD8K
bI/4vl0ihpCmtYE09bHQGKc36sUL4mGjkCaXvYQppYmuR82oqpUPR964wAW9u0cGe/l62ZandChf
VBXUvTrGia8uP3QVH8qOAqAZIoOBtJnBbA2xwErCTwQDBJQuYHyyfQYakCt1p2UKdxIKpn+GVZl/
P8B+JcGT2o3nTtiCGziTQlrgVqdveM5IgebDppqOS+Zv8wqbch3TCVRmvdPzLCv79d4TfYIPWvN7
1lQqG9qOWBxlzz21XN+nbVUBAubVdY6JKGlDehQ50O6cPqsfNfENFL7ME4XlpXTFInbeNX5x8exC
S4iCrFg+unT7RmdZyuhmESvdKZuPZlRoAp9iSvUjzYqFDtqeHHy+rWFDhTkcelCMCE1IS6uIARRF
D6S0TtoKAtlAKadaRbyAr9HqQHSJ60o9ERhzcoalUJWQfe5rDa6kxAPZ9bkCpB5WvEYDG0XGn133
fMUg4312vk9aMOOWXZldabEwtG2qzISfysLlz5E9I8gwkQ/TtiOdMEWAdGIkwWoLyqBvbPZdPPwu
iPBcOefu2co74UxC6NMSO8de9iHNJ+CnPlnGXjevHrComJIZMFqabgskp+O6+mnHs9kdUqRgDZCK
eojicwjDi1pKBBEYGBAbvpAIgMh6U3ytgDsuvXJEZ9nxkcp/T1rd9P6D3EPxghneI+knf4QAWPcV
rIYj77HBXWpl6SgBttu8y/4LpzO3XNXhaCYta6eCvthtjziMz7lMQg6rozcxX2qjW7ZFqpuPnMak
9/qGKsKEBM6/ldmrDU1Lifb7UC8YGmsi0O35vij0/NDHWCTCVxdjEcbwmXe1Jdxpw49Xml4b2xrT
9n/CCyj0enD+VfRNCz40HdTWkR28yQQv2xFpANPqE9s9ax1p+219OsYvLPTRD1Ihw87Cdcs4jEAz
a7yoGZBjAWAoF11EVBIquRRUiFDrDzrokuanIcjncc6jZ+tEcigqKwE+RysFOkm84Kz/GzLqfruC
TPUU4ycxo5I5iUfy4Pwc4yyEtyq8iPkHamcrRmoxVsNl8iytQfLf88GQWMbI7uh6SX8MuO1B6E4E
aaoIG9305Cpq4krA+pFGHHDqPHVMzW20Ltdt4Fh6i9vh8hgynX6mhHhNWgyZImdPIASxRHM4lj2M
O2y1mhiBK/67rM8pQQs8gQC07xsKmAXAo5+VvpxVfAdd7/8ae9omKok4WPJQGZToQtWWsxIDLE1a
o4HK4rcZae9D9UrXB6cuYLwEhjU0/9p8F82TkBsKu1UIuPk/9aoSWUSRvong5l5zAk4gNLeUcflF
KReGPUtNs74Xv5wq293Ix4M5dzJc7V1FxlcfSa6O12Gf3jIth3KQcH56a0dbhJkffOJAt9USdtB4
2If8BLbf6GTADg/UcxruSWyKmRpK8RqumWRt+s8pINUYrC8ByEn7caAJ17cgs7ZT1mOLToS7Jkwm
U08JDPT0+4cMXUeT+UNbMX4ZVuQ4Ki8aknB+RP55XCyJAhvkfxbA4dcbSB4gubHk9X8jUOGBkHA0
qLGneJbhcNhIXFpcQN2MD4VHq7ejYJZ6qHqqS/lhkPYjp4FyLRBfuXY23dpSyzIxB7TwnN+dP8Xd
OJKx4hz5Ogmt6gEhAHlS42GvbX+Wsk8GJz2d7V12eEa+b9Efe8h6xFGYmz4ewhu+hMY3/W6qH742
P+qAeuio93qhwTs5Sfhtiyb+XCr440Zofv7/KryPd4CKolgCyCislEQLEtDdsLXB+g/XE84XTq5B
xhSCuJsX2BlYiZ8dNkEKWBNEA4Xh6f+9+vAt3CpNr7jF+V2T8jiehWYczyBCgU1JcIVgEMa4XPDD
ULLDgFuQrtAWnAxWjCdnShRng/MRXa215T65UqQYvsYBm1IVmpIEEbOEmgaC8wpTr1Ai0bMMZgV/
VpkDXoDzSdPkfWVZUaRb0UpMF9IzEj4mum5zwtJjLBNVGPajKdJAtXiEuw9bb1IeSeyDiuwrpi2X
CDtlWq8Wkat3JZ/xUmF7zJb277a3H0lap5WvIWEFNSW5RRg/17GzZSZdcekErzR8TXO2+3Xxkfhv
hVUxSs9for+ajNpVdhIZzdEgeRboplval36vKGQ9dVsLmVT9Q8iFigNSApnD4Xcvh8kpBkkYNczY
q5pfRfXOO44pBQc9MVneu3eI5Lhvim7r83QYIO1J/+xIuTbm9w97JMOYumyEwN2crOJOTHqqOrU4
In14l3edY+sUhv6T4B6ASnMNvGkCbjagqMggu7VghnIqgiMi2G+WO1vrBDd3t5aE6ctRsKjBmWdz
GbuXUmdryoKwpwd3vhcbqWNjJk6r4lLBWjlx+lvJg1F97M0ujdtE5hpdn6uZv+GoaUX3AMUAyaiv
GbA6PottINM024CI8zbGJZV+0CBOiv1mdEJ3ChteCH1LZxBtNu7UA0QyEsHyIH9Z3N3UnXQUb/vU
FF2cYM4OipwKi/pBblKJluxZEE0IhPZ3xXpR/2LiLh3bE1oxgK+YZpF5C9yJQ323d2i2e6FNQ+HA
u8jncxGXBqC+xJvOmqrYwL6wyiRZPga/DWy5it6FqGetpKcVPY/HNaJjRb/vE5BFo4mY1TexTfWj
REtLtGnG1Y9D6fBZ+IHv3kH77MW6dX9ziexMH+ueMrkK4K1zwC1L0QhedZ8lBwdAL2QXuYmnAmjE
4btYTzpzVjCfB8fKsBNbUEnfv8J/JF0Kz7hsPx74B9h2+D3wb3OuTxTp636H85NYHCnqXHLrYrSR
8ToZbjEtD6FkyCAqIYCmgsd3PlauHMHXFnsPTCjUebg1wr1xWhJ0JRosPRjdL25Se20E9qA0hIqh
7F3/0HkEi5xy+9NfZMa7SIJD/Q0cH5bXE5pLFN3dfS/9tpnqnqgNrl5/6CZ5QNPvQO3+mXBbqYxd
x160WRoHGCdO542Lu1UC1nUowsjX4ZfM0AOHPeFpdxJjcp3Nk2oVT2FyZWX1XodVGdIXuau+T2PO
qUVEiC6XGld88HoxZHXVN1DZLRtO20xioopHHUxpohY+vn7TzTeOj3pxpUKszY2gKeJeZW8Q7mAs
U7KVOfEdMPVsQ5RZLXP79j01rnQXomiIgtIVqEQ/APRBJl6By9x6sjDrEb/M3ZnqOBdVYpnmvj1Y
idxGuJVLnzn9XB6vydOyvHivJTBL+n48PtiSDYzyHqZfEdRssz72Z1A9D7JCcuo6Ltan0TKMkHrQ
YmPQC8ywrfU6FESba+ldvhMC2QdrHumLAEcj5Y7QVIJaSHkqblWfGU4t4TZY+UGWUe8VkBMqWnmj
37i/UBibNu8Q6IaIIdQi4BqgfMT5dj3WaSseRIGcW7P+C657W5mnsoRBn1m2Y8cvkCwWJwyo7QpO
ALxk1p08mOlwT2MqkVh36Jbc8cZWjO5ofSl1AnLckQsenZrEhz8fBQrkvga+ZpcjiFvxxEyclTWf
MLNnzt3We5KHp/xQrluDQX1MV0ijjjKOy1zFaGfFoOqBb0IlyilsyTkBtJF/Q3utDLzgLAQcScoi
Rg7E3vmm0uMlFTGB437sNs/rifcVLI/sdrOiu8ArUlTP2tU7nuAr/JlvKF5j8WHQB7LlDEx9vCEw
sVgZIiOEH6SLWyf2kYmz3w9OIWW18KWnaY2pgmaQPgB08mlWTU38JB49Y/jmWhWpgH1OzasZ9eJW
NyHzVeWyLyZsJNJdszAp1gHqcWpiOYwJVOmnpuIfaI3fPEdv9/2N3nFbRoNtVv0U2BAjaPiI57KF
KClwQCLvV3PZhiSN7oPfymQz1m4SmAn/2wmn7JwGW7Gsh30ZY1Ft12o4DGbB05RcXXAeDO6EcXbp
wO7oFlmXqYGxcCIIK7U20XiYejGbI/WRp/BuLk5boG9zFgTrkCBwHKAfVrBAO/5JYgpUF8ymUIFO
2oTJPv9Y0V+JrWHetQLqlwv+R0dK4pn3NUZFiSlw1evx/u13PN0MTSM9O3vCD1HWT5Hq/CTch/zI
8mmHvT9Ip6qQoCPlTtp33evd1EhzKZx0Zb+5OXvBsS4SfwmaIBO/ZwjG8fbbuHpUSDXUmNblsKT/
F5vn+anK4TMYr+ja8L4XqvGZV0RJ7/rrxgbObMs0bkV2idhAhQYShJt9jlIdsM7OIolXV/ZRrSV2
J0aZGQYupPoCLnHlB+IqpGZKy+WwywZI/rxhKm6XMQusE1VvyxERj9AFwRFSYIiA4J+SGpISsrAR
UKJYb9qfjoeXi/03IcE9FTiFjeE8b62hXwesvtZhjRzjyDRhviir97/IcWx4SrW+Duann1GG6sH+
ogCUzq3fgLyLgCjXunkIyBmx4GRXsbHkPgAcZ60+Gd/rVc7+mNCuhDSulATJPtmFS9owparsGLai
onj4Re6Szm0fYspEv4amBOIGkOJyYOZcXog6b5eqLV9wRCd/yjEd5eBKVadXhJHa9D5FFmEP9gK1
EFAhE0+R9fDov139wBYZ9/0suJLYmRQEYBqGB5g6h97x4NLmvxhoACLF9ml2+Io3yOqw2TuvLwhg
erlJO4/+GV5NOey1KaDSRdh6N/G9waVe99eXhsNmPM4bzRmOhX5ds2lMvEXYhDuQheFColcbEUnj
/C4lB/O9umHL/5NOS4Co0fWEwjS4Qhi5DYw7M+oKUpDUaIEcMJzciTT1bgdZdl0pXKMlf5cI56/J
CWeEWInmPlYkWOmcMVmPtc72i9sZ1zTyKgxcOQCeyGhRLXYHAFpJufWbbg5Gcf2FVs0Wf8+w5ayy
xbo+k/CqAqwWBbeqrv0pIfeNxXARbKkj+C8W4Nt+5wafVW9UI8Xm9xMxJPMaf8sbYYQiH8NIO2Os
4emwMS5cd3DHC3NcVS/BdIWfXM5uukUPOP4EmN7uO8JrISegTIHt0n2B1Pm8nty/mLBB/FF9aCgC
molgGswRTQM1KX+/05posdNS60LfzZCVpoY7iCqgXXroLgU/Zl3vlxIuMT1uEtF7DP0ERqw2pRaF
Awtze0342wms8Rim1Vo6Slu3bkxq9YW0fPvwPx3qhF7IfJ/V9lmtMNcmCimsLlJaYvgnBAz+4Xvh
6wdomYrchq0pMdgspteFI9bpKSfNQcy7RWxXxQx3Gl7X4ikj7IAFnJFWOtoOJ9luKYn+/YXU6XBZ
DKVPYyXk1kyviXCmUxvSUD64UxojDrYsSB+LiDXFwtkEszxqCi5a8JpHLdX5YzwoOGtgEj9seWZv
VSNdOdQ6dEMnlc2BMbM3AEFTxBU0rVPfk5SHK6N2yq+VQXUjGk5TweCg4Ie2o0y/PUGtv1blsv39
61VOZqJJS81LoFgkZA27zsuAYVLaFQSShT/Ae8y66wxSL6CA2UmE6965+vDm3sKSpH8Q41+h3kFu
jNM77+sdhf29dDc6ANXaLQs1nJYeBUKFeonR4alDUhnf663e1EdCWrEYfrSUaDeXxwigFGQtn1xY
0IGFexgW30YNoOx3EGjo7nh3ZHMsei8SFpyNviTUnytZ0HPkVL9LtkDtVLOoH75BEOE4aFV+Tr/s
sibZn6bPOYXMewjqCQI8Hs1F6A6dwwEIx61NcIgAQPUlaiSkpHv4MvAeCUDWmTYAkYRqFrId5F3L
fVBW2N5y99OzQF9CuXhK9WSpQ+uPJ55i4TgqOvYyS3o4ee48Ubqfym+IpleqSV71tIgVGI43+0aE
BsE9gvBnNzXFd1sernajDrp6HLAmxzTcSPw46n+vNj6F+xTOxnX3uicK1dAt4svBydD9zccBvlO1
iZlpJo5jE4CUOXPN13Zce/KXfTMdSSP0WDySefCYvmsgOzDi9xEMA7TRIpZODHe60IiUNThoQGfk
zyw4WDd3yIIz7Hrz76y5MtIQfkF74VeA3Qmvf/Bta4cucz1vsn/A12/XVG+m/qsBJDJynYFYkqdE
s6bgQ8EbfVry2EY2UcI1gMFd56PwUo6sKNOGDChmYQbz3FVZEr+XD3gDnEEbYWpbSbKN92CLQ1p/
XP9a3EImzfPsbnvmWqTq2HX04mtAo7kFMiIZkkHgATGg9b2k+85B6Qd9YcbsfAONmg/GOmrHaO6a
ENQfieQyL4p1OHr8x8s4mQmt7vw5MJ+yQaR0Gl8S8DcwrlGAj7nBWPpbM9DAWBhOJAvfD9nAr/zh
0K5KeyTnAyB3Mq14Iga9P80AAn+SuzoDQGXynJ/14pCcxJLTZqCMniaqGJPPRea2ZvwuS/2z+llB
TBzXU7k0HYdo4nWuJ0YAkGrs3AMNqo0b++g5Gp8jjsGFWSJjoCMDC5CjZjCT9ESAoBJ2AZGhxn0j
YE+XepBWhUSJrDBf4TQ1ImGe+WMqUu+IBXW8JjwS7ZWOcqwEBQAmcvkwPA0+G7mC/NQhYoOYFv/c
8V9r+4lZGY3BB+FbN/zHp94Z191jxcWPl97H9I0w+wTifza/YNYaQADW1feFmw08ttFeGtwZ22tw
uXv6Iq5KJkI4+K0lBYdsCz824mFxaE/uPWyo767dLlvZLwu/WxEQAe2yw8VilYp3M/3OKSKmNFpD
qylG/G8yPeJI++U0NHqYKPw55KLaoza1v5iaoKS1fdcEFpZB88vSnro3cq2B0mCIwjYKgnfMgfeh
Zx1Wt+fckwyqvDnwzVut77RCvzqMuRh1VjgLSyCFHC43G3/g68pZD1qM4xrkI74zuOWs74/rhqG+
oiCNMtPxqC0ya20dJkdZB3K+pLEJWbL3p7XRb1SGihAqMfN76BxzFrO0FX1/+fNYA911xs0sRxkP
/WWdSOsUhUxh7dJLfdEQqVcD4HGpKC+2lJ2knTatcPySNqV0gIGFz92KlnogmCCiGiYT1rA7gROK
eb20+3Vs9r4JQuJGb5/GKNgN0FzNz9q1AI6Xq3Q9Ix24QvDocZybhM+M7cnsSaVRIXUI15FhcaSC
/lHGfl82NL3M0gRdfwQD+tg0/C3ND3TXQwWP9qF7KzP0nSHyGVyaEV7V2o5NOFgyvA/KBHRBW0mT
CZM40MfvXjfh+43Gy8JdJae3p0ctyt/FSp5kWX8IRz1nk0a0lNRM7OrCsffKqUCpnNDw02PCzfKh
Pw7u1N8dOV8ubKdC3gXXE9Rjb0RFfwKutRc7Tzhj36srp3taSSZ5Hq49mzfNU1p/m6PVeAfn8a7j
ctaAqDbl9rNCsohWk1nPBypo9r9f8sUFPlkJSapO4HSnk8HjrUSlIz6WWgdtLLOiWG9c2pCYM2h1
cd25EeVXMMlS0sCq6QvTQoqiyoFDSO0fmAzFbtYFFO7hBLQ4HXk1QY3SWmgqerOS/7Yu9U0Zqid5
xChR499j1aA7xdnvbQwo6uS8RwQc7vMDv/YP3GbQP7r8kGQoS8QbOB/pA4b6aBC34wawTMIyCdav
nNNfLlWiAqzxMSL1h8MGJTNgm1iRHBaOWJs+G0+hNnR+V6WoQZKJmRInQ/1yUsw2PAl6j20FPSGP
+DN8H5d0FWF/NvXPPkXS4aMiYaDv5QDPHPUcrcprvorQdoycO/yeMav4PdCHH9iPYMvdKxhm+snu
65hGJui53tqkLu08zu6j87tNJXukMFuIcPfxL+vAZNJx2i+i4J6lyyk3tmE1IsHC6LkrK9gohGyb
SljX13qQt4cqMsObi4dC9SATflO55shzpjwqPHhJUy8ZfLpRVulaHqOpiS9lIaaV3gAIq0h9QNlL
x3ykMUxZCcaQbUE2cYvo82LSGQW7tRP6Xap3TV/lQsghoe2t1HRlejmhF6CqVaPJ3emHscmImOrP
gvGx4SqEUM47mpqKkpeaf+gq/rqVNLgOYk/JRfKPsWSm7rWU9DAySdTIk1p7061NDEvfCoHYCm6X
XxEuF56HzxKPGbishbfvo63h6zW2JC68vvLM60gReM0ee3CrFWS+AILTEEbhBVKPEl36o3nANsMM
AQKqCiMp7Hsu6b/rxL/+s/uSidASGukA6tsGt22ZHTZdhtywhc9FQrOwbeQUmGHbIQowTK5+cgA6
u5nymGV5tadaugDazVkCG7oHPyYwsltMLFpbkdRfLj7WHBnufDoXguUp5JOHAs85Wh3QJ0Jowt7g
rbg46b4VgZofSE5J5XbzKa/btg0fnArrr1yBdzL46jmRByginS3Uj3Umal9oVYuyaSKoi1pHRwD8
vCRD8PCjWcxP0im20CJUUorryxod0yx+fGY/QEY1FY/viOhj/Vh6FTNh7j7eYgq8nv0x9JMKzgsW
6XBADUXtowjLbT/mrgTxnHvapuVjBKOEmVTP8JpUxoQ3B/8BPOpSBaOIJC9OGjpjwm0IXQvkGSXp
tynfEXP6Yqqdp5NtpclGNGyC0vZcMJKHbVXdpCxZU/VozsRnVxtjJUQGFfR4P6jheP5Cqc/Pb6Uz
5+l5srzqQPuKR6GcjVUCkE4XMtRcAaEW4RfKaCyXMuEVgZ9alloylTm8nwV1BWvG+VznD+T0grrM
1g36j+FF2UpQMKqEd6O36B9IL25SjFnVGm7Hb+E9SH/ovnPgRCp+wtCCgv8qpYOryV35Zziom0ch
ujEUs5hy3f9IgFd/evtJebWzB2VGwZqu8z4N9yAm2P2K6qA6s5qbUGUntuk3NFkUyrTxOcpbNrg4
JGGNtQPq9CA28AJHutCWw0rOhDxj0W7ViCpvZjq9zGvrdbNf9UQ1FvgrcIyztHTn+otTPAvTtqM5
U08FxTbe8q+YVPyAVQqcQ9+KrFAkha/RPO363HksrPSdnXojauPyN4VWhHj0xdr3SVmRfKLnVu62
rRfEl6FXmYQQKsupYFOQyU3hTBIHf6E7nXkRQdX0GFw8+CkGf8Gq/Su8SrrFbSwhRpPXzfz9ug6J
Zj/fgsBeZiCUuYjj9Ch1LWBGYDyNX49aYinqropRoL1OKD/hby17xnAKTuIWxbEj6YZZJfETfV+X
t5spiVONtLsphEtsah3qzK2MpXIMndyIPtKroiTkpDZZNQyUJBpMlqL8evAXakbJopknDF6DFqkg
71mgl3BzGN0DwqBbP+Ph+VCkILs5zGjAecyUjC3DGzzwtqGC1I/Dpqk8UFnUce993Nk3oSWgucJo
F/bhUFcFWuJWSIEiuRRclzB1r4qV0SgzlKtPSWjJ/nKsCTqGgDmxa1eKwLWvFLX/hx7XQCAn1hUI
fIJBmAW2k8qtBCsoqzZEyEMtH2Y/A/as+lOce6OOKQw+FUgPm9auaI0PAoD//75PC4GMzAWKb4Mg
RUHD+xLGky2aXiXrvYLl8GLlZTywq5T6M/DPoW27zlA9kNp0a868CY65lS7f+odlLzCEYKdHySrA
kJQzEtoF1Xw0pmwfRngOqy0X7M36PKSdZ7P4JrDZjVkPAbffkO42EKNAOdxoUjm7y4Q771JIcaJ5
8gPp1CZ4H7+KsfcQ8dSazLsm9HCdN2AVevYYNzFMovQxCKLzZf2AqiBJbB0z6NMHFnBXEFG4HohC
oncjQcO4Utp+WjRR/blnoIlAPFNHd6mbq8ulECl+azAEtaRdiaGQYvoiw7JdvWFBz3aoReLsJbMK
CrVLIZx9DM/VSbgeyGcCN+UkaFpzDH08UQyXxpl0mJ6JyP9gs9ker2qO5tBpjMBLMeRhJRpBqOec
qZEACv1DyuYSGFme4zDX3SENjgltR4CUx/rEZzJUj/e7EyncA43vZwjQ+o2BYE27MBkCib4ePJYs
7nIp/Ilc0YSLPghcg35SdlgIOKTNuKYAWSmuNUmyemd00hFo3s5NEHfL+TTFEe/4mPSa5mJ4rQNq
3Ik4sxVOFGbnx7XEKHlMXW55OGTVMg656vMxRh0YhTk9yQkbT2R92ynQ/XM7Q9O+8kFBQx1Yq+qH
W/cWlVssky9201L7/nyFMS3cIUHB4/11ZcXPcGPI6w6/4sqHREe3kR42e0z8PdE0gdVmQ60qQ4d3
FGoL4oi+59k3gELr7bco/1ziZPks+akR3ZBk6B9LKub4e/nH1+VEhu/7vwzh95JOSlYtpzF8ICYd
XQ1lE5y98uEvC41JWPimoyQZsrVTTWTm4rmgko/BG/M9Pmw/2Cg9c5GU5Wj7XxfdbyOtRsPj0mIG
BAnZRlKyMiwEZa24L+gDYhOk/Eiun7hk4E8rZjuvNH52N08EOIqi0CusSkg10Gvh46gnWi4XxyDT
6xI8J+Ebg5V0z1rAgJKJMFlE57mBadeFz/M3DlfCl2tVd3OooATbfjN4+gOQFl3fG3+h6MJUmiVV
iSDuLyteGN1II0/xP2kW9RQ9MuHgJtb/HqDXTo0Yehv6/T8iW7EbkTx2CV28nSImEljkbwRedwaE
jzIsfgXY5Pwoqf04YK+QWqfGtvU0x38jmZIC6YI0C04re/QwubIxwjwnK6ZNCpJzpBPuIZWrUjcj
vJ9mowZ8QX/hF3+Oeo6tDCZjWkSMGtUctaEWlA0lnifgX4jwEF/+5MldRYbf0KBmaB28ghCTyqLJ
ediULrAefwkItE/YbXaBM/FvFzv9KyOw2P12zXCmNhatyaMy1G3koVl2ShiiVFijmvwmYgX7EYo0
9IyaNkJLxyVqNHurLBOEi9qSKW5HwtUachJHzlmnyh6+hDMkNTsHsjfmxIvRtfvyu1yx9pgHEPR3
SmQgnJ3JY1mrSKFG06PDh87VshxtMzeHAW+dFGbkMj6fzjkpwKA2r8X3904gi7dxDQVi0iXrPuz9
5zMDiiDDJkmsHb5qLH+dBO4aHvi+eTXYyMfiB2BVexRS7VdfN9z28QFrWQp9QE2W9JtiHO8E7JfX
i1JDCzfWb8qS0I1GycLIT3VIzW4EMcc1hDQ8yrUrtC0952wQp3PRwSlKROPAlPBGeRaGfq91pB9l
g5HLxhIrGL35V4HoezRBu+KVnEmfesgdirRPblLShyALs1O9fpyQl6g3zg9MmsKpBtCDVuyYkS/D
EZ9HmMfmbuXFT1UrBmsYz/ueaQPzIW4XU4Sj4UQyhG9PL60ll8BCWWxa2ET8m9J8h4Bn+qBFOSTd
gXX7TwgFHJg2/6p4j8wd9frhbLVS8+NsSy2XxqtjKtK2xmKxp1Az/vX2ipxq7fVl+x7UUW9YwSzf
xflLsBV+WLOo0rw/ifwdO30ZDwWs9w9zYHnoxoDfHWBuBKpH9NXsyn9Pa4jpnCmWLFG3CG6HoAXT
oD9XKYglUxk29OovNzHQ+PPE6L57LP/5rJms2rkhs0lDjhZtosaUHkJ/iLGcB0EJg1wZmD/KBxAd
eZGkrZcwesnahYVJR1IeG9Rw5v8atspDInHMal2XAXNykiqJ4xMpLyrcqKxlxlvPGXPQ/dBCuwpx
hMtekSHA7YdZrndZ673lpBNnHFLo5DXvOALkA4IG0j/YuVq6hQiqo/1jUkGr1sR5qEaBJ7sjhdbJ
q5c8pRBFR3OUi3onOE7WW+SA/LNCynwPcus5Tcri04m3+nMPOwD9be5VA+QalLUYgS/y31CPC+tA
dxWZ96v05X/uSG+iR6b/QHIXqVJ/ylryzHxj8cnac7ipSxnBOoS9koRW9dl9KLn+OcnwFtMxlYSP
3smm/MZNWiRMAzDa3uZmSWyKT8PgWB2rjco/oRnRs4IAYvZly3hPuxXt/S8XJckWgbludJ59QEtS
ddMnmF+gVtpQn083HEEa9PqUnqm/rupQ3CyZujnx2DxbY0gULhmf0HWoqlnayZA2R/DQcvL5GyOq
fTUDiGKpUNzJzfp4AIf9had8WHZXrYYDWYQ/ojbSOK4L/3B+jB+L3jABIYZy/dC12PdaUupxzo/w
+12XyXGplMvP1egp7aVRKT8UOZkBfBWZHf96AVKmBlrxDiyIqtbhKFBnOm+d6/jLeqgaGrUIUpqo
HN3gTNrADFDsjqJ8LliUzIVNez6FFlPHB8Yv0QUlmfkdMVle1tNNMicJGGLqlf2a/NPToSZx80Bc
A7thOA7MUukftPNiS0iJZgMkPq8Xn1Su4kJf4EmnbNBG8mscWenX3vyktJ+vM0MMHi8Pl3ejJOxK
rM7ZyQ+RMkacCVFWyJzu/uXYlsPW3kTsSoKO/yH/il4nV80SBDo2vpcoZuu3szm9fWIByfFbFZEB
+t1PPS+Sp/1AQ001ET3ka/oPX0bYAX0YmXbz1HK/CjXASPiYvHRuyajBlXnOBUtkJRmaIgBCdQbN
u1k2IHYNmz+rqFmrBzpLYQeqb1EuFGh5XTyz3vttrU6n9NL7Dz7fWdm6jKBqlB8novgaJhm/QOqO
KPgxIKSA8xex3hsi09C0/TsNdijSn/OtJGQoulIUtuHftt7TRKYi/jTcwVORtYMTmR8ZwZRbFzP9
IYFS2gHB08AXtdEujhh3rgUjlx9EWaTelhCNM2uUbZ5xMpVruyiOQ9X7excbkMWgXQ4T/GTCGRK7
f8aIHz3QO85sPayV2g5JTccBtL8CLhGIf9OmcrRKn4iLX/aKC9Zy7z/qu3CNAKtzU2R2xYSQf8fL
HjPtNTzJmBd9JPQqfOWQ7wrh0RC5AHca15EfofIGfIMqftXJTXTgkfYbZBaIobF1lAHCubgBUwDW
NojlZwvd3hKBjXLHHHLpSJBBPcwhibUA9eQ2y5D8Qf1T5zg2cCcQ2TVKf/qYKTPUpgWxoYJakrPt
mRlM8cU3eXQ0JmfR0lwxg4wHxy/qHSbLsCpuHCXIuojRUtApReSswIuw5qSS/FN8tkhub0Ft4u/Z
aiLBkZubJblgH6jrhhYR3U3IeQ+qgJFeLydrK84chrRfxK1E0hww9MzOVXJPRb1m628j0zAUsT+s
QKs+pimDn1BhIJ1BfsdxXqItZOfmLiGSEpsBS2z0+Ph1M/3CDevWWuXt3WhSHPYgoKlz3kfS0+LB
6VgCiaOmbYgwKQ+10kEH64l1pmNWHadqrcfxFaWk019fG89kFjf1+IfX0IJvZ1gzjFDijyIMXa0a
/ztYrg7h/V+gGGqWL2Qgxz65K815HWXjzmr5iSr0Co2hHVH78iane7wzHsDr2NeaLEyJsiL6KVW7
oLFHggDly559Bvl2Pf7U6QYGfhjchQzlF+/qiVyDn/bv2jtGVEY0ecs2aE7Ku55xSRy8gG4Ml7GE
EVmiWwjfjNXoWOsBgLaDnHYN7cw7gXRMBdBkxJLyuCYGsL1tY/tXyDWTo36klwK2QJbPtNOZwNFp
5sOrQREXwHpnnwOVDm4vkAOpZuz1KWykyqJYK/lfnSvY019S/UZogjDB+n1GCTWaDqBmjKDB8bAI
U/wTE8054QW5pI2Ioot/LOvcFauKHFvOnWyX7RB2W106Rx2d2J2OcehgMa5mG0owrcuJfwBtWdPB
O/tILJP/63ear04CgIytf4hq7/GR5Rcj+7FNhaduBUPY3TGI/ZxK/CfB5I/BBR0zqvCf0ycT3mYD
310O9zxdGXZmrSpwiC3G2KalqqWQGv4BGoYgOChpsjq/z2jm7fHRwfqVyxV1aygq3a6jQaSBW7Do
7uQthvbJStNz7De13G320qa04C859sN2h6l9Od2RaZAlyb5XjRXKXxQWtPMVZj2zS8QvFHOLMax5
W84lWxbFw1KaonLf9iSb89igto7baFLRtOqSMGxWhCEzXigNjKubT/whp7k6NP4GrkSjHSXzOCTe
jvazuv2hQis8rVZfA+x4KDlpX+PQKhd8R4n6DeHjy2mJi9BSF+cRaTLZX4UmKtqAko5zvVmJA10w
IigkO0C9cpP7preE4zyJpFd5iuGXNZ4/NUnYcqbJbkPiD+oNMvmU0FI//xHQeqX3G9IBQAtEx1OJ
Bscj4JVZZoyOiGgWRKSiNhtCEDql4t+N6ROaqvmsOXAsJBZjRV7/KQt3ZTPRiuTALiAYx/wCUvu1
r7qcuKD/8Cy7x44p0rWpIiqUPVJ6D756CClul6Rd0si7KY9wjED5WUhwRP/TuLZkujFt4i/L8gyI
/Wmlj55m1flJh6UTfkGhfMOw+Lrg8r1K2YiEfX/MNFuAAfPyxOhuFxYoWl6XR9DYvQxVjCM9xGHJ
nuvOCoVQQ8bQD3DtWiAr/1oY3rtpFgReCCIjyF7bA4xLtRM/lTL7CZrGFR500yAie+EIQc3uIFDf
9c4Dy7nUAMPz4vuPoG1CSm2PF6Km1ICajz00ecjkaMqrFgyAo6J3B3cqWo7YEtZ49Swbp+6NyMjx
ijS2R533S6pfXRaBq0jKyNTbqUg/KAcVPcabXB9g9JLHLVplBtnVUFwUBs8u0G4wi5JVvI+UGi4w
vrxAQFQhzvjig9Xa5YR55ZGKe/iP0bhhJO7i8NQR4ZjocCboKzy+FKJjp3lNYOqgUj/Fp5KEVFrp
bhl1WMZER3B4WKwKgZ+GOx8oaB4ughUQlsrDiLVamEaKciTFdX9IqIuY+fkZ+lA3bUHgvGtpqKfW
DrDDMh5UEnqGVg/WieVDia3fxSIyNvqWDVVJBjw/XSi9bXb0y7fH6sIXh5VqahjcVwtoII5FGm1O
BPHT+am2s7IzdbcHceeP+v1xut2oVi1Z1sLHxh7PBS+bQg1zWwcfFU6fZw90ekWqnW4aePgip6pX
UAwbxdgXg193tStSeopS9rjc8Jcct8pBBISabMYZVQ/MAbjMmm6MWz2cxlGaDJE8k+ZeiUBCwZBl
hwA6aIxVgWD0eh/+A/Mr1MVstYWKpZETlx03aPT7OYQCPTxZ7PWzzPZ8iUmbyRi2srwP3A3y6pZh
xdxoVB1y1kTfJoqUsv/JpLujO6aIXddL126G0E0VqM9DGyZXAirQGai2nzb5qxSHUHQV1cIX4q26
k8P7Lq9KNavAmR4PHozEtr/mGQc3WiRjxGNWoFaN46A1P2XduLTFNiCqaISw25bRuL64s14Dd84c
LIekJPci0Ph0lBdidxSBmUU15WWgZ/hHp0ZYe1cjtUASICGO/UMUu1CeMhQSI+e8HERrWGffB/rt
iZqXihHbsB2TYxc13wr+GfP9UoxXI0FLmfyOhLxONRuU2Hqh2cpaIrTdoSZzJLGkB+WV7IqEfyZT
tfG5H9S2Ep/1uzAtJiFEbIAICaseVjoqlViRWcRYXwcyt85GZAQqk3qQgzzJIF4QjCrkUE+ifgfF
YOYJA8KQQDKZlvcK5QV5um+Hq2LOdGmARbY9TTrlEn5vdPm8Q29aPnrC4dDTviBs9sIlqS7t97Yw
lkQY3vDARuCJRUL2drzvMN07ceRnWm/UcsBV1pSUQA9zlKvOuvJ74M7bQ3YImMx/+PWKmnlUdy+H
cbDHGmLksGLY6uNntk2nDsHeXcBF3BBxQM/ULq3K4G4ZHAy/0PnUoRGQkXK6KBW1NaHJ2ekGwC68
ztFWZ+w+bF4KyDEdRXchsjRnv0z+f6kWuIlUfq9GKNn321jNKjiM3OIk7aPQGKhdKBvSH6Cc9DU7
2j/GURz1aoCyxaRoOp0M/43lUFoHvR1wp48f21zl8C19ytqV9GmMqm9rfxxQTodZ/DroAFYSVUOa
Mbq7ZqgAKZvtEJjr19z5ZrJJNtCb/sJtbkTN+PmO3nqgQApy7Ga/i31natC6PJhZ37dmrYQznQ1h
7CRA4WGz9H1HYbwcPK10MoROV8oRESkiE0GkeR7iRmHdID6m6GyIswGTWh2fzme/AH9QZB8GxECB
Q9Y2fCbNIYXCeOUHtrV0qCfX2tGZ2bdZ2G9g215KL34s+/z1m3u4N8OFmiQ4df4KLI2WQYsvlPmv
DszbgRBYW4dRdTwMpjoh2WpDZ1aZywVW1HZFP3TPd+9wOkW2rB/LdeirgROCDk8G46wzfyrxfuK8
5PwtjBGPEkbdyvWxponIHtc2SoYSLcnAkvRp+Xhz97VDEmXdA17yGIujvCHv6WUlOvtMZgeNUcpP
OkL8xQ22PzmmlNc1cGxNbLHKTy/I8ERrCM18HO+NdFA913iuI1ksQWzwPVkdX9c7cCtmXw85FSBH
2bzndO4K9Y4JUY4WbVRViCQ+t/v0bjnLSBCTfM556BQpYnkYVhMD4dEIKWJf+Efv2zPhS5a1m3tS
v1sX7yVNqYJuTAvBwocn1fQtqr6HB09xrR3vzKRVU046VU+3aXVFlarJ4IEROsSxmwRlg8VqRYZW
JEfPJSAghnphtSpzwTI/iTZIlR3cChExx5YETMxFD0hhKZtdCle0u1X0GTrN5y21iUJ7GfdBdbh+
CwDoVsnBEpOyCwng8Wl5/O9+Nc2W7XTaEerx+JR4UhCAht9jqxDLhOFZNVyb3H4CHvWmSWj9St2p
EgndAF5zffJn7GfiaoR0s5KCrQMnESGe9oSZQStq9k5iCrV4lqlBKd62IH8R+5/1PneQqdDw5X8D
xb+wbtKhWH2onpeVQbSOsfYpqkDm7m8IDLZgIKon8/ydF/G8L/I/zwDFKq0sXvbvgDMOXuPmt/VY
DuO38lJN+ZtZJfoLq3EadEigre2r1xwG77la1EMujqivDFys15ceWrDLQr5pU3TjemEzkY5+spCj
hnO6SOmD5poqnVuNXa/Y/OPxnqf4fv8eFPcAUbreD+q56V1Nt3CBoaqDWfhmsyvaSR/p97i0apvk
jz9X41PBdUixrLW/QuhUqCDKU9lCV92wmRUlVmwR03brXPNkiyURVTplYxVdcEL/66jmyNlWOslF
XG6Ml+IYx2xGN8ew0EMPyugN2nhy7nPzRXLj8eeIX46vw2zUf5DCyn3KN3vzM4sNd9NvdV1npRl1
+EXHuqodNvtz28h/yKc+hBY7nSLGgW19E7BAUwhv6mMRg5+oAHnX01L4WWkt5cbjAxv1Qpiy/vyK
1F5W3WF4/nYdiHEol4GhW58PtfBNnz2pyHm5yRnXLvxEET0AmAR+4hTQWOn/pPt/v/BHarZx/EaZ
PtWoCKeAtDnA7vzmSC1U7n0mNmacE9glT0RyFC43JRpQmDzpCB1Vo96v5AsjMVPGGMzx+KMrJrVq
PE0E2ckF7ZLV5/HEZ61Lwa9iKQBFyGL3rIStUAjHMdsKUBMVqSy1QzGDYVASxL20gNCnK47OLoLC
PYMyzKxq+h7huVG3ZtT0/2LYXRnHuw4FsX6EDfuTGLeDI0GsJKrAPiHGFSYuMvgMGNh9En8UR483
9KhJQuPQcm6xdWQLNzNBBxIcyxSA2GG2rEldYlsi7JI8HcKJp5rkUG6fBmnn2d1NxHuhoarLWp+t
pWmvZkOAjIAsdVDHh3E3fDvYwNL4Lzc1LEPmYaNnFr/Njp2pztm6NcMD17hloPoEV/0velQHZmqW
oex2yo8D+mae0Z95FXOp9F9fjVWs6w9BI9ZbZjKjmDN8QGYg1tLuDZ5h1JyURSWNgscVuh8EqDKF
qJLEHMxcDwrxZmAWRRKmJJ01r5cpl9yPDXADwYdDOE0mqeM0mm/slBDBYtwiu0/06v34TwGxOCF8
gcM2mYBZdU1vxQItdlMA4GVBVOH2FzdQaC4jWggoAdjduLpL86n761wHyqAIZcFI5L28y+FrXo2b
RYe3LfPPIdNt2GgsLRJN8SGHJKwlFs6BdqqtCTZlftwC3IRA4VjCIIlzcjlTsrhZdqKJNV84jybh
v27xFGmC0HqlhGpqJBS9FM8PIFPbBTpyYxOc0SbwoSwpiBgNeZbNlYMYK2KIhLsCDo/mAKRPXfca
iXzhQQ/pMSLRcTUW0auTpAq7xz1Hn6rg0ukLfArgjKPgtYVv3/EcviFc4VRP8gd7eNEGre2w2oIX
wyiDx/94Vkcm45xHD+hDS81PtOai0cPDxFch2npnlVsN+TWsoQ+dbaJ62km8Iskw6PryyPa1FJv7
+6eikZIMlCg0fLydTONtJPS1GZukgQJo5sK4GCj6h8JMbO9mvmuqYxZPxvj0V9zrVRn7ABJQ+2hA
2hggGCCPaQZ3G23XnETsBt5U8kzecLJZxFi2nJLhTQD3lypRBgWLMUzwJ7o7mRP9i+syZG+RCWdm
y8lfYAl8ntTXvnooq/bU3Icj8VJKmD8Bdzs/1S1hFMA92K9MSq4uMigP3yLIBvMHwrscEW2qKMqY
TktYL+UyZK7XTks2XQM4U6M9LGzj9Jow+pr03B5pl7RhJDnZ7xtuK8mBtJLIjp7Utp5zt4Xh6NGf
GzZ3ualc1uK611gd//Yb8AP7Kt/dRiY5NpdKfJlBRe5UF1RSr7MxjrcoYcHMooct7Xkz55bP6SBC
THbxMNZvaUYfTLjm+0PvtEosLDxXbEZB/BafOkN7o9iH9hc4xGuLV4flsCmQRnVwXwupSR0FRDUy
K1w0gWsdK1S0PNjG+FAO91B/oA4mORYoP4wKLGyNnxZBEfrZB1cOoqrf31FZh38C10AkSKXoberw
d93UQKYU7ribsXkTcdE4Mbc9+hTvazHFB56RN15M06VbF9sYkOvkuHrz1VCbWNE9yuupk27gBbSO
9tm0BbgNwF2lkkMXnPWbCEYSRuqaA2uj5SQswW3atT2zps7CoXMwsHoJtbXgvi24NIQaWF2Dr4Am
uGTwU/MReRCJrI9cNwZ9sX8WLeULk9RHampam7KimY77AwWb+gIUN8SBmsSZoUdOqbe7TNgtnBij
VI5izruHjMZ/9odoLzGYQJrqAgpSLMxOYZEwyOi1acTw8oBWh+mcdO8uXYcTXRqUMCNIF2g0PzkA
/eIgUM5haNqK2b7X4E/7Mo89qx1pjZNDwFXlfuRSnxzhlXaWwn6NCr/JGe0OwqWtYn72H52CxYVy
qjANF2xiUbv674rXpdQKcpRzRqar655mfKqoetv46FTxQi6dy1JqgwcZ7/J4scA+35u6+S0yBJZF
o73kHQSFe7CkSLtf3dyQTh1KQlr1vLI9kMc+dQLHyQHEpB/G1Z1Nk9yMk/JORTa5mRseSv2L2QEZ
PMqkae+pQSu2f0bGmu0S1JUpoyaLhbHvVeIox1hvunOL3q1fTpwLyrgQBCnuavnNDhzdt8TpfF3D
vdcxpBTuVEXXKdL1kN1+flcIqeN/no64DNL72MuF+c+DeY318XWlJc5n/ZetUNqR45L7FyaJY6nA
bjDT7dx6Te5zmTNnAfzzX60oqeQqu5XBnl39+QM7TPfUWdbPR0GWmqt6VLrQzfJ+7zBJ3wcrnjWq
nrxj4mNTgbFeBPX9QrF4SvvQ6OtbFLaK660JSCremCEQLXnWiQXpS2+p+d9GxzReKVVjzGvwBpLS
iOG95GyDQ+W/jMocY9ioOIh2udXmg+e6V/7bcZp0AL8hPoQhKhD558+esr25k2LQiLsDDAfgTXAK
AP2FsksQj7ZyrmlOD0+rJU1IcdquWNSUs+LjK2d+HMw+FH/3Fk8VLe1BEhFdbdchejwiGRPMAkPT
UfHVM3R7fAEjPDXpQAVzwIMW774Rdo0iKc4gcIuy9Z3cSh6SDTaBKyo6jIRkkmaYjGz7fB973b0V
6ILhiwzDsDbpm4khy4jtdLAz87Y5tFmP//B8fNT3puf6Gf2fqTTrSmWOysWLf1k78Pft/uWpzQ1s
5IaF7nXReR3Obf8Ce0XgKqZ0yCVZElDUKpN9MhLeP52xvwF4EWSrFWl6o5mkoKKNZcfO8Ozih2tW
EyLk8VjZJuDshwHjvXlWlS5xvdB3E0S2HJUtRmRBJYwQ6sK8CbD7YGXeLy4hfxvbMWMP0WTUBBjA
QYiBvQDLTF2dG5btEN8T+qFOuCvZxDbDAnJhWRXHqab21Ph7YtQbqxAratSJTGvR38mA37oHTEIc
C1wBiarWNAYhkaAloV5/YyhGlY5vlBVRPVtIRzq+eUZPy2yoQpNowmimpIe13VBG1uzp9PVEo2dd
az/3GkmIWtV9f5WiWM6ki3z7ixf2uM33f/iNn1n3vzAxUFJ8Tr9xh4wvfOibnI65/JHe/IFivopk
fHGiEOvCpHN+xY5tsC+SeBqvGmgyHNLEJDzIjUs8x3JnSXhbJ7LqFFK5SkESGqmGpe1Jq6bFykJt
mck4p1ouPKFduHCpYpQCY9gTUEGz/Hjuc4uD08qyclcWXzoTstQkIO2CmdnUxo6yaEWCMWK/b8MP
S9Lboyn8AHaqfghGg4S9UC5cLqXWpNnr5bGUoHhaPbqJEoYsdQGzd6wqpo+/axZVfQUG5s+Id6mm
h41SyT92VdoYHQTKa7tJWL+9W1deZ5Fw/F1sf30vRQ6SUDzJXHutgkANOyT6Y5FU4jm0jIwS2wJO
fpCyVuPedHDXdLIf8j2goz4p/rvzUJ5nbX3+L10lRDb2uqE2sL4m/avigiBgAwXwy8i8KoHQi2bp
wvEUg6ZxyfkVt6u4rJtM4pfZmRrEgc3H+XjmAowX3F1aFL1C4+ZbumKOCvmkR5ku3VQQGQ7vcwwj
vw4SbRLJcA3R9Xr7fsgTlNn+8azSEYY+fAIw4kbeLrFf072fb1n3faCPVxyWclMAEs1IFQLnbpoQ
EO4dP6X3PAZl6NFH2aAYUBHUzOL6Wy6QE4vcL4BXFFDfJscBmXQDJFJkTngkyhMv70fvv7Ce1vuo
6vY/rDw1/o1lXwuyErGugh5PgBxFfEF8MmA59l5cNM6LXyzOjPbb4SJXEazJVlNXH0MWglVdCSoG
JTb/R4BVKuAg41dMdDa+SIVNjdv9gsvVZ/c4SyWq3+BkyOZe5MXEjWsO3ogOyu6pAYIa5SArcK9w
oypqhZjfUu6rNTsWUbN7l8+3yiXtUgcUgrZALaxISj0kkai1Dmo/k9rLN9Iv+htt35CPBaBrHFrF
eHxfr1BPJlOc4DlCh/+YyOR3jqL6mI6nw4W0EMJ4CZIZ6HE8mnLIhC6G9eO7Q+K3ff0fY5aybep9
/wJorzrmCw4ryFDwIBWIfliBksp/2y5r3eLtMYQGTXrBb2AxJ8ZPSOcHMcG0najq8+OWHFNhgOeA
uvP+FpONNUWxJWeAogT0yzmDcBNsRWem5QtpneXPbYoMR9zFz+F5Ssn1cgMBCmuMPXyzN3M7uoPS
KoNuZ/oIlkoMHs9EC21Pp7MSNxZHgcxidi8y2fe8KazIbQJoFjycgxGEoOpyQolhrNm1tKP7PHCC
yjT1EHBMC5iDx5vWOpAURR409yE/bbLhcDgCkHy0VWR/WyAE+z2kHBdjF7Jbe+LDIKV8J2ZIdta5
dxLcOyo2Tq9s5AGzsnKOSFi0sOhvbirX2b7gJXT48Xfx+ZZjc/HbsisUT/TQFEqBlwGzcnsRpiNT
dD7ZuC2cW3f96S9vkKdcgFBQ8iNGwXq6cjQS2/TNpqwnA+Xu0ZMuUcEsMwdLorHIhiK8VTKlM4Az
ZAS1DxXWQBFsTHTqLAF66FqoGWAoizuXnmmJ+9Ori6w05V+xqrRBKqYoluD8iRIHprzOzBVTJTfD
6IGxcNXLW9yc9qK42jZAGKeieBJ1ZNo+eftkeM13Qtslz+TKoN8K9l3dRs5iuTsihq3kUr1N5/5L
FH+k12Ns0vfDLhuLyczvwP75vOZoYR6YyoJhw/2bnaI8c3s6sfCaOU17B3L0yY246avX5Ibv+ZNz
4+JtOvCxzfqQowPqHTkodDOpa8Esb6BM/mEIsZjlwFbnmoapNCswaP61PLv+kmpHDXNKCH5iO4G2
y/0GP6/DhnKyZjoJU6eTWF3FyGLeCXr3Y9xqZ27hdbSpgy7AvioCbsmQYozUyb9+GZjNU4M5RcVm
ASu6SSPdQ8GAGwXyQEiATLfb1jGteaU/5sDACSuIrqq0/p7EmLvU5Q54Cs3MtTOxMZmiGHH6d8iO
koxsydehMREDBJIH3cm2nfWtgV4ZTzjLPQ1f4RCk2fobpcW1uxVPl7gTE2dsMxf8QB2op8oA+KFs
TgZ+0O0ZZWWBO7oxoL+N7jUkaihsAUnYOEAJh1elb/5iwXu6QcMbrj6dwizp36e3kzydy3reRv8+
FXWz1aoSjaqBihxxRQwcTBF/bysLG9HM6M7T8jTUCMnevVDA0X7Rnvo6OAVpZTkRge/1H+vZMTnB
CHz8+sAc2rUejTSilJSFlCnz8o2ruS9f/6L7mgP8mKs12HfBTo+6otG+LyCOb08mzaIhmAIVPCY9
ylj/UZyPXfMEoOIg3Nn7wWAWVCtvFCrWcPNMoj4tSNJxNd8GWCWsG0eykzMtWlZ1cOvcQNyzvKuc
Ia+h4idKykNE4SzYH2/PhP9dBFmzDGzrotTF7ebZjeuoE27N0xguJInzM5JJsxqMIfgf9Jd7pgN9
KE0O9yQIb27LVo+oJ8I2R1KDiGUvr+oQanpaidvDPrdJuGETodJikpB469HycYCIdZq/GGFkJzSn
ttqcKjgLFGuGSO3HlhVTTc9u/D7x1guafe5b+wbt3Pm9BqQjXavfRiv+X280FOqru02rSW88UVBZ
Wjw6oqmxvxkMuB6nduWb7A6p3lTjDdvCj10tRln92tJdnNyCPE86Z9t6UdyX2DiMKXxG6LsWLmnB
V7QXUF8N1SdWxO+BMwsKQYL5Swgz0Q8EtjNe2+qzP3jdVpeS2wPcEKRRqBi3Nr5nq73LSVpknU/A
IShixcr7OLJV/JwydRGWQf/c8dylV49M0GUV0SzkpjJ6LXZIrePkWR3n6v88axoZepzdETdEKytG
irDWEtKj7zgZ4ts3hRucDh9JnnRCcDgHA3OveHsAERZ1o3iNBq65uygKgRyLN7Cetfy3IafSsKPj
+ZBqcrqREU1Il2KojcbbD2RjCXzlkUreNlTGLCGoBS4LG1u2VeZug2lklRBB01o2OWX6NBADs0xd
dbC1npq7o5GwWHJAqpl9E/yTZ8ZCJPvn1Tq82GJD++7qgVh0nTJILleMEZUSQOiqjSYT2bh5Xw5a
HSSxEuGuej36iwK+5q0hlSDxWR2M/Lyh4bYc2hOGA8vRbvBZIONBA8QanfbKY6cairoSntShUX7D
b4hEInEfuv+L9RepZ+28D5V7/Rcqqe08lhs7m+mrmjBCdvYba41rBBr1ERy8g7LPxjq17Z2rqE9m
tn5x17SUyzME9LCVcwVhkU/u3+KyEjAA2YwCFB/J3NTR2544qoJWmWYd447yPJpi5RhgUubWMdgU
3aUBgwwPeB6y0QWw1ajpHlv9FtAycVJ0vdXJdd36qf23dqAvzcfGwKCVY7Xyr/Mdkj6CsExkt3iD
4TuMPmyfTP+ipHiMA8qcRgK6z0ItPGSGizZ9pBUJuQ8R7TEyBPSGEvTi4hpaH+Fl+Dfhd89ZEIBZ
zTrLIRMww/pZVS4P349+vq63akvpqEk0a0L/GRyXJa65SdzorRNBAiv+g8bpBVYoFDizQnQsqxdd
F68I0WjzBo9fsGs2xRpjNDOfRkOTjeqHhkX1RfOOsQQ3VWO+dW2Y/xDySgNn8DYQHm/FanttjuGV
afij7QeMsDLCtG5RApoP7I9fHqZWnP4JtRscmJXVmm1yhpf7RTUlv9SnENZ3DVJRf2Vm2EaG+HmT
LCiQr8HzO7eCSy/I+ZpdHv+KXYQ64T0rkLhg9fgobRp1Vr8DfhX2U0duJbCr1cj7OKapsNp7Zsv/
/GT2NwY+nB2VjfZEmty4ZGIt4mPTVfYUwgl+JUhkLuL+QcSVON05psYccOalFrQAfvBxGTTjNjwU
jJIhawBX3BdOo4tqb1QoVsd+sUPWcWpE9zSElKrdw0eK8KeYY4YEIntUIGI4b37luj3tlXZxRqer
k8FoJFumzk6GwPQIewzBRVhM46SfP8/km+IT/XTnIURkZii0Is9KQ2NGL+TXhKeHWTKL624TiZuf
/atS/9jJ+hN6mBVNZQGsiemZXTjgq41i9bovun65MgCFvwKqUefk/x6XTbkdjmpvV5SnHmORy+mF
rOLULK6JyegrCy5yV9VXWqgk9t9j3MgWCjuFeifGc2gUBlIxM91MWdCQdaG8jj4Gya9t3eWNKW3D
lW+Cy/l67A01QKpHZnk2TNNkkajlXYU4E6/hwXKJW91gcxhlvA9kxK4eSNy0QdoBVrC1MIIEm8d/
IWCxFvm89LBnAlGkcEpLncunYQnxKl+Nud0u3NqnRZqA20iJYsHRdRuUG8/SJOGdCUc6tyvlGgLZ
V4WXBGsoeykCZnurdMIWgOQ9xTz8oH4ur7RVyjX5AFpvqArdISZPZHodavkYkWoGUfG2tomsvnP1
ntbCidiKiJD3Y2UyAHeaT3hTLo4ows8eSmJ2rL3Oqasnz+Bru65Q+N0EMTnIxGrHqwMOBHXj8hk1
O5Gf0P55P8/mXCR2YxsjjvH7wifz5fDRt0iQgWIQAtBAdbdcSxDYn8AKhEemlw2tudpR5bsFD4RZ
puOoifP1aOmuyE+W/eeHDnnO0RQa4M3rrKnbmQ6RPLo8euBwZmOePZ6YVTWmWK57Tg565MWT7s/1
//K4ey7DvcgFuuTFgDJrMmmB9l6nX90m5ICpeYN6K1mfS5yoLGOlPHhQ3l7d0gtrahCdIrf9I9Hm
w8PAbzLzrzEess1pj0Y4/ESFLfc6OK7kIQtaLsIS41UhsNnvAaZngu0f+VZbXYIPK415BexCdcGk
gJESJ2sWri9xstcuWXCkEczqEVt1VxBAhKNmo3nLYHkVQ1tbXTdrpWkoShawouFxg1X69oXV5dUz
ihQxkxNjAjlEBi8MNaRli2rFTYTvZ37OSTR2maWAmh+h1ukP1AThHUZf3Fl5vMXPfaE9Irns1cQ8
WWkQWuFCSFSnPIsgijov3O9WeC4y6FbICHn45ZNnhqMZ00ib+zSik5Rvhpa3X84aPBsR7z12cKV0
58rRPPQgGQePFV+e5McCk45IlTS8w4TQFXtY0AmTgZ3uHe/aVPaPhsPctCydj4UdLbSoIw7EoMTp
e8OZS3JrEtPwC4tSpYAEEwcc/7Ic+gdgZt0DRlSzIzwgRcInZ/3YlOSbPrJ07k0AQ8Gv8jWQ5n7Q
/uGbG/SgoQvUhEupFFt4M+hdP9EKzyEXF6R/oHYSQvymwi6hjLbVXQ21a+SmRGfxKmIBPwhRM4kM
WQktTIMAI889lvJNAfw4QYeZx7TmOnN5LY3OTbqOkPHdt5Vrc53RnP50WZQCuZZVv3s3muOq+9EZ
I/p7Fc3UAupgiFEDds8kXge6lNouf7DF2R8e//hyXA0RjwxGommzgzHznzQNUZuppTOZSLcap0Mg
J1199pdWbUEBxYZVN8jSlha0Km2dtccxv0ybOg2BGpjRYVUPB0YeSYiNSJbrpuBLE2u3l+Uunsss
f4E9l3Sd4sWxyYS1SdrZGAo8F4GEWrLainZQuU7hKK5N0wTDtoKpFbAXrAdMzzPSETPpXTpQxImD
/tEbF9cRYxMyJ1BHbgAJb9xoqbaceiLWLJYO43PCgNNaVxIlZP2ISp6rOLx6tAk2oarPr/FBdHYk
AhpytznrsIcUmv2D2rQ6TgPrQIl34FSr/zpqfBV6rLES8Ex6B/Em7fpxLY3BBSEoyunWKNoTsHKo
zs3mATf/XuNGDFk55WxA0DEJFGNlovgDKCDY7SQcwJAfOLyL58jjdeO3rOMYHo6hKmMplNvaMXfv
pRIQs/BfcsBjEy+uDjtWwvZrr7EpyekTxciE+qvjSH7tJ7bkFqULP1GKS8+ZB9Vs8nBFiVkrZI8e
VZYukKPfhgUCti7p0BOkQjBuhieOWsVcOaXxDfVc/0qeDDbRBiR2dyOXvLMWKomAH0DJ7I6q6Ich
r0iyi8/Yup6nGp+ww3meGa8hdYnxdA01KmrPEy3YJFcX9+s9XAdlKoDwlPI18BChYxNpNKdNCGFG
zDj5TaLYx5vgsxAKm4Go+PBpssK0IDNg4UNzDU/XndP5gC9vMsP54dbae/+mKlANdtUliRh05omg
lWNT2oNOzxPadaymWG133tHowHOV1uU6AuGADTRRmnqDxyRXCobe4hl19JnHiE/xWr4ZTted7Jre
BqWm0v+eIBs8f8VIqZQfELC1TTQ9qQVZvonbMv8HBEOkXpxAg/IyiuycvT6n5WJoHaM9/l7ZUOA3
VmKiUAvAarvF8kaG7kUbQkAvH+9vL0ismpva5xhR4K1N4+i80epl0hQwUdydCxH85M7kR/qFMXr6
0BqzHJlATqgFeSyH6DZRXWnuyorfNTIWjcI5DFMppAnGoC5R5DD5g6JtYj+LVnoZsQ/2AwSxo3dQ
GU9i3h3Jyqfv7/wAm+lU2hG3pFEZioOJ8JAhXzrN9wuV+lqrccQqPnH/aDdohzG2fL6n2ShkYjkB
Yv5bapDpXKuzca9kac5qyqlOQHGFk6oY1DSUM35vCC4iINpvl/Po1oE3kHC+5k7Xf90AChkEsNYZ
hCu0dJID8wZ114dgRFlTn8znVQ4WS1fWhP8MQjOv+fVEg+juYBqW+mUGzSm3y0bgZpuvMFbFiDeE
62cmeSeGmQzQQ7BBuGjB9i0182VcwLVwl3XDW9CcW1r17H+YYyY8WYa3bqaL7LOwC2BIjtLSuvzw
jsXGC3NIBUlY0s5H9lZA9+ZDDA4u5ACCRziAuZAL2EovhAKfLiUON67d2IfayUfDCigrZ/CwvD7z
yVtmBaUFs//wWrIQ/YFrnMH8eziepghhYXyp6ND7zYtlO8aphseyv5/wKpL5sKQr0TYAHJBy9p/u
2T8fql0824ankxe3iVBlOxKtTj8BxJekoQbGoJncXCUeTvEydZgH0WmzIbo3RCvtfsQles5WD4hL
rvNXZNSbKYFgI3Eti+h8pjNR4YKT5LXpKTsDiORcCSTOsmsX+AS1PZGtZOGAGWQV9kx/Q/7a9QDh
bP1s7B32mRlXBxt4l3HIRmc+5LmkfoIEPN5bIs6r37wCpv6KuT9gCQT9e6Z5P1qWEQRyWfZ2IrP4
RbZMYQWV1pu1yPIg4bLkI5wgUrujxs1sv6NZOgKvIwOLrxKH6Ydmlr+iCv6hXNvYZcnFHxjmrNxa
Tg4ek9UiV0j7F2JJeX1xjOgk5Fh4hOhr23BADiy3RH6ladB2t+6zJaZZZu2rqNkma5jU3ORqBVQ0
gfWq+BnZ98HKnx2iRKh3H7/lCyYzR4hwyS7N7WVh2AgHfaPv8pI8IFL3p2TbpyVeKAE+g+JbALqz
oXTpqcTsAMBnBah3HF/F7YTKvh3VxNQ5RPPyIYcNSCG94qNa0+L0UqjT9rcIdNCmpnS09jjL33ef
QjRCO7ZRuxf0q877pAcAOBb9n2/VcnfvC8UvvoZhE9yGJBj0khLkoKbejwg99cEIHXBD+NTPFm7d
S3jfjGyr4WG3saGPOK+aoUkOcTHDdQsGmmX7/UNMAkyZ91/V2P2Gy1yR+wOv3WiEIdHDAzfp5CpQ
jk0x0PuKsXz021xzrWXezdypZGB1xVZdI/cCqBp9h/hWVnzcIibvgDNH/DEmf/bjCSFjys9DJ32u
EZZdoGIl9ew0xV7QINsmq9xYLuXThC/eLbkwoeh3167f95ZMIBIEAqLhSrHFC+dD4jdObJqhfyfw
IjQFyYgSOkxvjy/AiCKUiO/XjIqkyoigaVk+5JGlSUrMMuAUJvLAOVgh2gPWRz3x5N2/6UqAaKsI
QBhaQq3FwMIXnkzymZHW87d6e7b0WQRgT1pzx88H9OzBuKtEbYIyw3TYDEUiy82GCJlU2H3EL5bI
K7yaJCkXbcX6jkd4Bch8aMPEOPlz+cMYJZDKT1wOsq7n10QbeXKtGIc7W12PM/uP3Nbg5xH6BT61
Q9hYc3M6a7jnd5dy/IWntns6qqIcwuJRZc0zt+br/k9VhpajUx76KX3anoDoGMymQtUgdzPLaV8B
hryFElTmV1up0h64xBwP4uUrKHIUpQXnmwm8Znwsf2bzDDTVJ85iCiSFfa9PD7Qj8NU1IydQZEdG
C70neX6yK7eHptjBN3WAWSXnWg3jWQw0OR1ZhE4yc6s6EbbGGDddosToThID3BjSOxjSji0VQZa2
6RLvE4Z6IYGB8TuLt9rs/dtO1/X+gykWAqHz0iOzMiUjy100n2vYkik0B4YrrfzEoXlZBMu4CwpX
KPc/weE93QTJ3nCqV9PJQJu46s87bnIG2iz8geXw1G0fRhEamKJIE52IrOh6SfF5Ka/scpqCoDdR
CpvUe/LZATJYeKBkLTisIyjHEI8pJ3twcLRT1M28+DTqXqlL0WFj7stCSWu1vMH+BsDy6G9UScvM
I07sn0gXWHhcjdGeWSWrXqrDSrWQjYK4eEFUqI17wB47wHCOhTUmi8OpVpUyLExqYhFQK1zvJ8NR
mRvl/zRuUQtVh1buJ1/g4brIaUge0N3Zb3DGlkUeWBS55HBPmUcz7Uyx7m0dUMEHWlcQQQypm+5G
lkDsh8Ng+ADl7+53GURreHcC9NyAi9kPoxaStsgydERmziLW70V6thuV/tnhRVSv8vdbwililS64
IZDveGy/Dongb8sfSYbheWV/qw3FixFJ1g+PPMKnd0iwl//l7fZav6C3jZBxITgE4HtykmoywNW4
kakhFYFxnKJUXWU+S2qhRbSpw8FD+8g6liylGibDHIHUNL7mwTuovzL8hds9LMsojvM+JaItNe28
CXIdGiPQMz0Vce7HDk0bmSuTwIqCDl5c41t34M8LH81/iWQ8FRlEfyggQCRqtUN+sfu5CZXUH5R8
4Qt5Q7C5Oi7J7rJlQswm+gjBSoXE/IxALROMgSJcknpD+icwRTUnHGZFWZsFgryCgTK5OjiF0wcO
5ysIV7Vq+Mq5LYyD6LJtKK7xZZxExHlNdSPZLKknp6ru24qhGYBnZpgVHXDcakB1Njb7OnRZeuKs
D2WMXfltQPSnilm+NRarn/676fd2LRIkMgyj57Jg3BGEKPVpmDeab3WfIYN4GBxq0qELuq4sMOqB
uTJkLAZWIHTBD7SHaAT4GLagz7cFc1nh4q7z3uvp7jKdYQygCmW2z/xeO3Piov0plFJnwKNKUrma
tnHEqzTALxW1szb3+pCZtFtrhS2gVOA2wP2rfkCzk6NpculVob1djeQ9d2l8FS7ixVjT1C7mWu2t
bNm0l0o020jW5B2OiwoOhxBCFAsP0wo1RFNTy2507AT0a7We8AXvd9wCg2bVg2o99yfivH1F55mS
/IHfAqaZGlilZ7WlTeUMeJHtG0vza0lOvpmyww+X/iZnchW3aOMhFPbgVxs2AP4xxy7M3wrXi7Vl
eBHegsQJxa8RU8yas4pCaAIQIMJLkYCFva7yN7az3UtzhypiVYr5CTsNkovyzGROiDlEworORtjJ
l5a6XHPb9XfuwHZGKCSGXTF2XaSbgjkmxoSbA2y56bVYzg0H60jYYTjePQw233f5tc7w8qxBL3dY
RF0Y5VCxoE5JFdfs42i4J53hdAufMFFuN9vj9n5G4g+iYEal4/+SZCL4RdPMNdd3YCBHvYiDfZYo
j6m/unSxbkuYuRE3tAApGCZVu1N46GlBV1tIu9G+aboTJEtxcum5M/Lgtv2bhWItv8VjJGzzlH1d
tFJt19qzryeM16HAqiD2ShgNe/p0WjeCelF3S/3X8Xi3BeUMXIk4DQf6F+RDcnF/MwKSBNPg/YkK
VnyZdMYDy9pHIZGYy1FI3d2umOlOhYfSEwyA4s6WT7jFH4JTrITRoxDzJBYWLM9AYEaoSf7QR+pa
XdlZ7aa5QyIhGKyzI/KAAW7/rjFaQ9lV0C9i2ab4bzXwGGc6rLGP8FTuYGn2JYDGigPP4l3u+YMB
ZCMDsuWWvVMhci13v/+jtbPzndX7h17KxRnrYjCxdS6BMwlo/CrmvmI1MYMLbKaYvWb7RUtMlxK0
tVTfDHmxFV6RkW6cBSs5pZ3DNXPqBEKojvQgxoiE2jccS/H5Ep4n47RjLghtYg1BM9HLy8bFsP/H
p6F/mknAHfaCnwdJqDFp2o96bKZul/9fBn9QDK6i1ckwA6FK1HsUVCbJ5bmRo62jWfWVxmYYGJxr
iUU4queiwXr4ETGCAxy4Msh2W3YijzSFtznLJPRw3JuSIZ4CxWQ78Be3AaAaObxxB8GplIfvbZv8
JLgdyAJ3RErEgVotpQvVBEUx4TyDRXRT1NCq3ap6GteO2gg8BJOO+Jq923bMeW/mo0GIHpAVlpC8
wKBhHojEHKVU0NlSUZ64y+vg+F9arLMNk7lNqEqM9OBIg1ypMt0+DypcDL75dvGPP8M6br12LDNw
WesxPSKdMJ9/wrblGnsNzquYM3O/VHqwKc1shVChod0GX52PfqNXgVV63jxooCtMM1MtPDRNmNzf
SYVR6AxmCfcNzGCc6MWrt5rK/WCAcHDQJ4yHqfEVsnl/c/dmk7J7NKiSXtWMYAxq7F78KG0Rjtkv
ywSV+3cHnxO4swDCdt6lsVwBXDrwvWigXLTYCk2cj29Y+F27YGUW5dLSqGNMIOxFZroYW/bglkUD
lshCHKOJwRL6+hHh8k5KrxyP52YmS1KBd9jzujQADNNNJsumgTjIL6T76OVA3aE8BVUZRU6qY6A7
zig4JwgSeHUKNPD99hgHvbxYhqcAAPsE9/vCYl8t/Mge1oq4w8ZHa4iSDrQWypbbN7sFmt/sd+rN
txrMKOv1BzXigELZNsBvBJbDm7a8vIeJ4fo5zWwy2BK98RiP1Tw4+EnkEFashUCKk1EZXFniHOkW
GHqy6S5WqT0RRaI1COfbPplHyI+gx0PRg9vpNKiQAcF45lFzikTBINZi8nYzI7iC61kXCfpEAODD
jppJb4EnZB0i45EX/WI+e1GKHdW97ZvC293aeUEDfUOjORfTxTG7x7WqDCH6SZFJuyaxKLXksSzG
iF28vSI8b5u0XPdKWq0hLqFF+/cfk1FlCyEEIkSxEhWgcEIZkiKCNUgSd301Nj8HBhjYHemfrKL7
jB7YEREZ3i1AvrQCE57qXK190a1vqsPAlEBvaDFUaVk2bL4JGbf8YwhLz7xvJAWrDwR31BrvskoD
602vqJ++TOXDVEu7bwcOyps80oz0KOzjyeAamY4duy/emJURAYQpX4aNXLh4HRnz/m14/q12ksLv
DT76SGyNPL+bWDhYSx9bJYOVrei/cWnwJWzBPEFGteTYak/v1bM9EJnoXhwaMD0ky/crPVyeLsBN
O9sXtl3DNb8j2WNgxLCh55tgLAvFa9LjtwBnlcQAlEnvSfiORYYr6Viy79KkwxQtIeQ6yIhY97Pq
yBHboPoGH6uS3MSH5mHXr8Mc2494WO4gIZ/AigJFEPuBzU/PugVmKRylUWRtcQ4zxvCO/HrseA8Z
6Ina/EvTcFUaSXjC00B0neL8ErSEqlip3fFWEOLSEMMvgUhmpzKNBgoh0+LsirMheeR2lTHAqXDh
pE69c6soHi9hKqT6i+mfH26wi1M7hfo2xBfwzYZA3JoAmL7/HjNPMO75h+trfwooKUr1gEkcLtHM
/zBN/+MK2aOwbTny2Y5JEDpobgWO1Xtk1feR/3qD7W/fVH5UJ58vfscaqxWVKyG0ugX/eWTbqhDl
lzySR19Hn5Gyte3izGxFWTFYEM8JAGVTqipoJqKuZ7E8vizNHnVVzBuTg3Z8OuJ/W1VIFfighxbx
dbeS3K874sA8OIKjnNRub8Fl16UCbBUdZQrc6Qe1fdk/eaT47IoBRlB5tf3ZEYphwJBZtNmgqwGs
oMQLAX028fvjBcRNd+ArpcR+Xzflfoaq+2ny7e9ZNKEbGV6hnZTjsDue7vd4hwMe7EPRYebQiUOH
6yA/nd7YDREGXjBRCdh5jersgZMPxGtGURTUp2TlI27sp+ogxCtRrtDBW6RLyNXtrzlQj4kCTP3G
U7DKbVu9zftgQcpKMVfBr9f/4P7CoPbfJnVjNfl4KnQ73bojxmkNjbM6dPgV59vUEvJO2UnwEX+W
nolRyJRuKVsWRquBeEGYsQ+rhdWaCwRRwcKDL/m14hDT75UsJMhjE/qnm8Ef6WSpbP6xgp7uEgBg
gtdprlYJ4XCaXFVNwIqpfQfbaBmoZu+J3zxIkXYW/akJC+1KIRC2/cat73EsPEGE9fRJBUST0eNJ
4wXmc5sT0cwIBWusjdKWH2LECvBJiFeqYFrS3vOEasO4Wr9damW0GayhFv+mqjXg1zQbj+tcWasd
KmdIWQqfwlVur8wD99EeVvEjbjOIy6H7F+CXHR06wWI9dFbXqth7XfIbyvwYWSSS1MqE+G7tgLWz
3JZXwEGrhp+1E8K4h2A63ua0fdpujG6cQdGzjCaJwI9bF6gQOmizWCfQc8KNlg/pQD20IA7HC/5c
18ldngOPFs13IDE8JPEzR/UlD24cW6ASNdoMHLNyaMN0C2ORzdytZB9ExP6ncRikTSEvm/Fk4hLj
czawsyvY3SiWuDe/NisnW50K9Nq5tAO7wxtBhGO1htIeVowBigp5bd73WAMuJ/EYVV4Zr8hjlQpH
mzCTighFUVNwC7043hzg2ii5hZiLbSj53TGxzu2wmdQ+yIB9RDDHJdfxAUpQ/AUPIaGV3MFYHpn2
k7uYQbyNhb2+Vb4Ao+cV5PA+fsRFidyl4zs3msAkosHz+7kYLqp8CNcrBWJ8LwGU51DrvU0JV7d6
O39Qxk9VTlFmSV6t1dItWs+xnEn00zkMNJjPnIQrSnkky7mjuc480gYYgE3ESruvI5DQStmlbVw5
XHmskUi0FoumQkeBN3Svz+7asU4F34esYq9nPoKaLTiPE/16Mgrx9najbJLz078l95whjsqUS3VJ
aRJ881YuAef3OLx4qZ8m6LeRwEkCTdg467yQG19zLLuPdBtGEDp8k9+Ksvve/AIfEsQ5R/1bVJdX
Sq7/vTfrOA8z5enZcbr4uZgf9RS4LWLIUv7s9nZbIbRmNagQi8Mkgk4mILP/sLsg6tc5yQzVT80s
J9hPObXnWv8huxnJZFreQenUF0QIOisEblBDA4EKkTRBVMkjWtbYpoWDmsO31sDAo+5ON/macHn0
rjvYrTX0916KiQAlq1OgisAbLBYeYZVyU+2lonneQOhG300VLJLkD4Tzb+j1cWc0I02IJuikKgKc
UfW1uZfdFpMX131bzOOr36hkLBfcmytKoteqvyJHfz/oEijLnm1jr9DMWIwLL++/dZgcxzNMvqzL
91aqWuVAbJc8CxU0XFF0CkmZtAHDYnKLujlWNM2O7UKx49aNONiy55Auhp76ZQxRv8k3rdWIUbfr
Ea5R6q4liaOH2zdtMfAAmDSs8AxTOgbH7xGxhhMeYzRbl+lB5M6sucBgQGhcZzYQhStqnOqSS0zU
AV0JARS2tKT/wOoMX42dfJVbfI0j94DG3A9vbF0plofGhuVg/YQlHbLbryqnmPb0fpQ3ozyLWQpT
nxdf3WzVGQ2L1bO1eAh0smhYew0tk+n9/SrzjLt5MY6t4IXnJOAnEYf8JjCua4To7cEyI8z0P9Lw
26PU3uN3EF1wijzW2ctMWVmg0S7/7A1/6quoDKdA83BdE5qEVKBYJ36PuTwCH+BhpL8ykPJAQBCZ
klV9VtMEk09kvF8RWa1nNzg9E+PGICjYsLBVz4Hu4442yVnZf8kT4FDUREza0CBvMQ9j8yIbfM8Q
c0isRXdovjUKFXK3N4fRro2NOBldE4oenwmE9CAvLln0AsBep++c7YcqjMYFdPaJi53JhmUoKnXZ
ZrxnLlv7tKtHmlq8Wm7MkJ7OSdjc/uOeuDFGz1HHg9EJF3K+xRVMrNYUBSvqBG1FYfLaOpbsZ54+
n89Hluh+1lhxcw5+IlwfM+L45qC5bNVokhMTOefvZy5L2DUcf88u9O+53q5AdmfDl3fUxLLSqKrV
1f0akQEh7idUymnCtRmx9qeInUhoOqXviuvxCbQ4FAQDDWg9VNUI8X+AUzwaxs+eDYYWvtihBJRn
muyKlZujKUMQgQFw8fBEMtlGPI8PjqBxZDg4wniJsrB8erxpFKbJ+pN+V5pYbArPkx7u73/RitGZ
8fvzEiYYLrgtlbuVK3axwW9KUyiAwOktILfRB8TfIiyeu4PwrfMbN3BuKxka41PVSUee+G+Almhn
hHfoXbQQzmm5cdOTXUO7x7f64AgknWb1Y6fvmpnbu6j7NOr9YI8DXzkL9h94k7L2dA7ItiIh+XnR
3MyBMC/TBWtQ5qzWAd7R3+Oo660b2aVivuuz/g6pYZCUFg8SdDJXGSmLj7Tm6kq11Pu466XfufLj
mHH5Umi6Q1Z5TGtqOMSXzx886DR4nT3BJWYWQIXJCjGrZUJuwkh1O4tirGWKevSBDUnldtyiMcDz
Gi38kyDjJogbzIg/MY9f4ib08CevIfkRXoUnJRm38m8Hq4PTzn8VyLFV6aGpaV8AYxxqiMlveswd
HYsP0NZjNcTS8YyEoI07jLHLJFZOSqF6LFiq7u4gXx9o+SwMPO06wfgNmA3IS2pLIsNjXhKTT0KI
55aCJTHkR+Caqv1uhni+FQihTJNsa9embFpdLLVRnIJclHIVnd4CVguLUMfOlx3nVgOy/YXkKvJx
0N6WPPmW5CPZo33Ka6HfeyCeLxiQgHpWlsXQKOke9Lgzcz/ikxMsdJvo+D9Za7lwOpxm9dFMkQIr
yeeHJPBLAH12JiRvKEO9Js8ysjzZDVhFzc6tfejOK6nz/PE/FxKiTXb86ms52q9XtFoLnaYU694q
DhXahQ8bwtmqacOsn2E2nUb/9TdGKJ6FPlKikYn7h4ykC0gJuFCfzfhAyKEbIBEDbVEjmiuvFq7l
K/KXWa0o+3RtDnp6cAIMZJMdyPB2KJ5GnfZMHeFvKkyw7EbrrGTDJFFUOlkiaJ/nw8c6A2F3UZve
Az+w+iLcVe8yQopszbR+4arheowolDhaO3vMdqiArV1w1cmfnd+xGZMB/NCP0ZMgm1igbTblV8/7
o97sCFWzj24vSNxs5mg2XCnzx/q0YzT8KIw8/dbNE5cO/mBhFYxXQclEUZfCdKjk/X+OCsQ21WqO
PFrU+FrJnZkpXCH5uCdG9PXB0eMuMo25TED2Fk4UrP0I9M/0kT79sx8fnJ/vK1ATMGQ+tW7s4kl/
4lkv2LlYTy7d4aa+dz4+KI5cxYdLcGkspKiJ/a90ypy/ceqsLPd+DH4jAWpj3JGew2ZpDbugGoOe
CQicYWGBIzoTy+aHVx+G04Q+snHZHymZqMZaKhLPdLjQqkZkETzblnCswnFFWsbvIseHyufi8IaY
fZz4oqWR/HR4R9oLi9NPHVCJe7s9pNxOjnJosnk3LgJ7H/FMB2OmS412tM8lCQncyRujuQOErlPu
9sOgjxhst1rPDzY2yaOboog7L8DZst7DVySvclFJdVxWnSYsOVxO1opSZk76RFlliiaD3bUd0XRd
wFH/vIxwa2IcGjB8AnPWiDtlVmQuTvc4I7wctIklJqnDvMGpudQ3iQ+ArPyU43N6AyQmPLlzk0mS
htyLtG/cIA8zGkPjZ1/yJJog5dkq426Sr0jf1sjSf7ZteCNl2SFICjCKOovX9HCrrUkRWrajqBjG
v5oB359aKtUd++/mh7n9wWFEcxNa55MyJEe7WeAgs0ZMXGl0FDfgX/jEdYelN9lh3qK7xGKlkfg0
CYJBfx9O6n3FqnDhAPfjm452uslUOKlzvvLunlli2VosEwKE7avSamXBV2G8X6N/CQD060vFg0Fp
KRJkjT1wQqSPp92q2GBt8z+fNEikW8x/+tAvx0DU+DwSn9jNhYpuqzKqpovTk1hJW5ZgPiP70WUv
Xr7Zv0H9WdgrbShUmpu0ZtWYqPWbu05GsKPzNbo6fJ2Ov0EMDAl0y0Xp7F/AAzsDvD+Vns75NPqt
PObTrd2Q42Pys0SMJpuUYOrKsVSHzS4wq/kKnOI5F6viBZ/0mZOhWNM9Gdp3TV6mAxw0Xz0iHXb5
Jp0biyLtPgJXAuXr8kU5qNXsLcWtkeGGCO3DcGyEa+FRyA/r3JhJ/DMeFksKTSFUSKGFlk14S/Vy
IhHs9vQ3UyDFXGe2q1sdri7PeCmzMr4kL/FXgwCERlTne7rXG3sGeIrbXArZoDq7j7rhkUDZaFHI
AKLu4LEvX60b3PtIiUqsa1TKlF+ESsH3hgKd974k/J9r4UyhdKq6LQNeMkIJ+VhlqLdlzLbmoL6Y
FbSKBDcgbhaToFFpuIzQLI3cqTo9xS59MOzUaUmMQZnc+6tq9rvOH1ujaXjBWc3o4py+Kzau8hWi
I7e/PHRyZ1KK/WbtYi/L+6LdXtb5c22z7NX9YtwwUWT4WAMLwUJFCM6r4N53PwNj+2bL8uPKLdxq
naNEeCaSYfaMQegN3pTeQ7lJkXR/+fRfHe9s+SvPbo0y3vsUkPN79GkKb/hAIQ6wiTMN/cVuIH8i
B+oz1woAK/TBQuFOSwrpYUfyoVE0fd4QAkBrGGu0P/4Ba2ruEgeytDsxxOgCUx1EA8FfOJbuxnHh
a/4Rpz1WXRhAi47O9f5CXYpYLFLRdwQTi5ZR4x2JvAFOEqamJbv2gZu53hWQRS7iXKRayYU9gn/E
Cv6sDasRkKeWo1LC6ZcY/vgfPH5mSo5vAlFUILaDKwHlbEOdv+9r4sfnBzzp4yxvCH8RZtttnYiz
hOn1ZhtjL3k78zsaJwq3MghyZRQ9+w03qbaQV2aV7koCKCWTZ38EJ6EyEAQ07gcrj5cK0XYouizc
V/wE+KwuEoNGgY2XFYqJRzJDrzzRNDgV7QfAbrsclDOapBv1OultVA+Zqx+G4Zp5Lwrp5AqAorpk
GotA/2N5eREYlIDyDcHNCjRX7bNWl06KgsVHtFDPzIF9Qvj4UxGJ8ykqy8mfsz+IhmnY8Xu+PJFS
wivhO/7Rc7mXFbRB7jKUnkAMNbcgMUE5G0qVL72JwqyK231vnuwN5gWduw4AP6yBXC8GiRqOrLcq
qQfM2x4pkx7wZJoLZqof7mSGJpPhmpUIv7ek+YX1tufcWqRVTBfn0WEPCerzR98lZi+HKCQrBQpr
F+30VpW+Ow5hcKrTQ/ZmGHfbrzcYiUUGJBWmtZs29gtd2QcMQ96hGLdUU1qlAyBHwXQvnux2uTKq
HXvnDr7UIbwBA3lNpvxxkTErVz7ZFYSklDnGgTFZq6TNIrig755LTzWun/7Zh33h6MDTEA6BFR6G
FAAAzZtHJ48eWt0qS4geuw7aZPdQZ134dCw4AYFB18X6z5TVFz6joqXosV7o6b7Aj2LrRFWNQaVI
MPNO+oZQVFKj9JLKRVdwtRmQiWlqPMoVMTxwJrDOPZQzR64PePbLH5pMhd6umXQ5Lmk37gQJ2hZE
ZB2IezudmPEBMBJYHPJQkZ1yipp48bBhsV1/C6ZEvgnSRC0subOCkgfcEshgoOiuVe77JdBeX/8u
luzQ5/I5Mvx18TiCaYXiaZjxt0douyA2Okv0oncbMszT9tfiqhpiXi7El1t35OmC2D1H4u8ADcmD
PTPzZwzeTyXDgvpMj+ebCili3qiqcPWzzqVZwQsqQXEiHMGkyD9IZ9WBQOCYP6TBSVm922k+VtKp
yaSLsLSSxNdnBV/svEWQ27v+SdXrtzWTwuKnaiWW0KtpgQUR3/BNQl/nvogIJzVJssGx1vmKB4Cl
ASctcwk4YEOSugm7niGBUeRHjXnS7ziibW5/kGPKRCYl/s5piN6nFfsfbZgddrnGFj19yc7ilClt
zt4Sh1xSrw0NfzIYmRxM15BSVSdIdPaJOjUf3nl3gIKRO0KQc0URAyogAkl1tqYeifTkfyvN1LPK
SofO6fvwwuu5cr0o6gcu8a/LUejJfm4J+Fa2TOYdVx69l+aXeAvcmMQehX1dsmaxK4XdIB7FZolf
WT5mKXijJE4LmxvFCecd5Tccqc8vDYv0vhMIL53ksOLN9s34mX8dNSEJ8sxlZCfx0f48PtVA2K/4
ryUvjqBPRWzvxP+i8H1rdEBJMElrg7Jab0YKepV7czib0JYydy0+HQEEtUNDUdAgLbixxiiYElH+
RdJd6pv8kyryQGbO4aJ+hAkGgy9J5dvIaemo8CD86MRfQsKTKXlMk13lok14KGrMmfFZvbg0tMO2
dqb6m85shNvWNSJ04+GUztNGVIIWDcaUfIm7BaIMVKRn1NZgL/Bl8uIFO2JRhQZZiBQ/jGXm6JKQ
oLsCNawbbnpnF0hVzxNW2Qvry1ZvgaeGS0XQuIbdDHSm6o/wtRU2GCq5UpW5r8FNoxwzxZBhsJmW
PApfjRyflMKjM1+ZlDDrBYmu5jJ9pluE1EG4N9Yfi5WZHgK4YFx3cYQGOrQZp9ODseYiAzpeXHYY
JQYlOsFg/VeeDnwFg6L2Oo/cLSxMs/g2GZghVig31xzuLOIMyc8oqX83DLsQ3xf3nCE8TZ/CErJy
oD12YB7pTNMxQdcesMJ2RCGFcrMsAf/VpvF4b9henqHZomfXlHfyB1b5I3ueSNDXGdsi6E/ih+3P
mf9qiwVQF7/U+9uaGGe4tG8P6Z8WeiUjxPgZI68ViQqxSVdpwKtMIplsTGfLVBiShZpEKbLalUZG
N4C7B4qH+jja6zP0OGyDaXTyjrIJUPFXnYYEqOPIVCeoQI5OXuuFy5onGc4uSy2ZAKz0ZKCGq2i+
o086EsL9TIDsp0ikqMygq1mQu4i84H8jJK0zcDEHpQbEK8536o0CcirXSrAkUnJYNYqrYj8DTUKS
XHzKoCPXSFfoeIh9SYQbEriZw72tlJQfz5jX7OY/oqLXR7xQrD/uXaVTRUnRQKdoLVCyDHrphbTE
3BmJZ7lKs8ehP2AvgFlOhsQmWTRx6e4s0ak+S0oQ44adQohLSw4TG/cKG6xbl+YBW1trFBb4KD7r
TxRxL2YbU0eWKxNvmq8ILQ0I2W4ncIzsGX4sO2BXg/sACQNzZXXUyW+bAOyLtITFUFLngzbX3BTc
1grNCsG7EN316vphyUWjkweyyGop8QECgj036rHbgI99sC+BX2SKVt2bHbMg7bEIh2RH/WBmS1Am
9jV3OW4Xtfb8Kd0SJSeaE1ikzYiyP7Rn75Lb7LvoNaeGXsQMlmNjf4nTdTpQFA/bIzOGk1v+YWp8
/G6XEJEfXTd6y2UI8GdBkzxUrkWhO0paVOt5PKKzesc6X3epStLw5kZtW1vMBWGAmmyoY+CsZdtf
mKUNzIU5Tg0/90TFIAnR59WSp3tZ32YrISj8YjPAfhQ7Nex/1eMnz9Kq5w9sazoPH8vbwjgZ9AwO
pbFT4YNid9GgKeET+B7Pg32ykGz2KwaDTx2zittBkbTIW4S1WTmVBSEBJPfFXHD2viFrZ+3ppmAk
JJIDbGIEUhr3JQV3bJps3PXiIpuLr0ZkXeSmfGJGOWuHIaN7fylrWybozs9szYXA8yR2s4j8dIHR
87Bl+shDKZCW+soxQfH2cVYHwWBd/Npd8WAarTfecNIbTTAPvBjUZxxDCmC9NcKoLJTdlMWLYjw2
Vv65wkIYNdk1FT2P73p05bN5Hw/MQNk1/foLddS18+kcccOB3ROZocHjVLUKLdD/uQ+fD/V/uTTY
AyJS9sLzaZ8G9VuEmCLjjtl9GQESwmAA25rDu4vegZA5kvygjO4JbhCYHTSUdsd1RT6SQ643DYGD
O2VJtmyCygQ2qkeQViOVcaBXZZBlEypXU6VZknW7P1KbrPeHQA5OTUQxMmoDH1dKCgO6bBxonkSf
Zl+mXxdcrGg+4urs4TXrye3MJW19PzXn3/TtJkv4l7WgRza9xOLl14Uoep6ZCMlAgl1g6MXNV20R
0kx0w1hdczwbpQicRiFcmXHC3ixMn/Q14ha1jKjYkzSP2j0yIK2OxACfbXDTEsnBMv+09apuJXvE
8o8yFTlbzhUG7QTzVvZ5ReMf8zoaCNlnJqjCx7L84l/fB/Grcl8yFMhLkDyV8UsCqGoDfjAPN/wG
uxq4j2FzMI+N6XcvLk+QlqDQZkr/t6HmCqjx/MXSL8Qxe0X2jJLOseQp1Ay7433DhRynfDb/agtg
YU9+r9sWf4yxmz2VVYuRz5ijy7zTQaWIMq6KCNgBU7LkH0z3NwH8HKhaiTO8wxYDIDT2bgYOwXnz
GBfOrS0dAW92dNxwzWsyh4P0axAbWfRtvEhHnisiAIIr8DOkf3fG9OLGFYzr+zuauvq3Blg7kJ9R
SKu0SlRAH4anmiDvA3HgARUjyTpuJbAtRzC0ymMeotrmA+66puGl6ideKoNlyhPGudqUYnBAGlR8
M+P/zOx4l+aek2aJYwrESlXgWx6QvXIWmyb5gbFvpmACp+rdS1cImh8nV0966CU+49owCvOjyFgU
5NDWf6XiKnmvpVThEkQhlUcq5nI1yJ9Jysj9XccNdTp1FD3IGASG2FBO2Xxhmr0p3Q+kkMSHyGbk
cTszGHCWNPbsoIoGg8PsReS0OBOvNaCknT0HkEFqZDQGCgqoB3Xj9T86lFoluhzUgjmsFODZJ/ex
TNn4bWhnQQT6pkwCw8dcW1TKWG+lkIejnz9RCVSyWHKgGm1GxvRly9aSIR6qKCzkKDgG2YWMyE3b
UpqjXX92nQzI8CQ8CZfq51L/0z+yMFZoWyy5K96Iyai4uA/qrAoTKX1oYQu5RKaoGa4m0M0rlMWx
s4YX95vWkjkfvK7BYsO/24N1WEHqxHIvqPKY7s7i9L/SH1cqI5leuwrfr7xhow0uv5jDr+ncT7EX
kzVNS+oE7k/FiYqIfe1rnqe3uPlp9ilKubT11DTMejuvoLIU83T2ga3ahDQnJ5FBcULwl2SlUbMx
RgP1eXK/9RsETH8rpLkAyrJxWHGBbARtXRSXn4FCspr0Fm1cHPoajtOPtKPP/sXrGt6ZZBfFaiFU
q3QT8p5K7VscuGG5O15+GXfQ2H5c2u9v8gLj2dpZ5u7BpVHjJHTCAjVX19FSeKIVdxlOOIBjBVPY
NnEfEWu4YjFLQO7TYZqVPI/HT4QfJfoglpTpWAVwGXw6xzzxjpbKsk43tLbp5KcjZbH9HLTwH/8t
2XGKRS33de2+dmCObKcdvWCuYiNaIEI+P6nNgIeERgYCsO/ed9amq6j8DIV56qJZ/3e3M1woax2T
6kbn/UGshJmOeowutBthDQTqfGEwZKvTyDKITwLXwj5pojnHENPRIWzX2Dqw/C5thlD2KglzQOQi
h0QdEXBGCH1Wc8YAGghqKEpOP1HvmxQOr7Ib9AYMlQIn20YeJYka4qiqrITpubFJa/2oPsTyaQ5W
HebtpS1uwIefQRIbprUIpApUXWNgN0jApHvCtk1sGVs+H8jJE9y3V74twXabeeA6B1M2tqtYRf79
/wA/+NtigVhnxrvc5tgjpma0oEN5LONOPRS479VhH/2SHQ1M0naYE6dMWf+IlTHkB6qIXnmO1659
x7r7SYg7sdl46pVgtIPgeV+WlwNXFENgceyah0G0l1HFBu8NJ3Aq/B7OwEYOhE4IA4oLTyKAXN1u
xpa133ICGOTN9d6jkOdeEXO2ubwn2xplQ2Vyn2cops3t0cI+ZNdO1NW36c/pIz+UCX4ShugroXNX
gulJZX/CJGzCA50deGBxUe1UQnnNgOyy12f0Iso+oXTOBnVN/N+hBIJC6z4PDpUNDr9qin2Z8Dwu
KI3wmqPfJjCvbK3UWyIGkb3Sb4jG+zQuFnbdtAd8z35TR1RUkohRmze9nojn2C+G29sFgDLEt5R0
SBKJ34YqOH2TtnbBKi2U1+WCjsjJYT8j8KeXVZCl4bjkErTbQrcmk4VEnTXHVLfGZosTUuPmMPlU
CuyunsSd/M2xPAD9f/z6+X/o8pctg5aJdyKuPMjLi10R3JBHK6Zx7pkAfv4IGKuJIw4F55/ZoXcp
8/JKisK5MEBfbA1gnGWZxgcKrG9tFqJs2IWyAwMz88KxaOLWDXqHatUHMlkp3GavezrY3ffQ5xuX
D9ais9Wo+/bLWeNOfz6U5uXAjcDhBwp3apnd/8gIOvcCfv9Mcu9XXVcCTg3dB7NhtCaVVpe+ZhyT
ynD/KY0asReFQZVwRoKA83G0nWsbHyra2K+SzE4PvrIBKfNZSrhdycc4oJkztiEM7pJvok6TWo5V
ewC5h1IZJ7ueHHH9l7V0+EuKUY6jp8cQ2yohgnkpm3cO621+aZkOU4dR/bQsYSeOCwMYCUDGOCtK
3pIZ5HmVf4p2WcXgoX1UPSOijIYEZt+xbQM3bKANwJaN53UEAEMH9ArShxdzlTeKV/92YYZbl16B
cUaZwaZ/SNO+QN+L4pKEoUmWDdZ/S3Uam7ZiEQXYR8h6XDd9XkV3zISsbbhSLAJSG9h2j2WNU4+R
LT4+xR7fAoHiiCcvXf7ryyPVduEFK5JlGUM2OUtoOZmPdZSmmGWheBNjw7Q/RQ86H1CgPetTLu3G
vd8L9jY3YZnW8V4e8sgUQi17Cf6oEoPlxmyNnPsF9F2U+JEcXgt+24LJBT8bB137/Q5GNTkeegpd
uUMM75Sc0+v9TnKWGXmyYFh7rWM1+DEUpiyJCA6j1tF8xgRMFrHBdPF6zOPwOq24WrtiwpTEO5o1
a8YamnWDog+tVUJ9Yd5dlRahbsngolTIBNsAAq21p30gD6O1+qwtgsxkiwBjw/K35jadLv7k9J2Q
0x6fv6yv5UOviWtUfmIfZdw5h+Tozw4iHLl+zNzSqy4DW9PzOZf8zAPrbCTYXBv4Tj3lY06PC9lM
u8WvJxNiSXPSXln9J81FyExioEouN+96DalkRCGjCNbYG8Ay//RKDNrcrrgbN2OZoZsl+VroGu1l
xT6poogVtV34e0/lkRxLckz7Eyhy2KOZkE970N7720/Z6Km+cUk58C8NL23lQ4FoASSTGNWePXs5
B+xCCv3dL3teSasQoChvGZCcUqU9zgpImQ9R9UEqjGcPiBqrAN3wsDEHTUgAGmrMgt0upDizQ/vh
vIAyP0TjDmsNFbSHSW/IAc3V2dbwrUvQtgQXb9B6HrcxnQoHc6wtjQurPsop552nriej7/XxuyQH
p7xnOOBB4aFYGLWw0Ak/RqaQT5qfLG3u8YRYnzerORSRqFc8ZHpaZpgGF/cCXAWvktLG8wKiXidd
6F999F9y1OMGiRb7Y6f9jBmQQx8RntWBHOGI3NXtQE3t/bYnUrFAQa69grwotGzwOlAg0gAuTAdF
brGz5X2U63CbjP7PlSkjbt4IRsiOGWwsMoOxdclg4j0lJw0fbX09C8IWvril2OXu38cKqtEIWaw8
yv2UxNzzgXzo2Vg8en/8Gfjb66n1a8kpI1idej2g5/PDk7X0ch9c1/BLBAdRQhhfktSQarlzIePb
+93duDAn7mSjbVif7exTLFY94QAV80xtonETN6NdZg5883rZrpFgod+pGmSUPDu7AnHUW0H1YAim
Y1Oag+39r7o3vu1MY3rf7Go5aWeBR5CdleQZPkxgNjTfDN2mkyZAUh+aT29lTGugMNDazIHKfXlc
iZDLYi+U0664gce4KDh19ENKCmWZVmAQhSaMyJoJoRj4GtT2fTYdNXa8CY/SGJHC77rhO1xOS3k7
voTpTeiE68j3y7nYMMcf252uLuiVqXOLCLc1J+eV7t5XSrlLxdO2YOe6Rj+iJmQlWJCECUd4m46s
djLgBBGcYkuuQn28YrKIhRc+H33LaIigERx7OuYwxd6HqtPcaurj17LS1ZYf4vwyYGTBhQZH+E51
VrqKHOu2hxcb0A3DK9+s3V7bQMuQ32DyrFB16wxO8JI5dWb5Bhy+b+iY7NG7ucQztKBi+JwhKfXE
Jq8XKNTTTDXuJyyipdWl+rlf/31Pq0OmZvfr3+hwRqlfuk0AeJvWMcQGAKzy+j5c1SIvQw9k74iK
tieGk5/quntQJ+xLwVOJgOjCz5w3ZQTm4oPLznmXKBFxSNmYhJkI5jMfGA+cNXliGj/xqOVpx4iH
KwcY7r75+sftYNP0M+ZZ5OOeJX27amnR7TnjY3MlwIlDhDsEjY7qiftphswk9XBKREIXzhqE4eFK
5LP4dTNESAlwLk5KZ+oKcWcvzILF71IV1lMOcLmRgkXfHesOjcpLyuTtooA8UPEi3jlSOzRmNnEN
y2WfRFMBI+8exZ/e9V/OYZhS1+AHlL+0ZwIfsDtVvi/tSPhzK3444sS9G6uvcdhNF2mZ8qVQ0OxM
YVbNWnby7W2KEeQPNvgvRrZ6wclQBRrLzqBneeXb3gflnSttZZexiAxufb8WjK5qs2IC2cknaTkF
Rz5vWAEQgjv94Prx1qpxJm5FOzpwCItOfY3H36CnFtQRuTHW1jAuApw3IUNJEqPvMU9GjJTvVhiU
2QYyT6bDtmDIKp2Xe7BGIWOMVg8jiE1CDgS6z7f5om6m7RLY5XCKZWinkwTW8h8xg8sq+2xbte10
GkLcxKh8Cf1Ac77IG7nmDuM44mDzuueoeey966Vd9v7cv+mFQfQAKErVJDWh1wrWPomqCULGLLsl
RdgG3T9qy9ODQe6NAhG5432O+2aJaJuQTMMxZSjYIbcz8Xi9mQ6Td22ihoK1GGBPQaJdW+tNUAYc
J/4w0NBvxZqjIu/vyAcHz0u1eGrluSXpNj6URjt8zXOvpHP1AfvIZBeJ4zF9QXpxRPoC2G5wkt9M
oF5+H6lw7g+qcTWj8GAYiQPpbuwbANFkp6iW8nop4AKq/IB9HUk5TfU8e38jUxVArA33ZF6Ch4YB
yNDOHlw+DwmWR7PEiJdEUUxBZLXo3h2HBesfX3wVXMKk8/eVdYVTGuEWykAU3M7jQl4uhFB3en1Q
ucCRX20sRtHWzgNcBy16ShNLlyx4xBhBasPsjj3KuPNZSsvRGb/K+5pB61ppkk+jp6o5L8hNT+6r
tazXq7StNqogNbrqMjzCwLlDwKbwJ/+ja7x2cpERFGtuqyqGUa0jU4oanROdBcjDNyXiE+S/G/A5
aoGzVGORW/fF1mH47zZf6zI4N8TTVya0cq3hehb+fgGVtkmVjzswb1sE0dHhRqLDYKfuznp/634r
Yxv7f2b/9dfhwaoiwOJAUGNAL8UQpzBlUufYaKSYO0/TUFrN3opHqRkcMgVAsVYNK6uR4w2oiZ6Q
TyB3Dokax14LXcANofHDTr4gSjffZ4UQJDuGrfbC7ValiTSJPvw5Klcuxm+gVo3ow3Sr7mVAniyr
x3smGJdXVBYoIp7APSEtH3nDCMAbOyKd1Mwl77xnJQ5hyD3WIQ4h/8Ee+E8jjVvVRCx+Tig08FFx
Bbrz6oDbw0vz/alQr8/p3cp/KMGQWlb4VSS7OWv9VclwjulaeeddJj6GFFvUljYmTGvS+cGFiZB/
x3Ew/oLKqFX3W4HU3Cbhl99H6b7ukmwIKsUKojGpq1pMvzRkVHjwSvbsycWOYqdHutpLgds9XTat
LFDPkhNRHJpYr8wKN9aEkq4drXzzny1q4w/oGSia+TqOc7E0jzWZRA49MjAQYk2qsz2VPaaRpjR1
5VE3erglN4QTGvGgste5v2huMj3rqVphVmhMQUiIM0o0UiQaaWx9G0NqUjuAlfEoYeM18DG7eRR2
PeeruqyNSzdFXw5bo+OxldyYDMmfY8EUAwlhogPHAoalmU/NgMb42M3WlMBdJ9IqbkKaQS2OJi+e
LjF9QUUGlFpjtKXaGydqdumLnQVnKkjr/BjgqzdkY6voIkz1m5jzRBiVuvr8/nriJjiIdzU0Ydsv
aq9OqUNHpyV3gFJTu8homihqB/9/uiVTHCJMf1kMYkUbm4q125dbE5Y3ii4fyq5G3nj5cyBvxX+q
Zkx6UAvqlAG1m2SJIEk5aOGz/ojIoOfm4Lgxi8YbppkcQNpGJYRregmc6BSbe8cby8rCVtknatS7
WjZGmFOY4sYmxPS4a+Bdcy9AzNBLALIzOYpV1+t4dIEIlCQH+oP7fZxVFtiGUMNLTMaAgc+KJcCi
BSIWEqXjoKmarEg9JVFswQzAfIhXi1q9yRYba8xWNYftHAam3WRwl0xIyVLPub6g0s0O4djYzk7E
BR8Yuyt4uW3uNEQkoijzA97E7REK/mlD3imZVZsIIBelfZtW0KAY43BAgtMNwzTBCPuQJ1hEOzhE
uWvWBWVS0iDCtq7sFVF8KnMf1y/N5xoBiRZGdsA5kIopZL2uRnyGpyvXh2mDvnqs0lG+9MOKybbF
9/J5qfM9BtY4BxmU/xtIZs9Vwhpv7+vw8psbH6R9sT1RulpwlHkjXCjDBbnpSanjWKNWX/O0erDA
40+fB/NU9Q1X4PMuFEoW9o5UrNkRM7HwuqjRU/kHMh34PSiCzVidZ2wXfYxC6WcX4zrBV9eJ/hPU
LRoBWmsPOdHxjcfeNgiRu3a4UNLEJDAq/yadBKt7otGPShiwZt1ax6sdrluAUxmpPihOidM71maW
G48QUAY6ZKA3Aspl9lruL0He98dtk2L5Bgl8PLDi9EhdQllooBz6Fx0pVp2edAm+bv7koBu1NfdS
8P7A0FBwRz5Qzk+gCI3R7QXrCkPr+5/q7obXQzsS4QQ9g5sshxbr4+kfRWVifa8Pz7bY3tqgswmt
sXcABFvZBg55kGSA4HqLgPUmLBhapZzS/T1XYiJ5qV+b4oTLr2yJ0n2cc4y6JMPNpQXvHS6T4E/I
rK7kA58JZr6Vk6G8SnDiz9hGIoR87aK6tpCvHJWD8CAHxTyHOLYxssDsL8P31qv+B7Tttsi4GECx
3+mf8tWiWmy3WbltiSLi8EsAAI/FTQNnzPQfFK6127TowEZG76Ue+/QYQO99+ZJ1NzIQ9SVNCdV8
HQ5DhH+XuDbmXrAj772BiyJGLMkLCRqSfxFgjH0/cVvjQgrQBFYZzhGatBYYyYz31ID2QDaiY0Lt
cFTlJoDyqmtuUgGLIFX2ucElhdo9eSN34JfqxmDJnZgEZYZRjoIBWXS0E8tvpXYHnGYFJvysTsgC
8991+2q8MnJtaUndYQOtAk+qRe3jC/dnLi471K+3Sm/5gg44H3DJKzFH7DpGpiZvJxLM/wsXYQtr
6dDLEBP1kySoynOj+9xw0nDHy+9toRdNvlMkc8vogbTdAtIOzypcBiyS0+fte7OX0QPhwYBkBR6t
sYP29ceIclkDnsL3KlmvyiQe+uRsXeS7k9ZVjdSfTLeS9ZDBtbxHPkm7xhagh0MCNyBUy8qk/zdy
UVS1W9ZHJHA+Ct1r4kf+Lz9uuA0h1PGwAUkYMT8ti/tmAud8lhurSRxK7AhcJXUUPrSj57k4iKw/
ka32DHZHIliAYsk+krIMEq2kCNXTwrW633ehRajd/IxYnMTbhsj+Rk24+pg2ZM65c5oZR03o8uQw
Kl1xf4VvhqB4lkz85aAGNRmnaBHw55WWQWE7RMmp8Fbn3x+r8g3kcnOls85dG6pCRlVv5y4nRelG
s3+Dzl4tth4eusrW2ZvGFpU/4hagehgXLCC/C9qjjG+Y9zCI7gdZ0f1/hrzd0mwLbjuLO6o6EAVz
AS+82h3rzK4wYi1jS+vZLq1wr+7VGPtTDJ/nec9+/xhATFwklKaIjvlrt6hOI8MRUg68fhuqjy27
bJGV5Tymqf8IW0pXvIg1yR+2AI86wTcxdW9ITXoT6r8sO38UD9+cQxXMTgR+wsEGWbq8ybjATQVt
jaspIlVAl4oTQs45sLWElXSD3+xCBy28m6vvoUsXMe2oykgZ0k29YcUxugYT9N+WRV0KRTAB70u4
s8Vn9uTtcNjWvDCJZeIemE1cC/dQMmuPhCigH7Na8ZR/yF4wjJfD16wnkOGVjL4VOWkOWqPYf39u
wFx2T/xqxttC69/waDot9mwuG5dEDMZNctPXoCENurFqvkZM6zO2VNzQMDMeupRDYav3UMHmUGXd
lz3tryGIsMnb7Yvbp+kkv5dFQbzc+PzTXzNr6AVf37SjILwtU/CDu2Qj6IWry62PfNy1nqU/E7rY
mRrRmCo9hgU4iO2i17NtvSwM/CliwnkG2hrD1exLnURRPIDAZ/90yWsYyTX3fizEhdH8uY536ePQ
5NhvKhRzgc/SXF63TjQqSwTlevyz41ZpMEQU+Vh6RcyrWM+qDNREJhnKN5WVizxhUWKWmEV5Rn6z
MzgjBe+VyNsn+vdnyU/xNz9eJ0fmD3BEFNzK3BKnBiSkwWmo0R6o+vG0OIgR2lGMZma9F3xyht54
Kop8pEH3mqFi8y13MWNnp48O9lABnpmanX6fBqMIVXn96kqWNystaqu60Eop9wUnIgtw9sXIZqKc
ciPGNeFsgTVi7i+jaWhVcYRSubi3XRcxNom2eB5MK4UhkI4Fd3YpTugTvggjhOj8GpXSfkMHh36M
uBWKlO/yQDu8Ypy264hz8KJBqCKLjSmrjmhVeFARSAB/iVZRIU/NvBCVJaPXaABtZF6m1y5sx71t
s59t9nXu0z+9ph58Yl8Ioln93G52Qdpo04wK2uHOIjmXuGJHAgZSuQ4vKKm613BaEHs8u0ab1FzA
IRvlofsF6bg7QLSBETAZjgUbe5AR7yqgyUOFqW7PbR6HMMcFnzN6S3cQnEoJ5alOwUlW5o59Lg2f
g5/KRk9bRD9h2p5C+HDAkn9EWiYSFDZ56NslwInTEUeHQ7Woo4fuLBKmtITAqyQ9NGT/qOU0sRex
S5oNewxTb6kQvwlkcLyLOlN2kuvpx7UhRA+EID3PMMNcD4NgfIretkT3cWp0rixVvfsHt53cFPR3
sBmw1mVXCCerPKC9axHt2lBMIt3t38CswuAGj0AU4SuGJdBKe1wttwH7V1cOqSoe9Q2or/mZd6Zv
zJvUe3jkFiMr7wf4nPjYDf3jAiFL2v3x8np/xoDxOzQQvvKP+JI8+lBUezZI4eKDewe/Se+8jufb
KdsfPgiqt2Z1x83QaB/YO2BUmGU0c60nQS1CKlm/qZgyzOFyVJRt4YZXuy2ecss+WAwJ80qgjMMA
63fm5ajOFznYxyKyrLIci0jvYzb+UmxtE7oHpkpzGsQjyG8ZjE8PUtGE1JPYx0z6niLDG4nTY+lM
7IGZCDLbsqRaKDyclvcoDL04ZKVgxs1TAXXotSJh/XIUKCdjZ0pEySCxbEVpnJzzs02itFfXK2Oy
oQHU4+AYgwSzq3n2dDQSyRodX5jTLW7KKlpDRZB+qLVXFZoZAw3frYQfD5oRBGPyfVPOJhUxGPA1
UhaVaL3+6Jx/J08+SfvW+zpBYcUeHjHr0NctwU6PbvvkipFsE5MjMwNGT+ML0eooUNPyk98GoUwn
htCGVYSOq3mQGsa5ASPh2RweP3H+uRK/w1ZaD1qPcMct4NCWOnSU45mquuKwXF4cX7rKqfye4b5O
Uvmvc7o2Gfl3LnVW4ThKgdEx4cfMOirYKoyQZPWIv9cnwJ1WM3JtoqoZvdWGbxmDgz2euVBdX3q0
Iul6QfF/Lsctv9Gqh+kb5uCmYJ4a9rzIktsfpVKY9gXKZiimHKoSJrfHZnb9SWsoDnjpouBWdVwJ
vF1JYFTTUL+M8oEEPoduXu/8zyeaD3Gp/AGCf8A2j1UWWJfz/8klRZ4ZZfc1AWqAU/EhWop6bddQ
lqu1P3hLkKXuuL0aV42MOvJ5BSPRZ5kYsFb9j4wLoC659AsWtK7w6Uc8CyqQqMETDXp01ct/MBmK
OfR9fxvppH97GYZXQUL94+jClt7onTRZpxAviV56Umi9A8JiHWGlMyqq+cckhO4XIXuaOLiP72I0
e32uNSkEeyNR0LAJkA21nnTVPktZE57tXevLDyX0bjVqCkgpKgvupQl8mBO/Q8VhTGL6REdmaFjN
CUSjGqV0xjEFn90F/c7BsyLdaQ77rpXT/c0t/yadLnlscAMgZlsn4J0LA2B/8u1otPBQYSevH38c
rDJs7ZN18bC+SAVMjToVpLMXP2zqMGGOaUpUQh33mMCRMZnNaehQpahnYaMy+gGCWOCXLTi3Nk+i
gli1F9ZF7puyHY9JOFISgPCGE6IFgketkLjCq8pNentz0MLfyzb6iZJlhg9Iu6q+hnKjEbKFgVLN
gG6N/43elYj2GwbUulUCrIWBBTRnPZvzP4p9P3A9g+MFutYofbFZksOmPrScUcdO+C56pp7koh99
RDjoVhNiq4ebfNGT51psSJQd4DjCmVe1AW0WHOG0ViQutjmVP2D0Nfomkcw01913bE3E0blwJZ5r
w4/G2/OqXfzn1k1wEZ8JxyVpLnqvSAqZ6OaLyQLzuswAvQOxLfZfEOCpiRh+69qOaODjEgtOiwfr
SihUaDHqaltHfth70dLqA1T5lThBdEoPQuDlgpFTt2UZRsUi8vRz+i+9FFKJduSNxXS/ZMCT7g7U
o7W/9C4kRjP3kTGjdHCWf4rwHidFCJoZfGOJVPq1QH+4FXKeAE+eAmxdbV+oZsvfYmctqIpG38OT
9MRAFrfOuWWWtEu8Ve3rekGf8Ml8XOkjzxZ2mYe/6xm7kL6av0NGLQ73/40rXpm4IVT2HeoFs2wR
BkWOhqpoW5X9oggQiOsSl34utZupSc4QJjvMVoldzUWi6jkEa0mrGZFw0i/1O3U7kIaHbYc4vkuD
pn2MZBzalVzeqOtfQy8IvH5eUEv7EYqMgvkbr8a/xjRZEGB5BA6yvBSmSEPUjJqxoC9zPdbiIW7X
aaMct4cTUvF0egXk0rBwMNafQHNBO7EIPRvCt3ZUeXe6C6csp2xI3qpn1JsXAqNF6us9hKLWBoRb
TjLf3U7hfvAqaffDuPIFCcNa1b0/D1tPfjSo3zH7GCzeFFzeEOBLrnQizsVhw5/goNKl3TDNYlNr
OWWeDHpm5+madh2HykrFn5hU0EubpX+JfQp4eRWOP+ARnr7aRQGl5YW6TFzEARl+wcO3dTp6buYc
35Xjx2tbgbFGSmR0tQAZZel0hbvcyemWyvuqObz/1OquBjvg4g8gotlx+pxm6XgtV77+l/PjCyQf
M2tWHjOnobJmI/9t2fQVXOBQsjWRhoiTPy3ZEaM/UUWbBF4nqw9/JW12hAhrmThHFR5oOxb0Yu8W
8xXsl5y3pfKQu865GcOS/gDUrgQaQaZHdbrYpH3cKrdKb+3AzQ8HdVDtZzSSK8Hr5asSSy7QAYcQ
M/lRvM0JTsCQamjyhurp1dClbI5RAF9OyJs6BrVgIhtASxoWrRiQmtj1EOwWj1jMjGm+IkdBZ/1L
lLtgh/NWBufJatYC9uHtWEBF7sullJLe+/pCsT7QWB08V6QZtHvvr/J9ceGgwD7GjsU3mlCrANiz
ky8lMbG/b4vI3RFzX7qg5B2pUTI0Qlo2xRoGCc7BxlgIUsUP+2r/lv3k585A71+MS9V6A6OnvqQB
kkdWzJQZkCIsPwcFKIVhmVYlMqlIR5PkJ6sZwILsKqvc7j1cBddOH2b0LVlqGyHwq8m1n+yarrir
SZG4IOiGDLU37sRZo2d4Yjc7hiLyAUau4MkIStj6I7R4rlzo9HFacipOyHo2Rdxmt/O3Nsfoa/49
eCfK6mtq6coQbiSnLklM5Sq472gPVhIXnhNPUN5Vaku7rmHAZRGBC532jaY4xdQdKoKaGnYQjOgx
SDzOLbkRr4Art8BuQgvy8/6EBAV95qgh+5hcvSJISv7RNne2JLSfg4ld9wjgEqKmCVi69tSjdXaB
ALmcZhh0zUsPkr/y3SnF8RbI2lb+xYOdBkpURfALMej+pYwidsbUe6ueF4IXsem/ri6p8qJdrWUD
KxVrZDwp+BcTtHXEK1opHb6oI7bKaTIqhIVW3MdevqIHpFCdWbLXK63xO4cC2VD22pWHxONc1xmD
7og6yyc0i04TB/WgEcdDqFimVVy709Mt7coAFmcisq8WpvRycBmUG3Hnhy5rYKdxpLWu1fqipoh/
HwBPqJ29vL8DDXBevI5pCKodUIx8Gul50LlyEuYX/IGFCeHVwjviRj+GstkPD9w7IzP/LzSGgV89
9bD9TszDpsqSJKfP9xC+9QmKqiFJnM8rRYO7jqWNpbxcEB7C1VA5T7Cc/cV0wG2Vsc727aYTTpQJ
ddjqMESzpfncQ7v5sxyGW3TW7iC4Ebc99McuGjqTTWcsYiZxYL+yVX9pOjtXCtPJlBjAqPup01Mw
ob+lD1pQM8xgSiKE6bDXqIRA8cx7Jx5w6e8D2xOCUmtoICmZf8ZGiVMNPHdaEZXsmddds8hH1V2V
x+919trTsiKUEQ/BiRVvlomjltaHrJTGd0gd655jsAHU66B2OUMKqYbSEThTtozkFiDJrhAsd5o9
wZmB7s16G8tin7+O7wWPxYSirVppmmlbuZqmk8ISQT7oc8E0a06RZF63tdYpuphjVKxRitY+raBP
8fmHdwVBExA+yTOO2DshDLKeWEj9OV23pC4FBKvPhaYyQoU6VfGwhWuPQ/7gLVi2S3vmE+wNPV0L
/sNzHBmSqUXmsXryU0pzfzkj4TROZfeheZJvN6u8F/fOQfxtkkQTaeSiWfybjv7N+R2B7M6QxiTy
+RkdgZm5d/Abc3xppIIw9d44Y3noVRdNNDk1J74Yw6VLAb5OjDHZB7FtKLfCxYY29Cfh848abBtr
QIU0/0CoaWsF9nzvaenmHbpEBh4Ix3Z3SRNutu4cnSi1kce7jjAJELhV5Vw4ED4jje6G4zDiYtHN
8x2kpGsXUyYOtvx9/EWWAKt0SKJJ0OJ5Np4Y0pJ+lAxiCq1zm/GUr9ECCfGezf8VrogdSbvKghq6
ZWZ765qDd8btKowdPJ1h1K8S82wQ/ih3e0uIa9nROWN2kWEyKqyYrvrum76DJ3TlUKDjeIrzpDJU
FDgcTcMRWvFK0YJNzZRTHQTM+h3kZ7y+AgyVsshR3i8gHMwMq/3jos+uysLY2uParNlgoIhiEgJT
2MCHEFFoAn1Ijg1iQhhWWE++PJc05e8MYgBJym1Dzp5d3ex3JwlvHlZP1zwof0TVr+Y83r58CkIp
un808HImI5KN8OWiDp8BxiOu6s04SvOWRF8Z+Tn04YjqJFUPC2o+lwf1gY+FghzJMKsi0r9zDVa+
OhrBw8ORcKXfdbgbmPo0QETWjuoFkKeubsGuee2t5YG/cN5U78mUBpjv2v0HxysvB6jGcDzD2BzW
3w/klLqveH1xaE4GMikPjOViWP/BNudhEtIPkcIF5hndLIAYUWjUxCXjQHcRtFNhkjgeobueAUQm
9bzmV3nFI5PVI5pEywTnb+WVPQ15VbEzJguD+6wnraa+9d0n4fqXii+RNJMRpG12Imlbyer/LE8w
DN8RxSqLilMAdZ8NMhrqgBv1t4lT/2O9sk75p243zaD4hCwcfehAAwSFNY7LlKa2IzGHaGJd94hc
JE7sa8duSQ8ZHMuAGBYufA1FEEPjb9p8AY7Gr1CFMjpTYk7NXF90GQ/R9Pd4CweuHw3p6hGXhjw5
dHrY8pEzuuGqtnD25o8556l/fJVsH/OxLSQD5gMLnlTjXAd9LoKDKCnb9iSRQEgJhIvXOe7UDONA
FgJwC8wiihal2tb5acr5JbKX4BvAJSP9V/lGl5dKQpbKa+a6r+V6F7ScFGercaqNAuvOsWkNlbEH
H4aVC8jq02A/SVhevGwFBQl9iBGrHACqkTgPtYp7dYSRj4EzBduTQS4GzoLwvslPxJN9HxLoT6BD
uxVYcn9cFuk3fzhYsK46KwQqtg9lebEOJ92tfI4VEExrrdHYh92bY4GogZK1CG2vDasqyhqU1y6m
NeNKMA2Al+CmIVjhuAXGX/D0kBch7xPD1mxnPHErzpdogS7ZAdC7N891zILvZdrlE3sKmrN3SegM
LWnHoKLlo+bVk7Yh7skEMLbQs8ZyAW07YJywueE3nmLJmbXB8h7xar8nnF1YZo2FMkxjwd3J3jyi
L7OMUvHpPH+QElZUTyY6VY7hRhjUXOqA6aAneLsljAh54sokaIjGNprrU12N0wvSL3qpczzmkMMz
RDMzlxK7xzKHWgT96JCskGMdsAdYfbG4gg1MeeEnTrEP3YDndTd7o7ODDHKISTkivVXrkrrFv/eq
oJIkMrmLAZoyDBwqL/mIu5hxPDuvLDLXsRSsKaiR/B4q2YUUAvl8XPXKPWby6rPCNYupKQWvUcpA
qoxaXvQ+sNjeYPJaIthKCmdIGZdzgYne7zA9MxQojVCs4dnM1FqDs7hwzMMHHNsMg+39RTNPc44j
R+sR0rVO9cNsjRfMtAfsZjz8hbWdZHzE2GkX9aTZWx6lHIoSx7cryMXsEDtpnEvTpM6fh851QRsW
RqeYw8wWqBsXzNU2RirTXcRIlpf1rJ6vqwNDAtbJu8KdYqRfphJ4eci47sqXSz2d8GmZVW3NcOdU
SIJWsOwdrJkT0QHC92E4arFBvL/h6Q4SsLt0J6Ka+n8gXG+DaLz5rY0MS08KArr/QXFODFknNyLx
iwfuHXdJY23xIOdCR1QO0jxMUChObV9bxSqy/VomeKzim23nPtZGHN2Oc6QXgRYXWI22l2vjT++a
h5jjBf5j/C4CSRZb0YekuWWY4b1FMPSTT6eUEy5xD9PnjRr3rQtrDJ8ivIqcADPxJ2DqesYJY4yX
mErjvWHqyGbvYIZ6LcwhyDJIC2atcVuA2XNxCnW6p0lpXCfdren7afuCe7SAJ7pcovIuGkNEYsWN
Jobuv02mxQJMBqF9jak7PG0ij6/p8vSupt2Gt+YlK4NySuZTYaAIfwZ2blOqx+qCQzs94E4KJofS
9+zT+PyzxRS6exYhRKBTs+f6bdWK32RGjetDsofm6cK22u2KC/hGFcPqBJ3TUDCG35AfDSgr/9K2
NDaNWonhY6Bj8L7Zk7GwXa9qL0k7NVdWprcQsfl730KR5DI0dolMvv8UsMp5/kMV155taCdC7OwK
oL5fQaKCoCasf/hD6NQP6Y3fl4DDNcsOFScFZDnlnibdvPO3tyHU8mrImy2Ypl73r8PxtTDySVuK
GnfLKpQl5yGwyICiTbsh4JaDuVZM6t/hSGUq812GSrrFxO1V5cU13rZm7TpF+FuAzuBW4bKt8H25
u6JJkOJ612gyJeiNVLi2iyQFqRScJ5GGkxKFNI1Y8SR3cMwEWa7yiHA+/qBreSZh36gFaJbPufMt
1L5MTN4947cln6UzBIYQrvOEy1FKWun4uG9zNenpp7GDI/iPaCK0z4Il2186DmA5d8JW9nGihKML
dkzXjAaaFhUTtRhYps9c6ZFkFlpgZj0i4RH+bSCSpJTSok871GdJcmkO+sgc2QMiMS+Y3JV3spNn
NrMkIFu4m4q3ain9+q+xp93ZcqSWSuR0fuyhRmrYCfEdnOf76rreyukoVDbfMqzdm7XNb5xNfIEA
8WO01NSxQbx1532bH26HdFsPuCla2IuGqEi/X6I+2QqQI4fz3oAvxDanLI/yJLXngSOP1EMyYxLA
EywH0+dH1+jlarFY7KBcVxC37P59C4Sg+u02rwuCyr/DN8131irfZsF/hBcj/iHEX9soHsxTT7EQ
XehmkfhRouGbaT3RcwbkF15pgP4Vpj/UDuKFcHy/NEzYQNBfXvRomgWwMRdQ2vD3Onu9KrFxwDUY
qho3F4SCotO+eL5LPer6dbM1ytQ6zw9coCXCgp85dkaufaQixW80/dedtAw8tjC7qB/vW4zDooDS
KwJayB9mHwZVe4k3KZ/1EBgZEPpUDq3giJ5n75/82RV0afKalNGW+PXhJ9w7pYrMSSWVgvtN1OuC
6/+MVjUsh2LUWQsRYfVCk1AeoTUP9hilL+iM5fWqKIMXBYPR1hJQ9thUtkFzHoPstcjZsYXaKXxo
BdsEvb+IdYfQSseQC1wNEWkAFBYr8fs9hPhlsNqrfLLFfI+eStvY4cbtQkXY/gAMmOILMvaIyldG
hJOSgswjhfa+EoiRLVQ4JibHLOFYPq/Ia7Xy3BDZp3WHAoq6FfZ0GgKaDK+2J8BAtvJHpsUX6K/5
dlBUErr2m1+kT0S3nNJVFT2RW26WsaVHkmhQUHxtSeDc0r06HttLztefdwpa9r/vzUtf+widrzOc
UxOqgzsWLOAO8gEOpG1cJS9j7+o8f2IQzvEXj80ZzJbVu0raE3AKcAjr65Q9i2MLegFb/GmKIG+u
xo/B5YJUQW42wLtC8o2l6gOfIZKL0+vzbMXdXevmft2ImXAtc2yrcujC2AYTl+cctuHer0WwP/hQ
IQnTgW0AeJOEwcpfJir1KV8fzTM4OmVWm7c3VHTcM1y7JDQxHWYCpYLbOkIIs4jG1KusrQIW8DIG
ForXjDY1FAnATCU0w76funt9wiLY6kPERbGRaS1FluxmGVKpeoCSFl3G4Uzq9++F7r+EhiUGmrIk
iULgHSxHuhnKE59EQIrSN1xFTB7X5fJr1jaXEsW7rLt+jlNybu3JH8tr1siZfVkjyz7FRVrQwDI/
7bvX1IHkmTZidmYLk6LDC/KHMCLwy66E8wV/Oz4cSGCi9dMuMjvncg8rc/l41Wy07Yuc90Z7pHEx
RWwCeDPRfQ4ZjnzYX3sgFaPS4qG/UV2N4adJFShUNGcdeKBBOcJoPQOx7rjtFXH/esTjIpWQQfVk
1Uq2CoL2WU9F6jLF166+ybl46S70clRODJ8iO7B8SwUiyAkVPIBLESsGHE/p9m7Mp3njdPcRO4kW
jvl0LR+4szRBEsZvc2fEU7wBv1vC3KbIetI5o34r/i6jTa3Me7LX+14RoDygJ7wnBtUYWSji+qjN
GKJsBg2wIOf67DY+y2Sv4N832layij2O634IuO4THa8TOO5zwJKrHv/KeTbQCaqVCSt+DfLaxLr5
NEjaJowcEepex1pXZY73/1raTs02DhIU2A+vkrMMYcoKC5Nct6rAVhcEZYyJgAYkzd8cjAlqTBRq
OO/aRdOs10fdkm/tj9Y+f9xHYqt+CqKYcNk4puRt+ClCEbE4DPrcRIXVc/4ZhlDBkOE6cydlPlRo
rWOmbqVVTqezr55jW6lFcye07+ltKdKE1z/I5YP6y0cytZa3BcJwXu5qYH+iOBomm4nPE7HGYPJQ
Iv+h40EnU/mEDuFcfxb4WStDzBDf5TnDV4ol9gnDh/TG8lmdbAzGkiRCrWG9qGq0/fQsB1Kug2/q
NZjNdNxuP1QGGXjVEFGeSRJoywVzb7Filst4ohXTGVQWqtOfTvWwzyfiuzJ2Xfcis0+ESzPmwRa9
zCQD/Gm6kXIrZW2s0JhLqwNqsULjwkjcUGNENwjZvryQgSChvUp8Rl7Jx5w4qvEmlPekOLdU9ofV
/wkyO6sjEptBQlfk1aBoDbNpak6kv5xFrN/jL+t+WN20v2ZXxbfIIHxsK+b96hKd7vCi3XzKtQQb
w0W435jqm1vpisBwNnate/if6QWkwy8aHcNmxNCV+9ndTAs4z57X87msnPN6BoVd6zskhdMt1Pfv
NTjK7vRP+vvV/fDBifhY/EgrVYvXQ6Rt5XvGEwXKkWicunm47qQDqhCHGl96gnxvAojfGzUPBCUF
F/WUMRwEraR+LzPMqr83JG6Bsao7+GVTiEWAvnHKOjOfu9UmDjD59qLT5SiTIozk/9prOX1mxRxH
A23Gk0EejEEhyQCUOUqCjg24bowhK2VGpc9KvnGyE3LyoE1PeJWA2IP2V2TurkNPwuRZeuW/IK9B
rnSW3/ZLIJEups8Wg96tCuOlgHU2J3bQ3fQH6vFVLtsQvCTLv3m31oSDmm1pNDqJVmyXTfZRB/r8
LTVoveEUIV2BwAR9/jxabz71imSY6Xwllbp/26j+tApKLsF1I3/W1pjqdBNrgkEvmyLCkoO0F452
69y1KUZhw62/VIg8Fxv7ixI8+66ej+YxvLNUUbBKOjQkAdX9R76X4UTKgmoxCPFq7W0azQE5eJ8u
5fmo9PHgcvxg4LHEGCkf3u/CKy3NaYCfmIys1FCFgnnsTP6KQJadxGbhjKfee4YKoTQjrgdDQhXk
68nvTMsDKJvwMn2TfZ5GgrzAai+YwFL5dlMzYT2idY4xiO5OYFViNrqO2onC4ltMUOTzsZqUeOCx
Qe998IKTxXXFm/nsdoeD29bMq9mMbFTdP4m1UNDu2MTRBxrbm63QCD7Z1rxubjj8ddqeI+VgZvSM
puXiAIRgwT9WAeDGl96sTOv4loMhSIoRcErLLzz7bVGX07mOi/t9kyGmWwpcRX/ZxSjfRhmCO5RO
SzJWMR0jKETq9hfEBVY/X6m9jrSvl8wT4hcAY1IigDXelBZZNJLSwBgvDJn7i8NxttmIEqK92lf8
jRsR61uwlZIkpZkzebpQwpm7wGC7Q3S8DCduE27Ot59I4+nyh6RoDoOpSngnYnKRvRwdK1Px0Swt
j+tOW6EcF1ph5a6imvWXdCId8y2HhPV/j1mmDj/sN0pGAvJK3dJhi/6FDeMJjPgd+OH6jd07q5cN
PVrudp9lecOBeiFohh6qn65HH5aaf8wa8fom2vEJhKq30nBOGk/w3OcdpqL7B2IaLxmYC/cPe3UW
K5fFOBosHP9HWHm5pyyiJ8HiTQTe5wsmNUJen5tWJN+6tbG5lY8DtWKzVLgmbgBoh8+T5ErssM/Q
3pb9Sg63O4dDOXoRyR1TALkiPISM92o80ey+EVbHRStbFbNVG/LnRcfYpEtGrE5ubgsVO0qwpUJL
NLuF65VAa3RgwvSERQ6kiXQpdt0Lq0v4V08aqCzG/jwcabiMLCt3EykXQMhTCnyUQVkeaCJCGU9R
p7ZaTNhrUtk213UeepKnYYx1sEzUCWz1ZnEeiXFmZKjtgsz+06mgEnohK0Zj/Y8bZ2eTny7Ci3RN
B5wVLcww+EoUKk18LEg1u//KPQi8+U7fZ4fnIlkzve5vFlG+aH/FQaBWQfkFDptB/Yfc5W6qgEKI
EzH1Utx8MFkRHOiIw4A+lAUo+GMvdAekQRN3YZ6kpS0N2iWGCQAKeKS/P5WlxhNWulVfBc5eFN5A
zdGizvNk6LYc7Be2z3ykUKhB8rKlvX3Qy4OibkXjV/iQ7m94yonY/61LCOQhvPCOm1/Z57yw+2dY
5K6p6I5cZGMiztBo59ecocgoPr7vkIzPe6YFAOxkc3JDUZSvh17Rwrz/Lmhse4YvaatqDTJvZzAS
spzWdiy3IAR6Z6eXvJfbu0y7RIYJ2FLzhHEYSOk7JBVr7VNFJIDrnJ9mQ5VXbD7R3kCXFsxUdgxE
F4sPYVtd4xkqOOOISqBsv7o7r4TLgteLH85GawvgrGp7WTJpwqy7e2BFCtqRKKcwZ+3gbZyVjDaE
QemuS0gmk6XhkeWTFp5a+K7bojaMaGi+g6rDrnJ6hsncg3GOCtc2IIr9/Z90J5ASSYeI2gmxZYxJ
leJM6Br9abVQ1LIGIpwpdK+1JhzbM6e48cvF5SIpv2qqv0EWvaDFr4qGsLiioFYAwmwqhsSmSPhc
OLkxVNjvkv5wr1rWZgfIcVvFVFnisGsecataNqH3dgrS1CgO5m8dHdpQbU12RzwQEvFVoL1AmnrF
LnhT5Ho2b3OewR29cHj6Heos14h5ND+oc4iUJiyQoR2iX2xEmRhxSSYZ+BK2TCheHSYpLQAsOdZS
BM8yS/ZrpwUt6QjST5AgjmH42AYQvz4iHdOI4KuY8Uh9p9qved/m8HQo7Ki7RWj2xx2cdQ6o6eL7
yhWpcV6uPoaOkrf/c4BRePm46+KMDWoyDg/mA5ogVmxl+v3qDWxyDbTqXTihathpkaYGBB07Nq6N
gq9Mm90eODkQjZAJO3WGaR7Im5tS+fI1VczWlWIq3TO1+ZVwyZGNrlXy2kqfwcmkqzAm+BaRdGpU
+JhE5mAjgHw6fyUpewQSTdgMPXzcPZet5UncR1q3gff/OpigPVygY8eW7qIWnRhHbYWrnuB31z1R
/2DyDFTpbOPdqfm/XrjGfRm2u0PzprMLRgaHhwzPUhrMHUDDc0uMWMd1Qm8bo0+8ffqtCzVvDU4Q
mRa3/VoNIS1w8UBruXUlCpDiLDlennxEC780HmyV74yNrPiEEXlqGoiDaRDiomzW9WMM+ILoix8r
7PVNrNeHPkvU+VfENAEqEdYwCfK09s5oLESRn9ZTz37jEWCxrPYMSexQjqvcrTKmC6j7yxi4gc1u
jciVqnN8hif4NK62C3zjKP84yHvvtL0qjE0oMFVbUekt5Czs/WMUlyg4x0PX7G7CxPvs3F9rVWqF
Y0D8mp7p15pNGOu/0N7O3AN039SAMvVWjiFjUG/1aBHL5CkEQWnbfbGhz6JRO2JPCyoaOpMS0Ic5
S2a0T9ApUAZYCCgx5h9xckmtm2Qti03/YRFZX/wUfyNTDGFKmuOMOrlXDI6uPiVB1McS73IKiYgb
D8kG6XJSsufikQTUQh3o5rJ/VsO3ACkpH9TVciycFYcPZoTBFKggQhGtPkE8fEEJ5aB3kUSyNbxO
ZKaj1mIisejd38XF9ZUz8NfcdTX2EYDKypujT3G3MMmlxZXwsOpkkFJeuFba7SPEH+F0iJxItnFT
jEy33OY+ztpE39Cgkon0cNv536OLAtrr6I5hvuRrk7Wqyq0TguQOnKBWJxK4/NWRrlZVhZqVgwwb
gjdFUoQOmvLEEquorZBx0lZz1N0pN8rqeRoqlZIU95oDfiUcfSIRG6po7FtL5GksNhUjFM/Yh7xR
/2b2A69IyHSPUFMRcT/NQcihlLh1S/PO9PGlBTQbCpOsGHdaoq3xkX35bS0Tsg/cf73HDkDX2qaa
QAgGPwZQwBDuy4nJXHzzf7Wy7TJ8eQ79IX9QoWNXCIRsyuGK26DCGa8ui9gFf5otgFaZXiZFvouh
3vdG+EwkqG330WKWTzMGMD5gZiELQTWwBurHOVXphFjmi6UN6l6rQbMqdOmku/BHDoq244P758S7
mBZ5UsJ8yqV800HwJsZemyoRYpU8ySc55rxXA+JDXJmrswctvNBaOWbOKpN62lTKphqofPpHwzUS
xqohDLQB4qbzMAOzsQ/StA7jeMTUNX2aMuBEq9fwWPbQCV12U+e0oDtUNLxtO8aAHrncUhEgtSAo
UH1WQAJwqJCjyFDMF7VQD2OnBTSN9j2j8aCuN+6gmxL+jzhqUjA/eJQ3YrbzrwOa8u5VReGKZiaj
Yic2wpfEtA/BFWYMqSbFeMnsTX8X+W7w2G0Q2fXsRCQrHH8MUuSn0KxkVryJw7Cf+KgN3WjBYVKH
H322cwy2347oA2WMpR0vtuhi4OUGjLOjYBlsF1Hl6m78GJPCll7poUF6sMAmFV4/St2pcIkJ/SBO
WVXRwhyOiKojziKJZMcqFfMSI4I11VRgneiJbMGPAyfyHFbKjAhBYXaQ7InvM6svj3UPgD835wJs
4V+llw9j/Ty76HfgLBpjLS1vrP1mNcZ4YBc4NB+kox81NH3P0ZPv/Qq6P2P3YrnBZq8U7SXyROD9
KZkI0jDNJUi6A96c0XkKzu9lHrQ88D4G5wF/MU5A+E7GsqiYy/Mb1UG+MFkTx+QojfurcK6O4tEs
o/SLjbfUvHv9r99m+pPfaw8F46ZOsWzwFGDAea5KJgmP+O1zFF7tNGlrMceHqskriOntBQjx1oFt
JaVPFaMLXNCKdqCzDcK4hsWa7zBlzutpqCeCdhKPhN6NrG+MIfVTxrehnTQ9j5SVSMH6pTJt7An0
IN9OWES3kkFO0WpIkoUUfQBtUqcnZpp9KaetARl0dxzJ76nd1xFTBMyYQxLF7oItKCb7bL2QSeiv
sNGREYU1dcS0/u9oXL/d8BJEXgBnuGgFAPD0SQufczSBCzQoeTf4YZMBTZYb10yHKmiamujurIRw
PCI9O35gwXYDXUZktuCJZNecUVdykjWNoxdCbL0IypbLiczR8+Ttb/PrsxUoWs1AFb0tp3fdY2nE
12fuWQ96ls35HxL9mr05K77ywqX3RKWXaZ/vLbsVwtmgP2g6sbDs0D9mceQdoa/HgKdGWeSSxAYc
J75+nqwAdN57to6YAaiH6fCiygXiFOXa2ATfjzLQYYk6uXSRpuAOfC1xACMJvDitAi6l1YyMS898
nQSWAsVo/mhYU/TvEIuifoPZRtOebtPf4vi8rHV7sIW71JI+WF+RdeLkV9Ro0PQj6GFVdgh5a03s
vQ5bKCAFnvDUPDW4hmvUl1lu7FLUsndmDIOlQ4mr+SHjx/Lipa3blIh+RoGvOUKpHz4PvPKHx+cT
7R31oQHgJMQoe9IKvhw6yKSNIkKMTbm+IJ/x4dj1RR/XEorgTs6XRnwbfPT14efGkQYQ/6F0T5Gg
14Uc5KDjzJfZHY6D9Ye/7NLUzboQ3If6tUHTxm4VdvPisTxFQ3yN8zrHFkr/38pin3cYL5KVmME1
wpYE7aqKq+W8vyn9gTmjZp8ZTMwVN0xKYs3ZPioV4IUCCmxs+bzB0+0dk1u9kf31dbYArjGIoMa3
zJ9a/biOaQp/+winLJ6H/r1+yDHPp8U/zrv2MQlVqrQRyOOKLFgQjNtH6fbklzJwGOgWE/vtvKQ5
6/h6+yZhpJOT6dVG9Op2x/A57Ut7cUR/bNDzIC4VYGlwrmUfcOU+zaEdJyccxoLi/6ld2vYEjK7K
YpOJlWj0daSlKQj+pDoLqXAtK2GzDMbbbDPAgY7Rw+1fLQ/dcRxE88T2ve9X52LgvrHHKjXH1Nve
A5teaTWiZ6eK5qQMvKx5FcHI1b/RIMcYoLR/0fqUjlFBhGoXTYMHOs3qdGRj21QEErZ5oTDLI45M
cshV5DNiah9QhY+U+X2lSGiAQ4s/5VBMgPdxtj+Yplq5VtbDKlf8agkYq5EtVBkuMeKfbWNXRajZ
9V796GTyxb7z1klS8HVMaZ+t9thynlutlrVuweY7g+63tGzAsrxkT58OM2Qf7NOH4wIRHjVho1g4
IAtYEblcOcsCJNjd9jQhtaq3kA7yOgve6x5bKW7BW8HSaLls6LXB6j3mA9dTL6woxY/3FEDcqxwj
4NxlewE8A0Ya9SW2q7fAdCFC4suUGI7Q8ka8o0JgiDqm/2teMbPJNCNpH74PSP7CTwi3C4Kqjk3u
rXaDfZeluJIGpfk59f664JNlPKE0LpUSIhRt8lfcz1KRzVyStKAVd8Bc2C2Nc9wSvRJqKMQStwxk
SDSFEIOXGQta6K7XI3zhWaHNsrsiiXByLht5qB/5rqAn1CN2fwqde6ei6Fo7HzXQYSWi+H4lI81B
LvcV8to3KQM/eOKC17xduJ9hzOlUyqmD4XnaJeUFkPF3arKUBFoiBMT4SU6K5H8gxh4b1BLxEf4a
94jf5iRdAKPiQLWJFjfJOM/JraxieMJN5eTui/baBL6Y0vJksv1iXM92jCKW0T+eO/qfa3Vc1dDo
hpE8GQ2ycg/GBPhm6fTmsf37rxYDry4GIJo894BEepV11ZBV9mO2OEbtkOjSvr/QRUjn5Lego5hI
4Gw/bpLvX2OpBx+EHqDppe1TZeaac4fzB6sYWBseufYGifaV5Ur8jSIomFouFwaqBRtCtiWXDYwk
lyi/QOJKKnLdYsJsw/i3dNClSrYln3kH3Wg/yrrjRRWZgQpJIj+9vsF1cBK27lD+4FsVTNHDJVFi
P2ZdpScUwDhq0kTEJXwWVoMc2TcMOWVNhLXgf5yPfGUGxDYNPGtliDmMCfcfkkRPduaeThpZG/06
uyFiwjAqlojWYajM4YxrkPS9DBNrjEytjlhR3Xs/gsr+vx1AouFa5aMV3vS4FQFfjIZHMuWTm277
nERezkf2GyU9h31nyBnrUE1u6tWSShSJBZhmSEfBMgxg+zBfPwQWvlc9O98Ozqi+cdN7yGjuDMZ2
NVcg78e9pEXKGS45EEBr8Jp8wKLJXkpxV82SwhuE3AmkJgceo7slQp7/aQfRCVeIj95W/e8fwloR
beul6skgGp5mp3QWnYYpM9LyNNwy+kt8xvvp9Peg7oMRktGwmZwl5ZZdPL73+FnhQQCAslRVV2Ng
ZGKo41KShdhI4US+ZHSqGqu1DAqB7mw8PhMVk32fzILlzOtph38u304Hyc2GcaPhTvX/phh2H/Dq
EwBCJH5pPmhvmucgPxvDsighOQnMKcDXuU0J4uq/SjO0SG2+TV4ba+RyVigdUgJJTCxPgEQOD+3w
Y/f+o99iI9pWRO+vlFYaWl4qh8ovgyleJLlLNnXLGpoiE64CevJrLb1UujJYZLrDg8Wu7jRDX3SU
9lN19ttna2fV0Q1z03y/YnM19vpj9P+79auSDD67DuoG50liPfrbq7+YgoCTiSJdwBZ+QaW5mAF6
J2fytJ+stGdk8XNIRwa6a18FMm0id9Dpcy7HnbtA3r4h9AtdZ3uDXlJSt72bsR44qaWgEclXW0rk
5zBLrtInCwjWVmAAoFrqR1f+MlOuY+jVUoO/neohvjOdFTYTE+f7E32h31wV0VnSzGCG7AsyQxkg
+YPbIjZqhaDdz3yCGRQxiWM5HCNeSoWwMG9tkCMivyq5cW01ox/OOqeYj1YfFzQFlN/CTCAHyI+9
tmSj3ArQ0rT0Xu9PV5Ks/KwXPP8eBsa0sRmvYSNc4tpJjxArULk5/FauSzU+JolkJHriKYLZVHJF
PsRtSGttrrfYg6doXeGm7KS1/dkLB+zBsT/6Q0kInlb0uJioGADoCUF/+aFCVm+cP6eMhgS9iJh5
amPSGwRwLzQGD19eUuB4qyHLhkv6ahAjy7ENCa60ZXoLVln282LAcJaxgUNxUpB1Oug16uPbXHiN
PeBAVd4WKXWAMiKDeIMi1+3/FpQKOwZXFm6lM1f6Hn5ymNyhESqGscqDJcBfatCbRnOWhDgfASj6
L/YjsLxhWdf89yCcV6Z7v+qPPKGxYhvcYXXFHBfFC4yeLPHTvYGc83NgvBuR3iUJig8d1sgKmskv
Bl9yt1TWU4Bd9R5xXwX74ImIvkwZvBMNTxGDiq2vnGLumEs/nPVLuAeTjh4pQZdsP92YHQIl1VsN
rY0U+vJwLviBOZnwZQEtBmoZ7RMwygOxKDAOHSjvZQ4pMMB/WFE5fgImQCL1u+ZI3WqHZGJn49eW
BYCk0xlYUMbU2XiQJbxoNCbmzKc1wUoQPCVfcjzx36K8zaf6Tzmgwt/8h7I0bsxo5xQ24Al5hMu3
vno3zpg1TRAYsx6kg8k0kXJASLUlnapLvPcwhuUPvugEQYSP5YTzk4eCMwT0fWia++wi/oCapOFm
8b1WFdWSNRd1qesP31Rf9Y37nY/J8k/hJULLSXVO5uWsYJ6wV/N8YlhtXpWNLVhq8TYsaMoAHEld
aNKOJ45priku7GEU7p37khQd1TJLEZ76pmClQXqTPtMJgf0teajx26y1/1SivLZ61azMEtLt6j/a
JFZq4wTtslDzd1p/eK8XE6y4pWE58JJkukfJwLE+eHl2Gwu7675Di6DcyLTzSkApCK5u6ELQKL3z
wOoCS9Hk/hhtxxIoMcluTfKxkZQoEFp9GXz4rDxlX5UIQKpJItTiOvkAASnT2GN0rZ8nAZVbL7yP
yuoqgTO/Pi7GFkylqpXkIM0UxEN9yrql3+JBp5UDkQS1NJvWMq4o+FiMLGyK2IFYZcEUWDAbNjy8
qaEZrMN9/qB8eqVtMdB7oZzwQpAxSf6FVA1RFZZYBfTmCIef0BhuRHf90jRF0LGyFarFxhAab20v
AGNqNqJeXVyAfUVkxN+cs0uSO+W+5qDv4ruvkTZtKmnV112tbP+PZyK/SuWGXpXBwWDxpw5irvzP
WcQozaa9Pu8LwzFk1jhDsyaKOidIac0dQdrH+gY+D1L4zedxgWpC3Z9LKPmrW1E0z+834jyynK9J
ShHnx/BunCdtHm+2dd8zP296nF7ofd/Ymdm9k7aDJtXAPf36s+2J1hOyJi1HccMye9yHqFW9QN4M
WS+6CTsRYa1dm93R7l8S7fQKH9fEY7pRvoy9i38dMzux7gUjVX5uCHQnpDtEvnTzTw6loXzkTQh3
It76ZtxtSGEnNN2+2ghgBw1uPugdkNiVS9G58TOJ5uOc9TnbduNOGlk+gvEfVDEwDAemRN4CrRD1
+cjmUqgIxO7Ewax3b/gldZPnMZTci+4rGrVe5UMRk06iv/WS5wGeUMbNHrbRCj3KT4MYFftMAuKE
RxkBv10Lf1X4d25v7K8GlYZ6tXvtnmJlz4OzhNBpYClgS8BUyTE0Fgmg41VnqWMt1ze2F5TvbeA0
xCIxxMoaUWMtD8SszGagbjajMcjrxeGPi3PXmjT+Y/iQAL1TIDuPXDcNHBz77bxo/ED6qCkwPIhL
c3whHU4EUkwqsePxv2ZSMBQOfEs598OCkcge997sFz457GKfvKCh5La+4do9rsb3xI03IBM5XMJa
i/yugt48ZEPqV55z953wNiasl0DlqUJJ2qxuSnpv7XPxC8WEpE86jbfzRxVvweFP7BBHQDFYf0b2
6Z8nT3f30ksJk5g7y92GQPLnLB54haTzVo+fQ5SrhlGTgiUv+kvhu1ZBAp9N1RCqHN6+QU64WOD0
N19rIzZKaA8A1PkfhxM0le2G3tCSJXSpYU/gMeooUyAwwtDP5uRfNGSFK5O1H5ZaZtZyXxkzrBFi
qB1XhPXHLYqv3o3eq+6Vtww86I9psRPBbfQom/K7pyf6ZQBKXB0bqUuDdBLoa0nk5owFDLNVXbUA
tzF07vIaCIPpM+Z6KCxpaAWla4iwSF1O1x6QjUw+6gE18/+ik2rT/L/oi91HWAd9f4z4bI6elU8g
DnGCI25pdQZSuiZkNk23YMRWza54rZBidT0Rn4dcuICHfu0VuOkXujf4qGcHbF5Q4GSn8MxNKunV
K2HxXaUGxGbiSbrLR3GVcF+G8UzhWt43prbvr0HDbkkCjne+UK5OIinU1a4SA+hm2xEYX/V07fJu
CMxlLTvCIEQYgzgqUwQtzO3V644RXJx6E7Z5V695cZMPzuhzbVof1wjQv+62RMzjm102CC5ytWmd
9sTkKna7uaJzF1mAC++2p2mpI8hg0vWr/aBy9Q16vCGJQAcyHkHd1VLHErmXNTA2LMSQJyJePpOy
T1nwD1mWaGvoDASJliiiOKK1aiKrVtjOIl9JN5pOCXMzzWOEnWMi6DkZ5VBqqyxUo6Va4tgHms1Q
0KG8u3gR+5Bz9N6s6dbNffDPDDDB29vO4PxR6Xvu439Ty3e9ZzG5LoYi34zxFvBAvyiRxIQ2qeR/
3wefPAfzssKlEsJctLzs3UmaYIsrvJ08P4wo6YNcCUn/gCoHM39qGabujQByVMTubZOF/WSC8gtg
vMU30YtQzy30IkAOL+ej/tyJK3JPxUynoRG8rhqDjr2IDNzXWYhSe5Do13u5TAh/GKd9irQAXvMF
nBCLQeZw+ADUgrjLHPxUQCa53ZoE6Ru7Ypx473yKE6gaCn85oZHGoZK+iuHGB/f8TxVJO+IcdRjP
bSxJX+HSg6DLAfZLpVlgE4LI71Kd5eFRXHmA7RcX9q2LJg9GZ8N5Uj+28vG6vJfl/GZHmzaLhhNh
cHCwhHvgZHUU8iPxDo/ydhO/VgLMqq4EN/oyRURhcZNJAvkNdN2GYXMlPxpOFgABsLz0HyO4Uz2r
WhebRjqUqHppvfFhlAoYO2yn4YKr/nCl0H02bof3bW29WfHdJv0djhSeSp5EVwui5SbFqEPnn1ex
V2gFTy2794X6t0tJ13QYyrMM+RRLPJu6CBuIrDx+OijhMQi1pesHgfTKtmtnly0SBISMJDZ1F3WZ
BtxJPrHRFyh3+MSf9zyx+Ij8BgFz5NgvWDvrC9QQ3PIg1PofyxL5zNe7pCO4Xv7bZhlzy7ZstlSZ
mVlMZ22VPNvzVd1DmpL2IQKPU4JLnuZ5O1Hi/38pjTV65rKwjbxXjfFO5wHf12T4IboyZMaOVgLl
5Ck4CQNH0u6OPDntEfMHbPTbYL9iZqPOmfAParDn8Ott0kDOhIRh5SBteERNsMbQHaN2CbuW61AZ
KbCFCe6jw51pMV3r8oMlLfTvzduG68ZDrgH1cFDqT1yoRp6euMnvsySDNoP/hrCkbyj/u7AnwRnL
637Sc3XEN3pZcYPSIH87iVGJRmn+04nxjmqJJJL2mL8nnBe+xKAR243ptlkgc3jHXFPZthProo8q
TYCCwS2mIQu+FK9vrpVohrmmSy/R/eey1YRJAIAxvE7tCycltV9dj1rMaqLW9z0msPYt0PInp5uQ
YXIFU4G8cHU1ahxUoyMMLuJdFFex7VMU1LqS1CVbEDZbt275TrSMetQm9F6jGyz452bNO3EcvK2Z
dio5SXRE9HjNZpNDU57cVRax1zzaQFtLbagyri+u9BKpi8NCFjJAtO9qwQ6GctI72SZTSyeqMd/4
ROkQygaVicP4GiwCccaK1WD/Wk+AiDNXp3WL8cSA0CkN08mMk8H0R7sDIDpTViXX9S4+DIxs+RcB
9hj27uDrlJ3Hz01Xjjsx5TINj0dYmJZnXpdHP9MFhvP82S++aCtYwvbGm43/r36fE+MxTWhdqW38
nriMU+1y2Hv1kTAI6KXt3YMaap2I07Zqe13EeXcJAajhZdApiuqJ78vomsorRYYTNGrDBa0rQft7
ESLZSSLw439JtqZU/YflI4ESy7rz4XMCNRvSyeNgatrsImsDZKetXiHFmPzJmxEWd2clgvK98+3h
A0jXPmJuMuX/RJXwPfhtYzAFml80keMyohBogvkd4+XNUSimeQKAfSKQDUGiXNelVyAluQa000Vn
Z83LcIvagtsT+a8SQq6djFWUoqSInAaITIVD7votWXpITGQkJtZNyARaUdnHSgXZUJpMkMqMpY8B
OY7rvUl1FA9Fjz8IfXlHpYov9o2XjlRZPxO7FtFru8L3qNYF8MszeaiE795p+ydHEFLFDuNZGLkK
5tBOiD6XlzKfDksd9Kkrsnq+wXQCLyJNioEPkAB5ZGL93Shu8WUmJ8A3KaMw52DpGWiHG7A/KsjG
myWxJ0ONsDj3DBnAtlEH1OQA8CIgEeV7XDZ4clPLrdmvotC0GbYHnR+TSR/nzQ3APbIdJn7eZzuM
kHuJMB1qgxp6KU1c7XFG0h2NZ8DIA7Ks4CftEYNnMBbF60TEjFc9A0uu/A6Ab8WRtu2TEtcnh72p
l3a+m0Mp2MH2+e4edVteeNfI+YNrTENPgrz/mLkJuxbkumVDbkAVaxKxCt82VBhr0uFDRFmDIWTN
fwZbvbipp6W+jOyYFYz0fSqMHkS4qWqX4wBQxskaaAnDkUNdkL2804VgRCC7mqorGONrwBTd97Uh
MwXzx0WtENkndlMEH5QoOVOk2X6Rj4uvhCpqOc0TCDw9LrGyVEo/8aU44zNMszNc3YSIA9Xdja+S
90Mlp563mDL06W1gdH5IbTfyQntvQySeKz1GNlYd1EmneIPaIWk6AZDYYENxsIaC7AUNsCOQDAYt
+L3L9H2IP6bd65+q6Hw1QLnEIjtJ2PGRKqF88G82KiqDFzUsl3TPf54s2B/+cdls6+DmXLPq5+pW
dKcnKEuwOUnKmB3be+DtYzf40c0zaWMPaZnSy344OU8AFqTCBPmas+MvYKbs5rFTmgMOuFm1DRAP
UT48/M9yJitcKqSHpCr4LRpwjUaOOiPHF6Nyc/WHdq5dbr4QAGbuHzkHEQfTb/UyAyGRCdFV2g7V
c7ayyjD4vd7Uj81MqtGQT3VijXCVX3iSyIsNed2j14f1+TbE3mZLPKhbN8hr0+/IzA/qU6YeLeSJ
FexBM7jNqFAEu5G/IKkJYVDlMGkm5JvkTGgaMTSxiimBlbNr6sextVi/mtNmWAFKsumSX6+cFmqM
RfF/qlfSoSn4OrOaKsEEMksw9Vsmv17vFw6bESzV8hW/gfRCjILr0Yte6RO4KLQYvLoIZZ3jUfaF
uQTQd5vVd7YPsg3b33mbUH/OW/TIq0MTFnYztOwzIh8sdQhIiuNW8Xh2C+ySmzXIhDAFGW0QbSbF
7EI73unoIc5urtGK6p/E/x1mvcwqPw6mPIvZ1u0q2tRWPe7y5Q2fjpM/zwrQhvfNV/hVq68HMFOW
ijBVebuNHp5KxQ2oyhtEnuNSF6Y52mfzjbfTC+eBbVplvOeIefKwm343ahVIzsv++Dsbbccsvh/8
niIlPmZu/tFyx4Zz5WM/cA6hdEg/S4CHp8R7ioz0lJKIGwBeDaJoJ4SD0KWGj96RMO4cUxzop0M7
oHZNY1HbXhvFjYjt5Q4EjYuEkz2NBw1s9PAjvyzpc8HisVb9TYcJZwuoxtOaodh5EmXzidCGY8q9
mxk9NEijJoeDTgb5lF7N+LmuwmsGyD3GjhqVkCNcdw0Ofz76Ox502bkjfxcwRJUqdbMhbIztMAWi
GlBLqCvfghRCpPtbV12IqHZKiiyY5rNG4xnwwqvV7o/BgRm01KGSa92HusJbfx/tZZ2ayBBaOxmu
SecJdYIBrxb2Vwg1KsExyGf502aeVcv6pDTcHKk7nD5UO6nscXO2KBXqMqkAYbnhIWoEziEdy86z
oGls7btjS0ayPnZEC8ft+F21f8PCWCOOfyRgtL3TKvKAyDo5ZJEFE9n70YWV42EHgVpG+EaXXcnn
JqH7XSa8F7vYAp8oWlSD+7TwE4rrzuRG7RNQPb+bR81WLQCvOXL7txhxoLZP7dgv3TT6W6ez7/lx
cCwBK1GIK0mF5mtMXU2kgp6g6zy2ZUbT/giayypveyNEsqIVZRwTbMXxDajLW/ov3NsK6qROB1x+
t8aqLPdXAy4N3fxUNRPhVLM+4GbSvtAFqcFlu4lohzXE+t/ULJHiBV9wlCTWYw9vLNWR32N/SXC2
jtyyMOosOLgcar9tdtw2/eJg4iKnKJYXgdGPPgKxOJE7R1tng8LAWhXL40JKL881n8FqeogPuUym
dQy/tZI6k6OBCsbMXOOvTgcgxgNet68IZG06RWPFp6UM92cRjOa/PfM+Ya5bVmwHQohDtQ2RRPuV
4h3ZNgNlXBo/mcZavduiidKit2MFnVcUFxLxzjjSRvdskfhDByqZd3jQUM+AThlM4s0SjZrWZ8w4
M27l/qk+/+11zG77NIAYXd4HPa5ZcSG+W7yRcO8BNpGhTmconNFND/kyjKscHlQciaw8tsgTOqRj
vjf8URXNXmrn9yJqrVDSsDuPTXE7/NLB0yKojhnt6gxU+4+FH2v6reUNSiByhescb6DvFB4g6+hD
9mrDnR98bTGwX3cl30acGupuAqXpJO5JMhm7llf+MhoAWbYP4paTUip804f0P0YA7uJ8NxbRfGAt
rPWdlzwBSt4p20q9uTjOuC3EtON5HRtqR3hKZ4B/B2dbplhh93+RdLVBdydjYqXIbiRImPTxpW/r
1Gx6Ndv/EnFOZZJmRBzY0iNTPW3+HEYfpWMUNZmWcEopvWE2l2YROAw8Ztgp8wV/TRzo33zKnS2a
L320tBXl3TD1ZihMeU/ANs+c8MHbxZjaTt2NZPoayiMpL6mB0cXMXvNr1OFyhPtBEF4QOvkefQ6R
mpldgxvwhjlIavZSTJ55lotGSuT4WrmHMKeQDHlT86b5y1G/g3ocX/dMUlA+VzU6Fsbj2Mq8u3w2
HegATVBxrsuZFSr6cTG+G1326II1DHcnt5AkJX9ziZCCr5IdyHdcPU0s4m0hVdUjsdFyeJ1sMRYZ
K5+7wz+UsYrRtKGQTefMKwL7dwyyGPHp+2uCsRl82WADX2CaamJsnl36l+GMJd4TUrRJpUat9Et2
qIYMakHEnMJUhpRb/Sqhdu7pMiTjQlAtfsAMQUtpRwpBX/Nhr4boCv0m8wGkqvUCVG+dY7aNDjTo
pM3keCEQrHZHO/ZPOQFTATAuQfQQ4ocZrfQTqtKx8N8yfZ5zD25EdfuXH/MoEEgWHgrOZuytn0dp
QoAWIwl99oj0HBpgGHyO4dzBrSKXZ+i34RvdK5zgoYrybz9PqlBLMj2Q2adFDnkmyrqwGL/JkTKE
0AhAzCNdVoapjK9URXK1zhixM0+StzEyhv6QXWZxOhvHr7tFwjePZ4lXk8N5B8ZsqsB4+pViNhUt
L0xNWJQtT6JEVcf1Xh5TcFmQTBsxO/oNA7324zSObnIvC99BKUFg3lLAGH5Zv79uSNwA/uHExANn
+G6s3rAao04J7weBp77Vtjxti0nWUfOqL3ySTD85xw8DITfPQq5tWX55BjHr4tEqfkOD/LL6PAb3
OvvFOcEZZPlAe46OkyLmr/04XfJYhzkk6X/SfbIjlPxRil2CBdXFHX8f7GdbCc5r0qpbenAaNOwn
5K9ekGjlQglwOLd6xCvdZ4v52etPn4GVyR/Ry/4ewYXpERpHoBYyxEtsCBXehtHrS1MS2xi8hfEb
7zQri6Q4L1aY8axkcF1IHTMBp940TfLbjT5fGlie/LRkkA8xohhW5shhoYSkCboF53X4jEXnOwcc
WpWj9C5oaWS8vZ0HsB8wEnXagMJrBrL7MJBjOK6ms25liwAmJAGsh08gyPRb3UURud/g5NTwxY4c
B17ScGsziOGFVCSnhb6tOfVQy/D+OZauom/6QAgaSEOCo/N6xURn1iynXKRNsOUgZPaRpDvz5U11
IA4o2NQIjYibstAbM28Q9ZSx0IkrRdgM9ga+FXfbAUTEyOyH0YRmV+MIzIK8F1xY72pow5jdwm+i
omGL1EYALAt8CV0sBdiM+XhQI3AQmRfBkyPeqpvPqepclXpZRmRJoMW2YEsJaVrT7+ALKFkWWvEj
VSGuAHwQSoFqSbd2faZJ63iLXooeXQcmyHKPteteZ2tcCXgEBqaXBW5ZmdB8e3W0IM784bw3kJm/
8txh4TftlPBxWnmgQrzsn1T+1sqTbloak3LJIgaL+cSshjEUVeoLOPYxDqeoSOT2I4Ck9f7iEQJy
8/MN4YOzmeg0UavQnWEePS3YA+brrEsa9WC4s1aCHqMlLkx8ayz1jO19LL3i56mC1+HIkdmj78hL
kBs++29bP5666xM6Vh9QhGq6gqL6lqXoCvjS8hUKYoKYS5qYMag5kicrdChdc6OF8LT/PCoXdXnQ
zIR6fjLjYbmrTiLfhT52gxKNkn7smiHHdYvqwTJQ4yxQj6AANcaizIv9sqpQnY66dk3fTzhQlEug
652+2JNL6X/5+R4OQyopTpQl+YSaWHNeJ6OCxKlkZ4q4fcLc1hHaxjA4627udMK2QuCcaEalngeS
3EzY1jexxqMrGfARUABBQ5+GWtZDFslsvqkGfcTNIsPyvy7CiR8IyMRx5xcAtk4HLUlBE0vd2VBS
u7Wv3oZMtdRCWjv6LJc+D0C6HRKK6vYKM1KgigeaUuyFLxEq+GuVWAZcREJcYvQpIRHusoMjgwmS
YNvRqRkJbJEYCiC3T8o0DfU38NtexcWM4TlYKzjeQSByb3TD+D8uOUYh5ltgmAzRFyfvtvFczS3W
55HD1kkLNAjZG0uTUyMGlHDPfxGG0bQbAdZ/sQZ6RCQUe/aJYGkcpoXxxFhXdxid7uXvNUyeCxm9
6gGrSBd56l08XTrPJDlWX6rsQyan07oJ0Dft4mhpe4pEZeVk94lbnOVLECGK4EvUhZwIu4wtozwE
j4dwGhvpeBm5o5xw3vb4Fc5rQtXWFE0qivNzuAS7sAZx3ct1BWrIgPXvX9rscBwWh4MuunRIosjx
hk4+szMxkRfp7QZK8+VRFgWfhs9TCXT7gUGIN27AEwkd7G1IQ29HQB3JEJpFDQE0QUE2NEAj8ge6
gWOTK7gZPHbJPLnfQTxcbtTiacAk/uimircVSzGchI+FtTVkUZrh0uUMxgo26qeJtmQDLr93skS6
XtiT3thisRUkoxV3hJONz0p1A9V1Al435mBlHgo9ZxUyN9vRWMhYuAGcPg+IyfNoyNSAJCJzUPyi
zpmDti1H7rSwrLiVndlOew9u1FB+T/RvPu7P19iQyfwuEJLJj7SU7H4nUS3GthuJLg/L262A9LZq
NSqMCGeAlH1856FhS7LcwAERcgisg6C2teChxRKxeule9mp785gHFylPXZ26va7CycL47PB8JJZa
yCWh4/QUIkEmg0oPOSkc0295hgwl/qMRSDXv0o4YTL0S6vzGt7mP2E3+vXlcP85Pwp+vQDcgBoqi
CfyyFzsqqOIM9frLauqsRA5dhqgrXFDlJgBS8jbtq25sijiZzAupQ/gshThYAfNh8iNYoiOQisd0
e5I2yyTMu3OvFJwUHF+qKTEmeoI4YKzZPaPDkbGji70WJ89jQQccsvX4adT10H67SpK90LVz36kx
QoUpv4qILtnkcXmLjNNpPD05LuLFX6nL2a5BcGySOHOws3s75D4iqTJW4aWtFbxJdPK9xKsyc/wh
sg3E5CBzmI4AS/Cu+/fuh/lYEdj6eTpTeV1ogR+7IaxUncXryFX9MTm38x8nJ9FwRDRbA6O05naU
I4gDOt4z6bKUd4NcW27ZWMU76BtOQWHVIVZady0rE22PlJf6Ojv8aSls8nN69MSJ+2jb7ak4Z7Ev
ew7RD2dr76Qf9V6Fnfdyz3F5ncyQw2DveDGeKfh0rz9Pym3Y4ZLIZ/kxrJcbhuAdiCB8djUpuiX4
4RYsOpZFgXT4BrB8mgxQApIuLUJjYv0riEOeJWpSsEjEzhl41nIGYsO5yUrjSFkgxBIvL1i+WVPz
IFfI+qfxYBi1yRBd5xXByylbFYO79e9lsEcYIo3il1vEMQhp2soJSY+hW3iv3H6INJ/zDNIjp2rn
Rwv9dyuomiSFO2ayPi0lWbhQG2WBxBF9Yu2YEnCKRlZL1vjrTnogbPdGiRx8ds6jq9Nntke+/VWL
mmHQkNDoatlTMhhA/gKz9aLs/T3Sps/F9AsX/T6qKl+f7Y5jHiwy23jUqKCT1YQhFF5D619/vcio
yqDvZWb4QWoOFd3S1yyQdH6XmSBmpaPr03LhHLh+fNkcSwHlaboljcBZzk/W1R71JUnT2yZXn5cs
RUlI2B68iH4aHJ2ITmfM8K4bff+YuqIFLOXSWD1aqxr3/SArfkdXnJa1AE3KiC8ZJpFA9O3j6HrA
d8X9ia/XgfS40bUtf94naM/g8I17+v72NoG0yfQb3YXOBnjhk6tmrTDk+1j/cUj4ou6JOdaaxQ78
6qzcu0koXO3a8SWOBtzYfQitm/NKp0vjMYgsc3uPWooyp0/epMrwpsXbqddAGBZDp1e62TkDhqEH
WbLjq5Sfm8BoKi6xMG48rJacN1gfI+J3EoFHtFvnrp5I34BpdcUO8g7PeRZyYtAmlTLeb0+ghoW4
JKHsgJKaaIbVn/C9IAF5wwqVEhDinbqK+CqRACzI0hP8wOB233QdXAS9iqYm82/zvjh4zJ3SgxZg
Y0/GHz5AAYLLsCWgh5AOUVv2tdoD6F8QIKkTRmO79BMpTaQLFIQk7ni4hK6eirAySSVfa00kMeeV
icGgIxjrc/KZsjIRDMCPwBV09vCOxnbT/2r92VdLYIWjE6S1vZfTTE36TNcFDHjy7AmnWOqRPG9h
VVDIHrTn7cK8V2QAooFYc0IqpPzXZNcC1GZnJu7J87viORNl4Jgq3WETeRZJHsG7WS4g9Wl5/ok/
ZNrVZi7Eh1I6yqIb8Fc2VDMwpMtJskSpqzU10I0CrSiUpYIPGftvFzBKqlPsB55vnpYCiPpZct9g
f5nAZQxjYF/lz4zZY/EJeYJNpVZK36y5tqhDNveE0vrHPWG4aHqAHvF7NvCrREnBiQbz5ORPObNX
T0RQbqnhXkJkf1VIwkHcs7sBHdD5nQ0u555ckcX7BUwBEGjJUuNCM4YPbtwtJQdJhRazh+4whbta
qgHlrkMqTvTqSr93a1izoYRoQoBJzFY7QOQaD7AlSLc9/0NNkaKRAtoXWzmHw5sbdvnAlzywE0B5
hQqIISaOHwPqY4RM/SqnOIhlgnMSZ1pxjzXjbKCH3wccqXzRMEI+s8Q9h/0uWI1lxc8b3qkuVttl
ij5+8g0tSqeJAudsadqit0/0Mxx0wbtUGl8+bmnX9Wsc8/jpf9Ciy1/4jMyCzL8C2R6/aVcBkH3c
k3w3M0mpVTjpqRl3q3A7kPslSbwMIqcat3lH+U0W5Dvcvzo/yZNvAA+ZG+U3WM8NDvOdd+aKnBwx
5KLGz1BzVvcXQiM7kGMXesW/wP/H5xebkctI81gKE4sWKPUrNkvbJNto++gP1EYN5N8miy47V6U8
95mpKD4Ofeg4GxNvMCz4Lwtbd3OVWsPwPWDODyNJiIGQI6fyW5weYPzdfloDg7m7GUsWTM6J8m7e
htNHV+IVI2JTcs9QGwbN7/VNdkJ2OmIUJwDyuwWveOU81MlIpstueucCKTRNd04tt0/p8h8s+f0x
Z+yNjU6CnR3o1gYA4P/8QexuDCuyNGQMDqUQ+WXz79heWJ3TlndeS8K1Gz8eco55W1kTyUbazsYN
wnrMBUgTo1Og5QvqL9n6ucTyap1xvXtZa88j+h0ac9oTWqK/vZgCU1D0J6v1lxX3u8WlPBBjQPXR
WT55ddMHDMAw55oF1fMNs3woEqLg3g9DbFFWdnAStT5Oyp4H7g0RRiRucg7OjQxfC/p8UQV7dvcW
AiRSrDTl5bu3jy3TU4g5b5W5uBTwWh3oMXVC1qJh/mfbR1jcRbnoFF0xkTxty4aCJO7gaGUAjkwl
yIbGhNdK3JRHGUl5UYaUZEA45T5ejmoACnOmRMK98qVsjAPwkh5MOSZqm/o57rqrhPDQS+FEG+jd
y3bf2yqMAb271IBquEDpJgSDVFfm83eoFDx7MjW9VbS5ahzFVRGj3VLNCz3p55zRonFXaaK4yDyv
/mmaM98GFQ48wTRHVxlcjGiTK+UcGLvrHn7VVSlCSZypBfpArd3J+pj+MEvy8aaOjNftRglihoKx
PkBnU54UliTLZ1kWW1Zz7LECgL68NIOD7QGWLcmYsHaqodqznjG/isBwlKmqOO7mi/WHcxnlu2C8
3rnCmw3N4nijYmkDf05lWijL/comkHRN7TxByY+7DZlbe6ZX6zZk+xn98RMIq356mJrWlXRjoIY7
FCbtz0A//fJ3mMDWo3cDKj3D81g15F62aihry/ZTTDBS6QP7XDFxhOgNjHTFwc0hzJ4qFqiew8GB
wGE3I0ABVA1/Kpfy0GQidDO7hrHGrZGcVOZCfFNgUWWOgZh2kSep3wSpmgd2i40mNOy6F7uN3iCQ
OuVBmsRZwe5DMx1VdCZAkmcU8zOKJE0q1eF5KU8tH4/V2FiMhKvRC/4JGkoXejObEeggnwN+fSXq
gXIUcx/di5MbWD41GRt2mwQOS2gqOAUEcn+b+N5YUJWxxZvhPbfmDGktIXNKL/Oy7w7aU01b/AuJ
73gjoNx6Jk6YMD8y9W3p0zJS4VvNuN35zk2WYPEApFkHdE6XabOU1NcDwC6BDdYBVk+4Feb1eBBC
+/0T31KgeOjBhbSFcj16TdZFM6AZJmONE7pbHKF1FhQ3OdzFPkVHuZ7wytzNsQ8UkACTzUbvxmHs
RFT4fJVDhhmh8DEftxnS4xrQxpqd/hfuVdRhYfrt9GxyTVWtunQGF0zsODJwm3htPzViq0/xt7jg
viUgud9IX25E+0c6+tkNUCeHurPS5pDmbH7EDzfZD4UoggAUu07w6f8IpCyiKOuk5FzWWAF70TXn
ZFSmX6e8HavliEoMAMMHpk4P2BJ/Eb81L1ZWkK+N0bqifMl275ZMUj/driG5SXByDGyR765nQ/Qm
HfeRY4Xcb5sEmaNZ2XgQwp/Qz8u0whfdnkuYpG5zacBm2ITq0EXY/0kGjfGfpdIoP+jl0w4cV6dx
bIrx5drQlhpqnXVb+cI75ytbWAxeUl/X8jXY3L/Vg/se9lLnls9lndhCGJmrvBYO6RMLZ/5yZgBz
UQ+cqXXU++DrWZRi4Rpt/NmI22kIsDDV9s5XlpEQfaeCjdHrejvcoFq5O304ZC6r4bgcgTRj7gQL
13YqWIVg8AGo/HtrYkQYGcmCxMHcRtmKG8971hBQArXhFlm0S6vPxlOsndV0bcwKr41RDNLngvX9
vsbGOeTNPg09ofQZPEmoZCtqSZLlF5aRHeMi4DyGh9oygU8bxIkK31D1UbavxdYe7BDNJA7iB9WW
vTZ0JW42B+hQurnbFhCMybVgqlg8P7HyYRjISnxfvMcKLB5PNhuMbwtKZ8S9ir/4H33Cs8dfw0ef
q56N/IxDqhq8/CTWKtTO7WM0/MvHxGLRJDjo1187HzwT2O03Mjbwl+/r7EVs6Za5BegNQ8iGO8iV
csFZ1e2PxS9loF9gkfIoLGVRwtqwTQCzmUypyfh8nT3+2RkxlLsN3iAMK4gfdAPxhrduJozWMZ6m
PYG/97H5uvNo0ZmHGYBdlSsT99jIQIc+KdSj1fjxgQMNnDXFIssFy31aKK+8Kx7oZJs+tyfjDCsJ
TuM3EmRZvDeLMXDQKj1nchzbmH1oDRjhRoQl9onAcx8FSz7fvHBNJQFb1kC7CP7tdAYBbmYEO3yy
e+xX6V6Rq6yQQbu0EJDbg9LXfRSeXsOewhDiII3deXj/qdNdxUQPvVHCvL/K125pVzXEDaKR/3E6
jxv4XbpnWuRxN7YbwxhNEez1+uAVPuSBL7hdlwabQLytUfXLE1kiBBxHPFCWgb1Y6fO4/0+fvNSt
QjpTAfc/HgPg39FJXBrRfimQroUA1vWPRPgem/VKPs4wPLPN3duKMBJ8xPVA7dbxP5gK0EvrCpjc
ZhgT9KgQgCtQyQKwzaxeyuGWXt7H0CcxbjhqjtsMp5ciHhT+cGZimcDxTORAsfgkMplIz3qkwZO/
ZtKXfUkm+y3Rdc2HCQsn97EKB2hQFLOxiHen+RDfZsOswfpQFtCgHNuhzNBqee08K3ePdnRKC5yL
n/ALz2xWF+xzL0wq+AnBE1elJ6ElEXamvq+7PJINh/RyiCeuqhJRDe8y+sB64rDuyteAqrCjmrlq
xXc9rjEcz6tCe+vJ2XNv7+foydqKVrCZ8uLE6NYxQR1Mj6hgMttCwShODY64alq4tNJdhhZPx+Um
cdP09JNN7Eh/7do17L0nm4IQjy8k4ZXtOFQacDk70G8O96V6E1pwhacEWTmwO0cOsOlcSIOfSZzc
qTGyKeQ96o8vsssc6ckAQILdmDJoTQdEvSFhlQTJWDfTodJwvbNjdHxS4elbUXFeV0oLn+VLlvdY
4GnL0hL3e/AGkmYvVUTIXn+2ZJz4F0QUIp0jp3n7X0mw03P0xVQV670j6+WXiRtFO6htn5xVN4G/
dfGYHIzS6f3CkvMVPqHiW3AjQC1EgUTKF58grLeBfN2zlXK9dcDAYPTtucRBHn7fgqSwTjGsKdHH
NKrSDmcXV09DE35EBO5FtSDdFOmZqE0moTpVvpbHLBmpLtwNa5ENLqqcRNNfHxlSsFV7PiCgQRlF
GgrJLPZJp+NyNx342jo2erwrtYRXOMwfKAFt6F7AVTSa+9+x2PqCqEQZUpl4PZttt0oHqyqAgrFm
mhINfOYAg2eBXZaykBi7H9bHbrWDeBRl4eBSl/Iz3DGPKov8TdHKhh8mGkbnmddVH0PK5+H8A7ym
/owPuhxWk/V3eKEp/r992yCYYKjzPEx8Ek1X8jOIS+XR3JcfEbYjZ2DT0LXK7r+16Xa2FvTr//dr
NsEuhbNGx0uXlOgCPBHnh37iCsI8i4fzksQUgm4LWoNXwIqW3GlmDxq9PJXJDtQ5sIh/qOZ6DpVi
vKxO58Jo3cfbOerFiGiKYUEgwBcgpNQH3wz68R5V6uiQzpCEhxZT70OdHNHHZTPt+OARk0x0jWRn
iqCgnHkavhCgfW2bfnNi6D7tBGK2XMLT5JcMczqn56CcsJsDtXWH+HlXRBC1ZuwG65JGhSOOuzdh
I+QgQK1o77fWbpPxkr0B6qUQv620/yw65l0SZdWanzC6fls/T+KVXCMk8a9YgTgbmNobMNkFFHkP
lyQe+LxR70ZJcmd5/+imRyNYhgwerUr0pAaMnCG3EcuwbPtLq07Z6xTu0jgridSNa+ePUdr8FBOP
D/AKUq7AB2SQHSfrMpWqRl3dLVg5xuIerXIX/NVkYnZpZOw0288YCa9WIZZCfJWhnVNkrh70hGuB
b5nUCr7QpPrQgCwEKhYewc+gPz14J/s3Y4t45g2/rjJfOsw7mqbU9+tVNv9CEtHvt3WXYImjkImC
YaGe7S17J8zt89GqdDquZu0aJGDmKXgGGRGXN1UmDHP4rAU7eepziZEfBB/ICbcW9zFZkDbRjypG
E7g/qKygNRsccSG3K1ekeIjNKuE0zkGUgR95kr5Sol4WSqrTU+1WHoNZIBi+B2xMSyxeVKiwFLTa
3w22J0g7HSmHbjH/S/1WW+i7ZjC41w3jPH9PIB62T7oa/x+DJLZ52I4QD7jGQqlkpTTYJVmOafOS
sRSr3GCywX17ZgS2A5KvzJgfEI6z3fIjhLJNddyw8XAP6x9aCVfkfVFie4dpj8DBWLs2PnHvt0Vy
N12rdDwwB1PvZGWc9ttRXLFu7lxLJ7JhV+W8N9+LKXHisPSNquNX+nqKBLHLd4maTSJ2i+zmN34M
bBiYfOyp2Ai1ZLUCyg0MH/2ri7H9B5e7HcVJaxfxyJKYei7gwZQY2VQ1wRXWx20NfGH9RfEeV3vx
MqHV5XMX+OZpDV0+UdGeE5Ye6xsfbC+meYEbnKG6bBYSSlONuByOzu+mm27SYaj+MYfF5Ltb2V79
ZTnXc7jpgbu4/GCVQmZdKjkN5hYhS3EwiMPqG8rgCmUywYMK7ehIXNlxqX/9vWOEhhVbFM4sjKg9
NeBsglj23gDq6sLyyU513RyHTepIm0shR59V8F+6koHvUIdo+xViZ7rUQGvjVhWoEXtiZaUyM0vU
nFLJrm+jUGU6N3w/X6qXBL5bTGHYXtl+UoY1YkmUlsNPmOA7kvMcTgyvHwItnHx8zuIeYGCOnCHh
/KYHhTfDKlHGpkWwiqb6fI0m1kYimMvgTmbdte7m37QNfsP/nSE0Pz5RmdeEf+1SqrXT4AASx+YA
U5oPf0PUysEvwXJlRjCbZZCzsiH7jcTddHJR0NSYIIVUWoRZZ0VV1e84xOwPRgAbLFOTxIzDv59U
2PYXdbjsbtbfta8Q8ZPATbk0lTPihM7e30DiIDSGcsHvQ/ogDE4sGHaGqh2aHuyN0gqrJ/o+dVUb
NXG3hzU5Vatjngs1ceToe+hVSoSUREbfaZJyf1SUrfM+OZSuDYuIfjd3C1gMp3l6dZBWjO9fNbIH
oMaBBS6QDo0YBE16QaZunynL8aEabuIhzWth4sAuJKvIuF2ngpDE6nxDwVENVK598lI0dxEt+JZy
VT6id6x1toDxYwk7aefH/mEq+DvvWkQLH6Gny45FTJPP/TrEYLmoAH9K2k0XV5Nz0DZxWGVSk4Gn
yFfLAENPu8WdWSEFINrddopsnvrm0yRpvoAORQP3rDx1Dob1yutwZgjmMltN0UjpB+384aXz7OWq
JPzMR490Q/EfhM+kmBJ6S4FkUPuqbVqqwk0AkU/nLEUv6Hd1uSzHx7Cnfpp2Gwt8vvD5+7Ul1bev
cJygPHPxZjQUbiNnr4ZGVAR2eBMSFd9SY64Ems1L3MEcB0V3/br/9vAYMECUsSnRGF8wFFBX8nvW
MFm+xIeGqNTbNpQzzSpYFIfja36Yf9g80D1j6fV+WUnpmesmkPi90ewI8WHhYQnz2N0/B5bsQNoS
y0T0538nEotnidZJuhKlmqMJK8JP8/8qyL6HbzQcR9l/f1E2DyZbGoy8H6bijBqbv/IHGquGYuy2
VsyX7zzxeF7vbd8xhBWxh70lfSvxJZYP1LE/xNJn4C6JkNspxkg1pl83mdIddiLhf+fBAbTgzeBf
aefPxBRbiCRthjqx1ncUvSTS/XbM943sFke4udB7fS1hnTiGzX8d6rwfYEtSD0Mr9Z+aH6Y92aO/
1cLM/u+VR5dZmCwAas+sEFcpgbEfQVge2ZdUnt+6jAuNgJfaAJo6abXAGqo5wCa6jJkvJdxyZuZm
G2TMdyt55jZWEA6zGt0YNlGR40ubbUb4I5DtF0Tzae+ofDf4HXn1RNJrDbV8CsVwWW94shDLWTxk
3kUZ/GdU+/rJ1G+vgl9TqFkfqY6cYC3stdmzQmc5ayHQnlLgLl+TxNu99z5TYYwEReGJExLBZrZs
/V9NWUVM8MfArGQZLoDq/Mm4vnHfz5ohn70FjkqCwQQIO5x0FNyD+MenGNz/PNzceAWjoWWRWMdl
2fLgb8ftUfKZa6piJy712IK9Kby0Zb2yA1qbyAi2mnNLya1GyuHhdpYdgu2RoKkWkUqi27bmuTGU
ijECeYHY9j+CeawraQ8GJgd7HRlY8RrpNR6Ufdsp9nxMNsPyXut7d8Qm0Ift03vuBPCdutl/1DgO
NEx+LqgP65pxCty7A+EhmjhJmOVHEE0VF8BOPhHPMTZedb0gTLS7F0slxZQM0HQeYGNFpaAPcetf
OohNxHTz3Os4bChX0sY5wjeTu+OH1NfGYq3Z6xlRdfx96wNocl3+E6RYuResOTQ1AyjzwuFO1C9t
Op7NYpbZe8nn4p7ydeSNo5piW/qg9UfKUDCdK4r/xYJ0jU0cSw9ch5CevYp7XHX8K/deF3NIbiqZ
0yRqS9fXN14ohrTSc/Fhihr8hoXDv5EGh2aGO/2CQXBSN1LOnGnJwKRt5FAQycYOl47AeAGCKLJR
erGTMofg9pw9BeuiTIJVmJOatbdXpu0pLLUrqCD152qPHO4n30CMzoPjs4V2ubG3JUpNIu5MKlkA
chN/m93TOxzDJXd8s9er7yT3vyKI/mp+9GjfJzBr0rF3pf4Ysj617p+rlrZU97LrYlpqUFgjXsQT
4hxE/PEl6s/s2S9Xon0VqbCRRmR60j+Vq8pc8EivtMPGYA+CjstbwUxBDA0tpvEe/RgfpkDZ0AbI
2bheBFEqh3nz337a2V5Frb5GCLoUsOAUwm+I0hov6vrNCM0zmuA7QOqTt3W4bZKSetWlmZs5z6q0
7uxQnuPBOPyz2jBIh1mq+R53MtJ8AEa/zo6JQEMvyMYf0wUBsyczDsNmheeOzBTPioq8LzNjEn3/
8UeRVtjtvcz6bf4Blvbbdjuty98s7aVM7s/CBcgOZ5dOPA0lt0iPbOs2OURFNVfvUW+7nBetBLhk
PnUKR2likJSh9wMlvKhNDXbBo/fVHuOSBl7fZTVvvTaKW+yOApZKTJTQawy/aeyf5SFygWmhOdmF
Vjx0YYTvnUgl0ODhmOmDySSObqVIBYIAoOIQKcGh0fu7y6WMPf8vlpdWgJPA9MD/9TtbWQcfO47A
wgtWsfMMHqVGrNCkh7gnxgh/CJwNNLmbng+EMuAs2vUizpKtE4SCrHsJ1IzL8fq8j7eBEcZFx6JN
f4GXMBDoI7GalLFVALgbMgeftaFV4BqJipdB6D9u0O+A73m5Zg4X/JjVfECEAtCpogMNuIDrN/8A
VB1FcwGSZHJ/1WGi5mSUOi16egyQOpsF1dn9/tfPhKVNyCB7WeLbMM8KS9IWSd4ca84Ls0zi2/4X
57ln0ToaSp3hnCzk9lBEX/4n/XuUTFeZry09+tIQhQw3OMpI7/8nU6WuBc4kaonoFyuXVUjUZHdz
l5e8utyI2DbApdrXUtl3VfwR1epzj2DsvvDPEb/pqbQG0G5IkdlG9ZetPdjOFBcnqL1Cmkp9v3FQ
Tow9h9IXGvS667vYljDUEhU/Tv8irv5sWNeblbbgHcqgziCg2IsbU9woi70NAIoJkRTaQgXvw7QQ
bbrVNUbbNU+Bj2iKBlCcdX7rKkkCL9csZZhzQKsz0NpS8hIZ9QGUudGM6cWEHnrXRVEH2vQCNdD/
5CnspgH9XbTA8YDgEQFqaRe8t7mg+VaqoDHNfuwINWnkdyli4EAkM1AcMqvRYvy+V9vQjQKWwvVX
NX72OmnF8M6X+5hxlePU16og7GKXEg+k4HwFxQFzKroZuvrD2vVeaEbafG2pDsSpRHz73ADaeZyR
8O+IvQBvL6mxr/ihNPVkbZTIjSqGjF5PjWrEBYM/dMs+yuVwSJ0xWobGdpU3J4549S4/yUR9rpJL
Ikt0Cs27ZzM2ab3RUEZfzcPaM8hsn/xvvCIYcvM1i8PsPO67WE137T3g7lw2FywI4kIDuMgKOcg0
YTRIsmI+3xDKim0UNvAO8VkVBMRFvspEAQPC5YA8v5CNTvZ2odlnVY7mEwoyAdt2tbzu/m+P5x+F
z/r2BZYNVHA9TXsfFoov3TL5joVyG7WwIPryyfyCsDsBZDoDLVetqUHhm4ULBO0IqGoKkvfBUfgI
UrJuIOc1M9dF2o8y2aXvh8sRTw7POuhc5MTmv6CxIvPikYJq6OZG4WiQ6olso32gyCOu5fUU+rrA
MbHnifxbpSnUkfFODFXcB3VAxgsJFNqh6Kaut956p1i6WuXbVjmV9PndOks4zEcyK+ePY3cr3V0V
HQ5svodev2J9GSY8n8DeKqJFGusE0wPDV9Cj7+UAMKC5tqc38dN2VYrnOrG8MZznMlQGosmWswr5
l3u5NTqJsYEf+WGpoJZyT2gIQYBZrasKa0wDYeO6C4gRoiUzhJ1JKx4G614pSl3EPu0yY3xmaSoj
1ys2ZO5VN+Iy9gcIm1qaIk7dKneSoTgoAW0MlpWcDUPRsJ9JWs3C85DibxtNi/6qsjPTix1qTs0I
W6QXrDj7h7K6jJrPtKOKwXLPwok8QSKaMYz8q9CRdNU/JoiO9cE5bqRFo/WPO4XsX5aqwf/+lnyP
fpLy104ipEKAYchCej8HNxPwI324sKlHnb2+RzfN+Tjy6sw9lSVUazHejgqOQZhm8NVauH6eQJ4O
6ynEYp2fPmywT5BvvWttFOXbpnvRZjae3S4SHmywjnE2K8sPTW3VlD3Efxro4CGaEkqLT+pzaO3/
FVC/nVaFBVw9ddgFJBT2R8VeUxAbYWdaWozZQBe9hUrTWM8KMECnQc9YG3KYPFkBvEkDeD7A0mAr
L8XZy2It4MDGfK1fOHHOEpnAgGOWmIp02PoKYLeS0ZE9d11K/w+g1IrEv0ON+p9mQ4lrSD+y0zoG
nnCi+O/lvb1yQ3tHZBsKV5HnN0DvoHWljvBG6axks8yo/J4LXmSkliLn7ZZ7aTF9RB1qOLrct+Aa
Oa1unVPqc8u3Ht3wzEDDguWb1AMsDCix96aJ9A128Ko8t/f3Y0jI/XhltJdsEcmPrh7+gznjplDf
7MXrDkUos9d73pgfrWp7B7jS4FEfY/v+n4kzShXN6hohOQ9FVcGrrl7Wha0zkE5UJkYs/2Kgs0rf
Jm7/cEQp+kOotR2sdMjHfvHifVHR3a1wIsxeAMF3p/5jmDyp1+j9N+SroT7st6c5RGwB8rK2a0oX
bUSYoPDl+brvniToWzPdxR/E8+Tnfa30xOuo2mUqLQkob0llWVXXQNTfBNljMdnjjY0WJDSNiOrK
Z8lieYyF9ibqa72Pc/ZPo+S5OP8h3FySp311CCYpUsriFIbFVaOfppNJN3W0RhgkDdUa8vLgWll8
Qx/9RAySlEvnHh8y1jg8Y9lrhePT9cJCAG0O1tFwi/ETCWHnHHLv0/CGX+zyeBigrXxD2Rte+rMV
ABwNXPjov5FUiIEFA/UZZA8cEVqalHbgpxdhuarDbSHV386eRcyj3DKa/8Ebnc5SfMVMAq/8pXXx
/BdmcLFo4A4Ibz6QTms6qikqwyds9EO+LjtaS6BZL4dmS2a1JubWGv19l+LPClu6dQk16e1V84kM
5ApJC5qhL56X+6mkVIDMRhSo9EsMD9AIGfPzJbKLOh7Vp4riWZ4UjD1geYvv+0IHzhFi2BMM9l3z
JV+0z//YwC1T6eQuMtyDqFRSTwJPZZkB4ZuGFqCFw4ARD0qY5EdVDO5AEtLVvMN1XP5zQBs0p9U2
XtP4UPy5CBiZ6CQBgsWeMSfPP9RzoRkz0RSacxyBtTG5BOywL14uifIpkU0aZAbK+hv5VRSkNqJo
K7ARgHjnuKHE/um0X1ca7zTGQYS3egzM85sPfeFVaZ3j+O3YZYMRGrs+FTMszDa49fEwkscttrq1
TPPdofw1WRbpDG8SFBkjnBYtOoKvETM8rpsLQD0VozW9TjCWkZf/CwmYTWxVZ9fJxSAGHFdziebB
vh/8u72s82ZM5YrJLX+F19AcA6qW8HnYni9pKMVSPpTKXr2l0p5Q5u/VU8ZrvbE5VRNQizpMHB8c
k2kSip/sYkAiewguB6WSZEE3IvCPmevKE4XlHhcpA79s2hd8msS1ylqQYvWXmBo4NWP01yKjRei2
xLaFTcWtZZZSysMFKi5Yw3Y+n661IJB5MqC2seUeUH/2KWROuUJCzxy79iFKuvLMdMSpb8XV5LsO
4tmDQ3A8EgNLiUeLMXEr8jUu64LywoCiBNJkZBad4B1RXx4kDDjtbWbBB0uD21yvLwpKVsfdsv2o
zw/Vmyxl4dOpHgoZSiAbWCQe2RjZx47RODpwPZmqonD1Zk/yizuYa+sWgQKl64kP/aOMkBfc2/BZ
Z6fkPWlWUhWkoJrhkMBCHHvRzeP582XMQVgY5HkCAYpjAicmMV510KgQhmHh98GX2enDjtC44o6g
1l9ogKrDArhfvlV6HGndf8WSW3roGUz2y+wCgjz6REksI0kK2rzSfGJvErigF0HnelLAIggKMKJ/
NuXR41fXBuzlP58YPkZ4dU40FSU/PORfX7ZZAmW7DMSuYl/BCYly1cA3HuebTDUK+5mOEt8bdQ1u
PSKMA3ta2/HMUPDHRVOlxf8PoZVegzwYyLLp89GvkOgPJDllvrvtsu+S6u4JMakTf4cDfgkNoe+7
2UI4FncUyAE5/onWeL1/TV/ZHyRGJhYiUeKPyP/LGAePxw7RQSfZH9BHF/nmOkRW8ejMe1WvKMY8
fNn67SG8dfAshmQ8UTwV8FA885bZu6oMdJ04NY+YGVJZ0eyFOJIe/EsXkBluugQ4X0jQeeaVit4Z
UYjsqKbVbNp1OK38tVtJv0FJgBvafSx6ddFXe+CGCDhBuYBFVgVboxIc5zHn/SYscOkjZ8yj14D3
C5zUxczjivsbLV6eY3bxwbzvR/nhajqiLsj1ExMORPUz0Q5rwkkNoHh/1s372gb/jVxvXl0Yf9JR
V/3F1zxQMxZPfO/UMquKM6umyLlDXkIczUnnRjhNHS1m+3wW/uEyOq5Wy+8DEsEEQ5SnSdVxRSKu
BcVFLqFLiBUXMRzOw9IMVcnsMKYH3nTmzRAXlqf4607UXQrrvV4x1oqESt4LSxSSB0aD/kf5vIG2
03OgbM4NeCkWwfVVykOYyT927HzbCfFJN8rZJb6F4xI5bqVyV3esjI3nxmpDfye9S9qsdE9JnxH4
3JWnEFueFQWMM8AQiRSDxN/1N8Mepz4jqnuRVVTJm4yhTdFo//z980LfEggvYwqb+egbS5/Oat2P
NhtOZvqD1iTA6+QyxDA+Gln8ZXOSKPT6eWAzmPh8he8u5RfkGLfxSOHHBX6kGfONfXKdbJ1yyeTh
VtCK+3x9RzmH5srCDI6u48M9WcxPdnAn9C4ZlQQuQ62OdcHe0gA/S1agHiAYEAJBl4J1+1j5Skb+
2yAdTfXfmZfgbGTWPieQySjW6CHd0U0jB+g3M+IkTLOmmXOcZllX8PKVcwOA4x+KxaJI0h0TFX5Y
K2wWAEEFuhRPgHpUpdAxjB3C/70dx1DtIbPgCYSCud/8Hr6pPwNqHVpLo5F1wTIiOyXMPib6mfQK
LDHOC2qT0O/0b9VG1Z6jAVu4TN5BTD0SvgMxHQ/a6YWyF/4xduUWt5VRiERLfkGOxAF+xHNfKS7j
arYU2tk6s7ja7fLlLpFGnb4J1Q0Z9CATz727If7m7O2gvfmyuD7+RsQVPKElSe4Oae7HK8RNZxHe
+U7k/u9ofpo+hhhHKAOV4VFFHbKGo/s7r12LaOmkrlI8c216JgJ+pgi1UDE5woxpsfBvgu8Ia/P0
O8db6DBuhUccxEHsNT2ORsqXng4yK1Vu3fUCW00C1A4lp9+ihTTzxfijGfN4MEUWpcIIUjeHz1+h
ZT4qdQxAIMJmhy+lI5BRA4WUVCb6MW7akNntQVF+8pt6s778RkjSvBwffX22Fop66oGMJsDdFG9k
Q9fMS+h0xz1C3uF+ksNMF5ugQNM9Jqtwf0EXu23qEMjZcqpgCVRN5+gOUXDysZffJCbWEyQD46U+
pBzcMzJvWxhoLcpSmkhsulpQGfZa3jMBkm00lARs+0oN7oXzD/T7odnlp2xiRxZzErnK+m5tQOCm
rm6tE0Bf7/mb0N1iMGaPuJrR0MmldA+mOqfzSrCmNVvLULHJxfz8++LwBmFbD3rvHoEYY2Cc7Xqi
G6B+z6D9uVVdQLKT394b0imEMwudIHPwLMuyVjmLGGEexiA/prJGLTrcetgwxLP+G0MU4lcxXVeE
wrwkr/BFvTyxq+XosNnQ69K/ai6BUjW4YEabkpmWSKjIjTXmQo6ay024OEmV/o/ABJf1m1mJ309x
jTI+yPirZed7Ud3nnTPnAwq9+TQSShh+iRwgyMaApkVye7q7RlApDAyUzgrxTi0BtsEespzBZS2m
tPJiQv9jZkybLdlmCr09StPnaMR2jaNiTyYcwhkrr8FaOsb0o4zxC+xi12x28cCYpfghmwy1UldE
IvRANFguOvZ5WTh6Hx0/Qgq9670qy5YPBQbm28DsjwDh1r/qC3P69Ai+ppPqKJY5B8pEDosDlxW9
gr459fCSkPokhQw5Iytg91JpS7bLxG1W/VavudWijmGAGtolyNlurzXaIP/HHgGGgNEOfgbagqJ5
t9wjsWaJIid0hEzJW85hhpe7iHw4d2f+hF1fvtCbsqTz9S2LPxv8557/TZZ0dJK3NUfP/gPt9W+k
t/MW3qZE4W4i0vrcPihqvDJI+8ca7Fag2OeJAYwjkL14xdMu9X43WmZAGa+vplEZHV17is3GQam7
6B8UuxKwU7xf4U9x75HHLfveUcsKK6LNMaB7ENGS/h75ycQWMAIzvIy6C5qprToyY3K1u1urd1qc
wlx3mLS1CFj1LCJKYskfqiJRvnic4+W+/FeP9Azt7OFXsv8hlqFwE8uFgPvG2cq43VzkuFI1mq8L
gA18P/xZQZoFnwIlHOJIkqTUgLBRwh70LxFfeuksNjhibTLT18nJtjZgUDLaiyQzGxQa8VDB1x37
6dYdPNj6Zx80GENF3tN6jrpECVwKlrRp82ea9HpnOJi08j44iuzEaE2SPK+TxaD4ZBTBynnyau1p
HL3gMmQAyfYsCXqYzd8GFw0Rsyr6qKZlqQ2CfMoVJ5qtyQBc1AcKA7j4lDNBlf9+t/qkA4KIWHo7
zKCPsIwSvvDjz1TN4+DvsSD8SgMNpt9rDsBh+oCwsk+xIUwIUNfTdI4RSMlE2U+R2JjExZRQgl7f
l6WrqYHlsdBeKDt68oBHB4SjmY3tQlKe7ZSXk/V6X+FZM//GGySh6nJajDjnBW22i83oIulSokkJ
R9HHdbsbqQv0uRCnJ4OcIaXLa92szDNhgz194pqhzNpyNV+yqYtOUUlIyKeE97H9JulzI/OH34C/
DQ3XOjQsAqwFbe3zf7PeuYF7/qwxmnmnfi+flFchyKqVGxMn1BI8GhPOZVJeCPGaw3ELe3JJ62jH
xjtyVkn3Z/EF5zvLEPv7ExK8eBU+5pd2hdiGYqrS4dlKHjgz3zlWTYB9h1bmOHHAjOoDoRWcwipJ
sZwOdL5lhpjAaQz06wc/x3NvDNEdfUwfZNsCOTXtNEBCOrotbFPnDOaBLck/4KhSSlejqeXPXWnr
iDHcwzoWQREcujs4NiHNUYu7RUqvBggtFmKwzqk2H1UK/gBlYkrs5pDjdrwTG8kaSAnrJYYtUk0w
YP0Wr8E8cNOhfRn0T8PscKEYRzhwo5VZmHG4arYPrvMy3Se8rx3W7JhY5qmm7Gd7s5f6DGyYuqlk
Jr8+0HFyHZrT5p/CIN1/Sss6t8EEOJG2gNsPSQ3jyQDsvwsjVWAylzaGJ2iEBXdf8As+60U/nOUC
a+ZhSazoYlxY63MHU9M4blYzbuh9sh6IAEH86+tDO2ejBdwvfCaYDmRJGiA3pifsdnfNyfwFffCS
kIA+b05f5y9DkWI62frbyyDnTx0Ud3V5tHR5AFmggsZQjXyshoyRCIgC5wvVErQM5TSWigivhleV
dpig806g2lB3Q+EJcwmi1BZeDqGNpkJs7eL5CcvsvBzM+HCWjvfg1nGtZkrC6gV85ANvhFktdc1/
UeYGTL5WBFUu1HWULoW5rfPgOO5KjT76Qz+o3icDuzvgcYlENBykxG+TnCHb5C6aR+XUTpi3cHEW
77fvD9quKmq93r0++Rc2Q1T567F8rVgXyk0Do6g1Bk80Fl/IsAcvAJGYXVMEurhPfN1PWsOKFyYw
azGwo0VLrlWwOPw3NLt91i8wkS5XQ03hWuLAeqipEnedVyPQg6wndQmt6Ibojztbru2pJumAhjBC
Oe+1lnYJs7U0f+AFja4ItVIl53WX8Yhtyn6Fex7cInZ034TaYUDylEf/jh5qtDwZfRxCkUOTtsXM
iVb3Dkyi9b16kerTKA6gd4TkoFQa4EdYCprRshsPFmno7U/nfVcvoFTMI6XPvchsBjtrfX/49Jnx
eWyRCUdDPwiCJ01BMtw1uqL+Zshn2Tys6Lw0stMmjByUjLRoVfJAH7Oza95KQzLq+CeDc9nOXR3D
E4L4p7pvTsBXX7UZlWnIe5L1Z3bzF93ZSLPycQQZ9ASGI45+TybwnbMK28Pg8Ux12c4sTtt9nkPu
yF0rLqHf8jK3rOh1pPtg34ciNeGUH++8rANTq1irnMoG8RZbP8kaNkDILjLboETQMX0chOK2krD9
8mwnm7yTX2E5blh2Ux4yy/+//r9F42ClX4hpPh7BkErwBa0+ueA99xSCDs14AUQMp/kUcPBvj68Y
xW390hx4nH3HATZNKayi9K5XdpgBB8fcyrSx6MFrGlykM5lO9wGpBgL0xh077CY1mpaVPRWolzCK
zTJqSbAgukn3IktGD2EfkCTrykLaLumcB9och2ENuk1JL2RhbIazIvkszN26GdZlvP9oWxOCESMu
yLRtfH7GlmCqiBSEC2zajOI9QoyNorSxYkU01lWMLfkl/zHHK3l3dlfOaEow9ffiN3szuXwtzbGX
0mYEZ2h54onRrf+dj68d73Jkslx6MXhuX1oB/vGCvPh46OTm41E8uC3lC1qvvKUg+rIjJs52e/qo
/MkjTLK/25MQ3jkw1lWB4jN9UWh1nPFPEkSXga24B/TfS1oUDQhpeFCVzCdeMDRNHL9Zt9RsCmNg
i7W074/PWsWEGVtLXHGaEgjWfK14r2dzV9sGO1cUl9jYSDtyEVtERrojGmxtpjkyztruTiWc1wxu
Gyfe4NikHOVmFbwgb2UlogScAkfxeKcn7xi3atpG4JaeCroj3rabLWoVj76nYDnFiW+fPbrdpZa6
Ll1lRp/7Zl+sUBEnYtGKGRka7T2PzC9DcCHrc/ewFkl9KDjJV++4/GqmGY9Q1r4XNMvAYxESxlRJ
1mV01LUxYrhpCF7LoUg7+9bvKxIz/BaGFEFbrkNgMT/ipdRyszZUocq1/u9+SamxVBZQPRcXv8pI
YvzA2eQEztgZGgor3LBef6dctQvm3awSDbuP7h56wGZy4r6XJ+VK2dKL4zhMWoeyJadGMDvpHOeT
IcPqvWbJ4xRNJEIiyCuaVFSuGuTLBPC3Copirr1PNaQEU56/5Xjkhyh55WgyYCDwrEpuRJpU0dDS
b8dyga+alwVWh2PJvelAcZCS5poqOD8TNa7EtYB+rlhB0nEHNusZ3YaoSgFTE6ZAf2zi70xB4rHz
tMbVNKRIcVUj9iJ6fCvmm+pGKt8JwUj9wLLfR6hCrTweDIOPGoN0meHcYeLb4vwXsq4rvi6rZSsO
yAL8drRsdLLqnce2VIXjc04ij6FAqeqad4e/ZQ1Jj4kZgk0wvu1aQ1WtUjWh1xW1YyfNEXhictAq
zRMieRa6uEt18jHA85me+8GSmO59rX42KGmZ1LWkICWQr2vn+dFuzFCcXVol5rHY3EQX5U9AExGd
5heJy9+rjlzvYZmF9+deBGq5BqzuT8dW0OBEgU5MMlX2PBAs5NqKCzMMK3Cqot1cI5h7Q+3V6M7W
SruYuRH7TQWEAv9FBO62Yw65BSrMqF/47AFmE4Qzppnaq/iXtEZnHuuVi60KPWa5hQFV5ts79X+n
MMhUtvimtLCtGtgcHOgOytouf2N+2RsAf+cH4/JVN11NMieo58waX5Yc7ZyvBRS/syFR1Kl44jIl
yt3bW5RR0WQP7kPEiTA5QbX1PKUFxuWEnwITOHTLD8X69AV8EdlXrzOYFSB9ZA7kwU+vk2noY0cq
AsLPxnP7ZWrmdWC/IHFbEOrA0pbODovGEEIQQko3XocLSrex/5fr0rTdmydeAdrC6WcI+vDzAuRh
ifytT2wWc+6RdsbqY8yVNkKzZvtOOdWbvf3p6r8DZJ9Xxp2lQWRK338s65ub8rHIGaeVwkm3QvxB
iITsuzWQlY017EEtoEuuBYNwUaAwg5iIKyK+6DE34MUeJQzAqb9AunPXD9QYIYkCuIr+M0zlweNQ
b9xvP4UowYPLVZ1X28OEmBiiD2Iua4NL2ntOwMd1B5YE9KHkjy+FKwQCitzWy/WRr3AUptEt263m
tGx6QXNpY/PPWSL9EhvHs3qYNUbrnUUPVbqF6zPL2xVhPg+s537Zvsa27+LQYcxgnVAkCIxrizMK
U6YubatooDFXl/iHB3yfmsGx5KNn1qybYMpf9b7KpfOOamqcOKH9oWoO3+BGVld4lE6FEy8/jmYx
umYPEbjLEz8iZKiTMliMxbBM5SzsHtXKi5Ddyg7Y4YxakS9v8PxXT+5rnoS4IFvSSEVlgV8aiXZ1
h4c79Qv/Ld/58VJdXcOjWpd5afEi/DYbAnbOPHPKkECrkfdJrJwDqSmEs/PHzyc7DsGz9FfBZIn9
BjlEY3mt4dgl1RgSzt8g8G5vQq31MuX6WwMoiPM6rXFiOgIWlFk1p+5Ge/E2wf+uI+wKpjaFqTRb
6c67vEA09Yk3Tpt6fBRO1t4Hfj7gN17puAA4WCN9+RKKfTI4yZ7dGflMMhSlvc/ZIwNscdAcTxEo
iDdBi8u3NYPfYaDXEQfxRgWMMpcmzPelecjq4oSmrqyK7U0jodrf7pDRpiWYt9bAiweHAJ4H0tVZ
hlIN53MpvJF9bkijiqGw+MZSkaimIJwDSQPnxB3rNTqNXmwfWL4GIbpIwlPsN41PhE+H0SIjbtC2
m/feoq3rnmXl2b7+KMOgFnKKC6gMgXPbOkg7UPjDHV69XQh6U/pl2H+ucY+7rQqFvuxUSwdlgJH3
yChC7YptrU+IPXAoK4nKGKAcepNowInCeTerWnuKlWLTK06TMEpTVWRT7K+IW9cH7La1PJH3ETFR
iv15g3XxnidNAqcwnia8FzZxTSuehNLDJ8YSD6DF1Ppj+BI2cHtv64qJD3ST42GtsvulkCa1ZoE+
aVwnYhRYa2dtQw8K1mqSHbY8HFqFTSSQRiRWfalRO0PZes1p2CJMqG3bJpxq9jqGMqESYFbuBsXp
b8wMB6OVg91QOKQXUYRRqZZ/fIQkXwZGNjMGSLbE3kNAytcYtK97BJZUgjzKEIWUh4fpoPIjl5hL
k4gG9YBp4VB1u25zzo2Sz6b3326TdV+7TtrCOua933EzoVwP/oiLDuIRahewqkijgL0zRzni3MLO
NKpnaOjgYrTePD9nlyUnHRjRnnHenZpHRLYk5iPZ24/hntf07S98lakY4oGaNBcFXrcS2HIKb8bZ
0AftqIjzU3ZULLRSqWo5HcJhA7qjFFaCWS66hLZSHWUVvL3MdiFsEBBtOX/ht6v7w2Oi/k0K0quB
FqWpKsocJRpiD6bSGz/nC3nG4IK2d6zMSRZCoxwkpAkIG5R/Tl2KqhiwXNYBwZFNHI1giJIpaUXw
dTw58LsKEFy1/7GNacxszXJdI7inpm4qhOHWwMT5EAamublVEHH+nPgfTX2jVoGuOFDGXrdr6oYH
WmAanJ49F3kgutexR2qiF/+NLOJy4MJ0S+jxpaRSfptM9+TYaiS4wRwAJPG82eIL5rE5zJbwzaeS
OD5v3hZUf4B+uq2YiMNkAVyTd/IaP4wcvg6W21jthf8y23HniIaZk4HTpgJoz4qBXs8sU3NbgI8w
2p9Z2+6qI2q+V/O78txJoX38IDg5ZRJHkmHf5lEq07zdBgRVaOl1HpiFuacTovgS5rv23CHh5l+3
jjhCG9E4myq0l9PYY/6gJIR1/85guEskpFyZd6SpAAvsktf7I/Bn+IQGC8YdwAIQA3I8U5DOn8Bg
gE4qvG5VP/Fngt/Y4KPTPBBgjMsaUXfdgfzcrF1NPbScVb6cPOSFx3M7s2mwKXdiDiGXnZ5ZXW2L
UGjH9BXzZPpD2RSyS0vvOf7JRGEmyXwkyBCkuhMn58mLOyDUg8N5Lqs+xc4ubMIOzAScrAtRGX6c
vZ8HfrtYCqCFuxgTFTZW/IlPQqKLdPD3hd2xAgVVnRbtrCxJxxlGaDO9vUJLd1hnSNUySY2SSgi3
FOj0gOSHucw4T+2uDv7lo/fmh0b0/dO7L9Za3bs4xXKnnUxczuzLwkYP9JXgs9nULWwq09WD909c
c6Lx7RlhppvYsGg2FX6YFA9Lp9SN5DvoXSFTVseZ+iZqUN78hn+lqRxgZ1Lpcu5Ex6EHbx1Ptk5Y
u4INM9ZnQQhHiMSihHELTxo26u2WfwcBaI2xHGbAGfK2eivILuY/rd3lJkCipTxGfma9XF74PQi0
z8A8Ot+D9cduvX5JiUmLKvPu4mz3NJysBhmb7u8uI0XoKKKl822dpYe0wBJ2+uZVJwUVSK1764ok
4u74STs6CegpQ6LqDu9B5t46IY+oMgugCOCxwwxjNi5Zz4/WsewDkmPkW1JdiUO61u9iOJiji1xP
fEkZ/cruLi+2F0NtBHl5FvOTawJEC9fMdH4pFp8cLYVoIySJm8M0f9CqYTqauw8ZJKYdWltk2f+b
aXMjUjKPlZZBvVH/DpwG9s7mbf6TDKol6OmnIJaLgTuWnoKkAtKQQ+W3GwvMC47LCHeHAc3Ks1Mh
LIQ+JYlmCZh4siF7N4DsjjsvIgTa5wqlWFwn0ba4BNw6UebLSbQcQCCm1Imp0IaopBAtaZ+772sR
GDNZ2AJUl/0UGDO1V/PLbeNWkFniULor1Z9akgk2udYevB9v/e8/3k/LQU5ZCfJ1wWvQqWDmjQ9X
BXF82ojrLbLD+aPzsQsi6j2jHlClsqQgmRpk+APNyU+UcTdVPi8iBFQj0/H69UFrYSJGciq4RxzL
pwn+RlOt3Nz8wssA00SsvGBWvIrPe1W/QxL50JbtJdRGa3W8BW9JLTN9jzzZ0dZyPjWDneL9I+YT
C/FVLoblHB7CmoGAfGle35C5deW6c6AB9lshimUuxXk19p0OgDCppvA4S8MJ+r6KOlKXuXq321ex
rXLsNByx2L+ZC/UE2kPmyD6CV0xmopzaN8b6rpEY8XizIjqu+Jcq2iUv2aXhE5FWz8xt8eQpW/CQ
ZIUKpKoJQ1GmsB/sMMxwvlN2AIYj0Ll6hYjJjZpN0iE4Ed0hSfUJqIRFr3tNKyZLqlMlu+X0HgWM
NRm4BHbx9qqExPlb4YHK2tD4m7PK1SXr8qWoZ3ZpNAomS0xxvsXuBhGR/d1cWxGH8KHl5F8EdtNn
KwUKkNdCs+T1Iiliso1ejCo+NFKiRPwNLu5ewqwl2fFh3vwhN40y+xEyN9Bg4qSCl+oexTpLJTZI
8H41eTp5KIkmvh1zJpjBdHYEyoqCnMxq7vTYw6ubVKbDziV2hRwvrRaQykQDUMroO13dlicGz6dI
uNv+Y0NeRQbQ9sDCUROpC0kJ/njmN1Pb6bBORVKjB4zWzOX+SbnA20L152w7YlPiSZDnhhP8zoqi
+peCujLefHHfSGP24UXrNAf/YEAcV8JZvkgUh87QTMrSAOJ/y3TLNXWrQXwR+CB5wkQ08UpZlLHS
M+RMOphRbIzxGexIkXecUddZmjLF5Po5CoBhG2AcgpA2AZHsqc2jj8Y6UtI9rWhBHKKXtqE7lMnd
HbD+GvuOYDIW2YFxwfWxMx7Ecy+OVQE+izQDhoLByVPvZjHEAcltE4Ojiq7P92ls/brd+YELuWYT
bV34SylPZ0OQwFz1n5dzYbYom7x07kNwdJvS3JgEIAQReo6NAkMaYL29Aj+edJijDZGFzlKN2gr2
RNwXpMiooq8k/ARIZSZxXQEv0zHkHmuLknd5tYC9/PkdD7MQVFzl5dIPQ5DjLsh4eohZHjtIZR2t
BvyqHe9cwNABEl/qDTx5TOeo9mq/r5XIQWm1spl2+D/28pDchy8xkykahqxj+/engV/6q7iw838E
XeW4JvXUGpVMCcAtBQiFxSdge0y71MlzMPwjPAlCafuBfKeTzIr2SMuWARTllFDE8GbXAPzQY1Yd
qWroUM9/WLdVyf107HkVI+I2C84bBztXWhejRWoSOwFVCP1Eayg1tsORGURnx4HBoDyzt4sZybLZ
A+uSuGG2xH001gQqJIcaLs2MBbY1ijNrPn34Wwr3Ica1OnwIC0M3iXJgOzsLE8Z2uAdhCoavT7gx
RMGDdyCzlbeUoOqiXS8eEowoY3yDOwyti3JMaUhCgQMIv0NWdPAsX59J51J+CDiJfoam00jbcq75
+42APb5UtMmNhnWjrLv9Tj62nqI/0TQtwv+T0IgXkpj2K3XAt4cZMvYqfak5aA/HbRdzpGNb93mj
E5DSCrrM35o2EDrl09D5wBUG6gP0uNTJf44nHikC53jwLoBUiFAXQXN6I0/NVycUbvh14HvVr0Sp
MgCq5fTIAJZzbMBK+abi9oEYJH/sixH/Uf2i1fzNuxCwgHycYXu/Es3P586Uf5dz9Kn9ylfmzcNE
x+0lBpnL9xD/eE9UhrtWvZ4iQlxBm+qhGnwArjIaVfTQ06T166I/fpL+LyiZccoKB3vhZAXSlIkJ
Oaeos5I7SnV/Jt+fii6VGlwV42ospGdlHTte1V0vYDt4qvNTUH/hOBsFntiWG2GBQU1u4MvuJthg
btnMK6U+jvnztLzKhruM/nWZsKxZodXODZqGJIVA42bwSsusFUrQHf+kN7LdG6xyb+Rh6rrohkS6
jEHD6iSjcEycBzD0DgFCAydSwaf2ib7LRX0mXIk03FrhLsg3rOozQCmAPUAzS0VUQsYsU7vnp2VI
q6Kp4aA6rbmIIGJ5J1B3w9VnPpUDnOAmG0diruLAHCX02DJYMP1HUrfWuWZoWnDWexGc7fk3MccZ
VtIkcMJAqwbTtXpldtyQg8ShpoaZLnTMvDk/DkZwIp8VYPWq5uIrcUUxG5TEMffirwL032FbANAO
QJ8BB7zvRisZqtm/1VT2lLHdlpNlpL+JgcbZ3WwoOxGkr4pouqMYgdX9iQYGnDjpUGUP0sN5EvdK
VbFUu87cYRyUvNbaTrAYvQo3KUCDDds+nSvPviYNLhc3g/MRrtILBHH7Q3YfcWJLt4IfYkvOwZJj
EtWo/MtJ6rP93UBWXBpwU9vWZFKtoj9P83/yY4OsW4jwt5RksJC6Y0vVKwDTdFKcyF/6pF41Dh37
/H/ECa6C/soIhEtbuqRQGS86tdXPHOwg/Ropg9aoDQqYj1vQ22CQvqEPwJLkVYyur+Pegp1VVm1P
MQqY7XV3EPzd6aQWVzN0/R3JJjOO4GsV5q0Qg+YQG9/NWiWgbr6UYuKzrWqo5PvapISa+HBZGWlH
OvSQt1RH8zpYzpJ52/h0RSkLUHL89I4H54r6ubDqdk80QMqasy6Q2C5yMh9Ne7t3/K7Gl7JouSJw
laSHjvYM69AKTylsqQFKJZWh7Gbwhs4ZHGHyYTTF9i6FgIzmGZtq8bEVWkC0J6fLLXFJAlyjuA3J
8dMw9O2f4HZlX42vooeAMMS/7PWbDE+Z9Iv1zUtw+IkKY264BJgEy1DZ3Wfm0VPHTj0sFXW9nFg5
H3n5ZeR3Yl7k/1/4FVcUnPLCRnx6h8uHHuRVIStVgB1rU3psyWNfmsQIDngyty6xDUSkbc6C2juS
Ss36/JNVNc5yFVjvT9/rAN+hYnJN6PbWotsPUHjFQSH7n+B2PAxd7LEeizxAh+UjMZues13fe5KS
DfBkYBJwolVl4yz3+h6bC8ZAxZdP/Jigp/wo2HSUtpnabF/h+4scrLI+kVqzmBowEU6QtSAZNj2e
CSkKRQ9DSJ2TxC7nl0rWOi8BGIjXcJevVC+d69+AcIBa4Pciss/+jv+8Wkx82XJMZpwhVLGDXs47
fsOSoS19CVR9ExsKVzklrPcDnEq/9jGs9b/HMV59Mn9QvBWzp+mHxpGbSOa8ph1sPFw+Uwf4mq+R
iV1IMf1acGPVRYgriHgGu+oWpUOsZfGaM1ocuenm6rIBNIeOUn0YLBaJeTz857Na/g/LPIEATkx6
jzdlUbn4vA6sAqvRXLA9PZ/Lk9yV02H5AFQ7/0Iw2uuYajDbhPMP2NW2zR8KK1MD87OGoGaO4WP5
a2LFdFpKAGgBxcv2BfZvhk6s5iiH/A+PRM5R6KDpY1vPR2VNU5DrAwZzIN1+va3vE1SwUupv2mSX
yJTlCIaMQ/rj/MWlCCyeoV5aSU0FmI0ZSlxkKFHEx+BXP7kWAObJwOmp0zc0NPr3UNGLACsBaS8r
iiKbTmg3gt6AoEVsxczJkFyOB5jpIW8VL2v2LdI7umHVKu9ncEkvmMu7yK4owetjVA90dLlEH+Sr
MGulr1Vxqlr4I0sqyyS3A1V578AHb8Q5I9ExBrDNcdTqUTUeDYY9XV9lr6zdMHG8gowdCgHCV4pd
C+qqkFyTaJDO6b8OV+YK0OCNoJIU3nZk8WExknpmzLpWfCp815+SvVFFCGZ6Zni6gBKEnO7tY0nD
W/OdGLBHuU58fPuD+EpYCDXL+QqCUOQjjye3yvMghrDeEJnmDF/RwnpP71tl7JT2NJBlNXGQy/T4
1zZVDDELhq/sVtTkUo5pvqcT/h03jeJAfig0iZfTj4yZA+rzYEynxOJ2xkT8e+aMumz4ijn3FLnF
wgpMVD4gs+NMgomJHiC+7n3pb4WNoBslc7SWKaX1kU2p1u4+PW6UPm3xjuwtC8Ysb44VV7JLE2PG
kaiC0WGY3798xlSoN4VWqt6vrPymSi1bdg06vX9bahut2oGcR5opbVigrxVqxN6h9DMOvk65/+cN
R/1xOx42BGOrRAJR9dW6mzcYMEBLY3PdWtI2y/Rm69/FYO1PWnJwovKKn15mqRAKyrBoL9HWXQqt
mjeb3EiooFQ18p+tHQg0c4Lv9EMpoWS5gNHCGe+eOdS9jStpbKKiq4CGR2ZxDh0jkmuzz1LdVK8T
M/S1isenXz3XDGCWPrc2t76ejeA8DqXFLgc0Yps0Yc3LSSqtdJU6vqUttYX1Po4SFq/CVGAt0dG/
vy897rlxgs7BKZRg93Qjzv09oeO9KxUXu+XLPQYx4022CSylbb4pmB3VC8qiFi9KUL8jhVlJqk5V
koYNOm7SplcgLDAWi6CQKw5+MCpSmnd8IMHocw/MrCnllf+9xXiIu6IK6waeZY/zdY3zDWwmmf3m
MF+FAAoPR4dFobLD3GxOKuOIwUnql7QlyxXR8d5yi2v1DFY9XWtGAyM+/LRf0G7BLLkkNtjEfsj2
OXRuy1CzranIFd2+8zT3FNQele8sNGMc23x8ezNnzodH2ON9uQ844IBx97WS73wYUMNcoFwo3uRN
86BpPCY9vdWNozEoxz/+oqyisqLXZZ3z9A3esAIYJ/fasoe0aPM2iM8C+KVkdoaoWMh8cOOXQP/x
Wshv361yS8/eNbha10zPSyDOh61U2HoEfirj4Dcl/7+/dS7048TD8jKJiQcifmQqqApWoRLC/G1i
LLKAqzZ7Glu/Nr146sMpA5shYw3X7uAuw7tjwURlSd0KyTrjlJy5nlouDn7BsqhAKThr7Vf161ic
Q1CHG79uNq13UVNXSIdpLxNFx9Q7QyBJgT+WDJCAUp8QYPiXI9Jh1tbqlG2BbNLRGg/wer0fi++Y
3VlNPxstCU3+WahtiO6AO9TGne4l4GoblVFOv5oHkIe8zyUeVceoEVrMIY0yCzp3+QIvXLJ2SSqo
HJEdbszR1nxf1BZMjufAmTeHvL6un0pBMCiL5CNiDDRMYPOmkawatMwLxfAGLI5qFzVmPY8i+QmO
Hl+u+iNCqMbxKfF3brn8NkAqett3pVxGo18723A+N6KRaLTyzORTslItcsKHAwo4gPGf5LjxvwTF
KsSVt7oirNpYlPt8VKZ7Itjk08Fw2s1ZDBpF8xGna0WPjoSPjCMmJtcaSw0/LmADabEvloD9sqyQ
KKkEXbzlMxytPdz9qNygPoXKnvgDUX8LsxSvPQTKU124WPPqTlZlGdOWHMyvWAa2Hue7sdDg+EHl
eypMNcI40zuqY4L0uiL3rxIoHYZEIg/QVTcqGIHdd7viJSyls4K4d85q05/LE1WRnL7OK4HxYcPh
il7BEOBabQ7Ljz/8PdAEhe/d2H7YAWy2sRgIl8UfK5j979P2G6Ier2rynNjYTa+1PNGYEePmj3+S
kJeq1kP1qv0yXRC0keenhIcArSSWER0qrdmzCzdjRMmK+XFVq0ByVsCqwodfcsrjS0FLjkix+V81
8AN0zjGx4irdjuuYG9LdkEWnW+fo9ci13crDYTUw+cM5s0RHl5C2BlJTaQbJUQ4/ylaYG3QlFb5m
HDTldQjUq3kr9xgTrchguEtuXjQNB5uEwktAnV3KII2MMTQotf5Cja0FWpAj6BW47FsuP4ZXZKiK
4gyONVuAwNEYTiGF8Vh6gtssNxajA2Usbbt1NjXtNmUFJOG/PPrJiJHdCe8aoT6McdJ9RizCyOfj
k42Qsse2N6CbcTDdDFvvb8uZRB2GgkVWpcNYCWtUItubbb6VrhE7HuicgYVODiL+bOYdcnQv7y/s
BLieRFbLEox6ikkLCEVVlJD+3q1mHgl3E25JjTYET95lztnq0GVRj5kHG+fkbufAbQARd/dJ9xJW
cRmdnW7ZICjEHtNBhmBrRtuvzYC1jbuSlTyVcbz050c6VhZbOBsI4B71X6hNEkROReNwNh9M8zQN
BOogwc3IlVM/HZudqKeZYgxgbs/3RirxMv5OesgzJycdwfKQw8I9R8Qz4htFfrMqKxuHcmeyypC8
s4y1cEj/wEPKdy501pb6yclmisPBg02+D5RT7Gg63IU4Kld9Y696ui4CP2zNKYLd1e7FY3lKAloi
kY8dXuMMyUimo8lvoePFUzSB5kFQ/tgw+SxBjXlVwZVg2PvJrnydfYPxXy7mjA6p+TNRwSGTLMJL
TWGfGzCWpMd0fte4QfMovl+UW8nxRUrCNQ2aLfLNdPVmlHzxTkRO0dk5Wh4r3U66XVLXq/xEnM6h
ZjnbNkf4oKpOwwckXuEtmItFyZxP/FE2ESVRgltWtqp0BXJwMLTCsI/S/rZDtLzJ1cXUKG/u5y2l
ezwChMrpM6eLZLzvjQA50T+8LYiDYBhElpSBm31Pzj2uXDxGDC71dGEd6AP9oka9tGnR7bV24xQl
mR+17v0t5wusjQ66xi824r5DYGZR+Dxzgv98tMHu+7vwiBUuk0Iyo1Y7u4V7V0kGEOLahLxoDiPA
Gm0XOPtVNSUoq79kwiOc/mPoCPeN7TDR8K5U5ygOp8xruGTZULlg1Re03v9Kwxu93kFXxxNMbuN7
BrKpHH4QcVqbFF2K17FHYIreteDA2GUtxBzodj9JSW9/fXD7hkBYWs0J/N4etp7MN2/aQdwgJguW
BMgfHpcn/Qwklruk1pw2jirppwh8hHOMwvnnY5p4rW9bquS3KZ2OE932K4D7ltWp4Ug9Cj8bk+Z8
Fh6hPtiYw8NuMQ42roQCnX5V7uuSEIj23AQKIggpapwkSveQswTROuSS3kj27TOGzurnLLCTgeYy
s3J4bu260U1C91Uc7YVplRVTI3zxg2CG67XlmULItO9KKbUVsckZIhYfBXWP5DBiq7x+mxzeieX9
y3dVeaS1G2tRiUpDcEdk6hQ0Y+ylgkzQ1aXk5+mq+aPqPDR45kMaPh3CzOwm0vNqmCdPP+HUoz99
oiY0BiSDI1CCAre7QTlbMdZCRHa6EeS76qEDkdc7Zdx0jRpmQhnkcCVXb8Mmhub4+M4U0uo1NYBl
MF+l0KYcn9fw4LrR3XpO+WQUGJNAVGNaq4fTCUiV83mIQwmfDnl3Ohh1+43Mhlw58FPPUeivDjKa
UgS62DLHwhwrt1GAES+An56dNXk6JMWteUYbxSAohvBfpIql7g+/8wcwQrylCbPeFhF9zMWiQE2z
dXVNOVjSijES13NVstV1PXAUucJQxISs3ApWXKi6b9jQyylla4myDDtHzwQKBB43X6EFVSe0L3gG
1jfMhdDCyMF9BBlS41p0v95xXL8s7YwfJ+bE89QAVUai9YJyXH2oHp47XjMeW6bUV1XftqgCRmKy
6sdfutL6H5SHqjjfgpHCghL8WSG60o4ZEnsz+JitLa6O9EM5qCTugOv3vT4NBg5uAwN6Fb5Wxe/L
X2pWJCOIDb6bY8S+EmsPK8tOZbzqxECvXgs3Lkqj162Q8jLZYATL7IRI7gmiMLPvYGujnkX44yIL
ZyxqGVFP9iVSffuniC2mORMjtogiM31KadRccBWB+4rYuZnJEUa92iphXK8oHXARayk1/UexxiT0
5Rpd2IAHJY3DBipYDm9pnoqNurqEVVnb4vSp7+AYC113/7GokwC82NZdDbpm3dVSHLy5RflDWsN1
XXLmZpLuV4Quci5RmAw0hyHVlhp1V6Rb6FMWGWxa4k9buTBcDumsiUCDyiBz8P5SWaqj2h2F5SOB
q0t1LBYJ4kyUGPSF4viy8t0nK9VIEP0JHSYkr3JOtBIwTwaSTZw0uFh3w2qO59NUyJa39GWbg1Rh
DRUR2pGhPkQi11V9/tPD1Qzd0hwhFU1yUGwFVMHonc7dklbgGLTdtX5/8nkQtIduXwhsKvdC0S8A
Sm/PHELe+Ns9R2QTxvwZ7P2vjUZqQD/c4vDvUldQeXhLKGJ7H/nArIip5AZbM+FlMIS6lsPljBfy
9uuJc2bHkAQXAo5s4zxX2IQgmERmwnwRHgffZb8j0VEj8V35q36fwJ67hMsG3Gv1x458AqmR21Nm
pX+gdIUCo1kWfiMx+vD9K26G3DtfgARoRGRy5WVnSbJ9NvS+fH3e+OkMHJkvLiNMOwx0BoG1b4AY
+EVTsy9sx0EVIv4dRmCwuDtvRp145GI1ZjOECs68T+c/ogRtMVflvIO+Kw2mRAdLWcS31nEkhA1e
FTMnPJ3JuRo97t8omNXveT9dEc33AX99ig09yreH1ZXec8GtPJccOFG5QTKREOwYFZmvyoJ8/Mxg
7TQUvRaqlNChh7uCsr9WL50Lw0zItcDXKKRMieMgDqagIxMMO7mA/biusQBjj8G2bx6Woszg3Y73
tM4R+338ApCYq2NUB59sLAzxNe5AYwzkt+VUKWfVOcrkGRkQHnebYV/3f2WTpdMSmZ4ZkD+vUgsS
/W5ozN5nwoVmDWLVvgCujGG32ctOuaHbDvL3cEWfP45g0/tSQjo6Ji1w8J8t2Wtv0n05Wd24wH+b
4Ag5mB9wwhglzeJbk8IDRu5QifV+l4cVM97PG4TprqlRWqY8gpwFujpLygAGJjDdZCQoVC36wEnS
gNDMntdJ8c/x7xKmLhLWuv7wrsJBK4MgusuFx0Tv3h2NdJ+qPnG19u4QM0PHEJFPAcZJH+vJmHbb
9v1tIbgtXxB2Y01684KBOjGBItvLEDX2PUwvRctTPTzPJsHlCGuUSvy9RVxGCltqg0YCEMrKpdez
KH71eIZIdoXvOd/OtKHgSkWgBDY6/Rez04Gqeo9Q5rwjhSkg+QA9EeHMyOneblbARo3pLbxahVnr
sLjxciySTOvfpzsqa9XBKwugoiH2t+NGNo7CwOXjWHAS1k5EbhupFM2i0nSSuVWy7SGFoRdtvNsZ
Ij4yQtld21pfcvl8emPl6iCUZsfilZqlAqhi1oMr1oPdmI0TnYqGeXu3Ieqer7ibqcH0n0yNWUTX
c/pSlysdsQNEHFeZAjA+7SaFKPShLl8vqIpML83Z8IU4ydc5wEWGGED83B/HRX5TJ1H6Mzez9WGJ
Hg3Rk+SFUwBRYHs8PDVjyWmfyLpCe/zNNeO186FOkDmnhh26qV431iFVo7qjH3szQVyW/XZkmEGD
rlN93gcXeh5yTX499GHSEnByzZfZhYMRcbmO0KChQJkvUm/zfCUC4nnCJX/dRKk0ZHQ5FCVjcMpz
8G0IqUwkX85JH9Tn9pVdXwSFPYljlcPPWpq9yrqlZAcgJR7/eLPKDEnMREWyPI0i9yJEeARbSm4M
gP9tfJbseO33rwqIkq1wNWqc1HhPO6mUj+CUSLRqwRthpYkjo1cwrtAf/kWSMgqOqZ3tWu/fQvHb
7NampVnme9m5fAQjuY8f2sV8Xw36wEXiNbSEGFWx8hd6HpqF0ozLbuQ2GWXM/MFbS8PJq+14M+c2
Zmp8IbiS8nhgiNx5OZH8UBAMLLSl8AtATmPIcT+xLgDgFDnxjkZ9uoA+F41RbbHJdt+M836XLgL8
kGt3qvn4ny55fzco0dipNXrjh8qyM4fm2MNw5jxYqtHDdnFY1UcXWd95g17cTvNjTIjgjYuuUXXq
74UL0RU6slOKXkOrRhsTlwtsonL3b7pHtJIj9fHh+OT+MWojS/j1bnneSXY+CuRlt3EB2AHIkkTa
bUaR5HbFeLL3ALKMn9qvNsuph3ZPUBlwHigvhl35TgvimwJf1C90Ul+oLlhDqRswBvpfGBwwA4hX
cgNtkYozq6MTNxVq4oT0nh0ke8pKFgpszzcyCFzxo2OM3Pl4n/oJEx1q8uGkCuwk0pdCz4teiVSH
Dn6RERGNx/4D088RALYon1qnjeBYjGFVqs/QvAsUKFwTUya3f2PSlon44D+k7AVogeirnOBPQtm0
qx35e/KmNNOYOJuBwDnH+4a92j/G/RoomQOh3ngFOBcLQ7ccBUh7JM+19M5RSgAWkPAcQqMq6Aa+
Pnm8Cb3+756/vSNcjbVPXTkcKC9VsElsAJ8RmNQ/fzxVch/F26yDVe+V55gGBFeb6GcpoM4+6+oK
HDQCqk64ci13MXJM0Wft8I7KB61xPyVZVYqwne06nDr6Xfyvr8vlotBO2AyErGGZ4R3XJecj9OIS
H71JIo0aHBIbctCYhCZaWdSXj+xg7mQ56Yg1DJijuzqhtaHONvENmIhppnZagxXfeIxZk6fWwspD
r1FhB0RfTF0I9eUEEzNdk4zaQ9l4zT3VVuNV/Bczum4kvOEKnYUekF+WMmVEYVSafNAboe3A7ZJ2
nFKl3R7UI52D3uJNVT0wDhAH1l1oppp0EOUwLKDTLVeZpeHQ2oyHnqfzibjXGDwz6D5G4lPMG+bn
tyU6QqKzNSO2J2CfbrimwdZOL81odjXxpYUvDWR2SEnKtBht2Dp+3yBpvbNCSfFw2MIdpSYTDX2A
ujIbciC44jD3f5NqqqtUMVV7T8lyUb1qqP60ASv0SVljv1SQEBBVQeX2f2o51t1CW5Kh9oV5KAQg
uql4eAZHzEbCRk76u5VO8dMRj0INkYcrC38aTUXv78trct8d1ys0vmk6Lq6GWW5E+1tBEzucZb1x
Q1e6uvaNTGb/ikaTkgRMKIrilvcswRU+nrZ1RlOpKnJid+iXfS3fQUfBBCA9cws1nsBPT/3qzzlK
tIg3+ZGRwZC7PgHuifjLs21jesBPXt6pIzdOtYk8YqeAzUPbUt5hEP5CzIcg1SmFuG/vNr31JXxO
KPYww7wAaLCNdPfM/fn9SAMwB4nyZgGOLlbxN5FPMzGIgX37kDYCMfMkwkH3crU5GSB3e4tkOgFf
M4x3WV53LoJd2kAwcigIpmq67RIC2dSbG6JMukGTRI9r0eszRqRjGjP2bj6MDwtrdoqCIqGjz+Q9
6wfGmJ1PrGcORynjSkJvaGkb02eiIN6uMMOkfn+mu6ylIUVL3CskzNG7f616SD2Qvq9P0ltTSC0d
YCcC3Uo610F0r7fVIzx4yQMsZig0B8yUwsWDZHzlt1lSk82OoZLZwCGYd2OAMHnZEp2HESKNQKYB
37j1h0agTeYSM7KlLH0/zbEasktuzAHacqTFpbgirHIz5zLpczSV8k2spKlOX1yNsVYMgoavGg6Y
/AYvA2bsHKzVqihORSH39Gq6YEjzb59w816e1lIS+/kML2F0B+XJzMPjmWMD7o3Yo7+PkY8TdKoS
hCgdnw2Ji9/tdcqkTnCRV5DPxvkSprNNtQ0S0WdJ4AYmwA8yo/i00uNFZ/NUdVFkNMjR9mnjXOGZ
MGcYIu1fs3x4Ugz98RIIn9wz+mC7womUvImDY7v4DSDpXSXHKAFsjRYW2PzcXtHZhCwvhRh5V5M+
6rwru7aJiFGXtEsyWLUVpyB6t4IaGxrhg7yPrgPjzVmv6tyU56KmqqhRgsVzyUW+KzbygLHD/GPH
6KqZSF7cJUfrmGLj4qmulLBgKKX2BokC0HmVSLfF0945zBJ6QetlQa9+NVJYyPZVLQ41aDnwIX73
F1lts9Bze/epix/5Kd8Blc5zgR/o/5GBjjYXDChCwUBtS2MpB+NHkKM7R0ZfqmGOJO+lsOZfD/KE
vbuCFUVbZHa3+hHcyJGyYVEs1zdIMsE+6vucBwes4G/vhk87Sr3Y2UIoVdfQYeFEl85ZmytcE4/l
m7QpwCFM9fgffSmp3+qWsmkxmYwAfsa+ESY98rlGqbyWJRufexX/A58yLQ8t1gYLrIoFw/cpSHka
+7/S9wumaZ9yMnlIZZAxdped6atNVK22efHktyLz0z0N22mLOs/dh8F4+NkLq74Thax/YrxJwgSO
47NXVFjP+/bVpakSc+g9/Yugk88R+eAylvoOfay3uz0jXiJZSeEwGwqodUahygJKC4sY/m3OU5N5
S53dDzQcWXhE3tqFRnqNCuyl+n117LyepOL5xX7GZkUDg+j3xrJNZgAF9ZvhlkXVzKGxW1kPC/Ac
6GcKz3aOeOwRsMXiYAwKQm6YvYyAGOSWwVZTqo8UVfa0mXNn2EwlLIVK3PFQ08XrLuPTaAzKHrsG
Q5UbJOq1yulF2fBf9SDrYc/qokzJGh4SCZZ7imZL0wakwSxIAZ5cY7jJShgLPP4OKgEKhQLYe2/J
lKpZCWrIi1/V6cC140Le9eZsT4yJUTzbUAJpxjSTo6b38TYR7Rq0Wdj2WKjTPdB6hU/IVQjmBclZ
2dFb5MT7+km8Dncedm8F1cWTc++GTZJojJGfKut9Id8xblGi7Nr1NpEolGxEJvd3Dh+isNE6EonI
o8XPLo9bedUdrInoJAyopoMHEP2rzFRMQxRWfaEF3/g8PlYxgdwRsNo9BHHqFsS32JbXvNbO8qUi
rKiUTOpem3klDtksqc8BECimPphVts9KhfyYginx+xR9/AHXU7PgTWIrWE50HspiJp8anIkNxomF
eIyNun+Ip+5IhntkoRE44XbVEvz1Qvh9JykBdeCEhTD5XzBrRio1bAlwWdv3R1fgeVG1eG9NxMwO
cOGeMe/as0zqI70/vRJqjjNVQTU7hHEuejg20ZArGvkYaUnq+zW9BF6astQd14ijvnqUJzGgkPaq
BaLVlNUEAqMDPPj50WxoUus/zG8nnKVYPZxuEjdZ1BNqRCe+1C31bVBtMFi+wXEQPoHU4g/1bX0M
J3KdaGA9KaBz38Y+lwFBCVrulwU1dkc5R9lR0RiYKI5dFnWmbJkahy5FXSniya+lQr1PKpPAN/5z
OvzZoWk9A+wqmQk+aQhzRCb6qCLHT2nZ/jlttLvOG3QJL3P/MNBQbOtL+62bpQrqVLrFnlZZvRSu
SJwemPG8JVBILYJvlLWKGzDl3L09vCHbrhnPe19zGtzxWYsymS4QqAmbyTa+dOgluWgNZLc4Rljs
OUJIwyZroVrpWXKLOBjvUPj3dm7XBndmeZqCSdNak3YnZMu9DFrgltfx6aiHNoGiJMk/qwNsxskj
tPLRm7Vnf6IwgY1UnTLlvxzYjMB9S5z5uYzLU216BFk3TEBm45xMgOe6mY8xTYjXqA7Yt2FOG90x
p6uiGdu5Bmy63Z2pGDrOjgugWHNWkC+oEjDP+AQ5wBHtaf+bWG+zXQAB9+RmEbJKe+EiBV6W4Xw9
bgPdaxjT+og8aYyRUypB2D2Jh9dfTz+ajmC2ggzckUcFnmSy/EM1qVlV7r6qylHGoleEsSjCQRjG
jQmvOGtcJlJKD540PgwdWvX4hfuWgsZu+EB5C8LO19X5TsiK+0PH/jAMWtbHJhALoIegPnY6smPq
nSS1adEdI0MHzkhCSg0MP4mGhyUahGE0mDsWo543aOh/NRT82T1pdGTysT7bd0sgTbP6iYtHuQ2S
3ucKUFdNyedEFdDwKRDS28Ou65G0Bbgw2zPiIBFwx+l7v7s437Z1i3sjHNcDc9vIIhROT0dI4G17
gdJ/cPBqZJJfABekNWa4Tj5MdXtFIOB+DGnPcdGirf6Tn5BT1/Dc/jrvtoTD2D2DDaVFWaVb3P25
KcTQAJNa4XsDiL2Ytofq9vRB80tpCsPRh4EcC3V3n7Kx3D86MtrcWwmBwwT88eFb8QU0l+GWTbFq
59yuI5ixr4CKy1Zx4zju5jq5TKrO4gihtxlQ2vUhr/16zwJsNHUDR77kooTl37dNg+szkuHNNAvS
jgQCGWx/dJ2zCfmpzRo7Mi70gxQUODKj5ayvmYGRyTH1EWE6CCSsn8pW1y4JxkK4E3XsBb6YJU7g
MV/YcdB7GPFTn2enGK/aJmVm/zfpQP+EPZvqETRlk4n7fFwK5SQpkQ+YtNvBm0Qj/a5WTGhgPsCb
tuh14RhWeloiyngVIKxc5b0Et3pt4JD/4faUqUkeC60AzTfqBF0pgMM4C3HNp0eOBtYhWhBRjL1I
5zZznqArguZwXY5Zp+dUD0jQvAqAnj7E36IyeCrRCj62Ogh0hDWrW0cbSMt8j401rWNcgWAgcwFu
8vyWVUGEgC5s22rDXYr7s0VDN5VdKRLjXg3qFHPZwSOC1RzTHuKVt5jcH9Uq+5gdBsjly1WNrbQS
0PcJGJRlga19qHa7gxTscHgTSb6/FvOSvSo57vL9aPqQxsUBjQabBbgebxE+cmwSkRSrT7N5t7ez
SzahGhfw90vMV68cjoCjvpTu89AoDeve5hCXOOVQr1CN9ULGatSfOkvc8W38l3aa8u9lQipUDKIN
rb/X1jCd3P+B3K8dg3rTEWeqJY0kbL8bx7YflYNluF3/IKwlTc0qbThs7XNLf19ELVEtTPO7lVGz
Az0yZI/eQtiv799ycmnb6ZVM5WZ4o0X3zzFIhcklo/7qxdT0BCO8Ha1fEhRnktxGeh74QGaGIwRa
dNclJqFyKQBPr8hpaHJhsHrR58ziPU4YrOTHlU8lLEqKTDTiB209Occa+VEr9CtXXgtwJX/HTs/U
VTWnGpRHw6XCmbw8z9v0QgTTqoGt5G6cOVkwkU6gTiHglJ4ZPGwDZ8go9/tQKiLxuS5Nm/TZxPZr
HJkJ0r1oxRycRXgS4Dokd74OngDAb/NuCVG6Wuv2LqMpHuZSbuxD7lMiGr8iX1S4ADcama55sAS7
2B9wN/R7F7k5cccEYRJ6/TJRGgnjcfnM7mg/vrW8FyRB+2aAKfN5A/416OwV2u4tjEqUqBbUS745
VRTCQLvYSwkdRNUwjiadvd3y8Lg6+zc36fx1LqfAHhfTgJQjLCRg9pFvAwVx7OrYrSzzBw8oi/Mg
6WkNT7un3idgc7Y7fSywQDwznl7HPex1DvzHjmKzJdjqGD8LDIfnGkiWBHlRKcQPTy97wWJbwzfT
xOYMW8nVPMPYvO5MnY8ga0diPHYqPJW0vidfTsRKymt0S9TiL3itFCAa0s6qFrcy/W5Orw6Fd+ZF
wNiNk/uzi6ikpohlkV1P1X6n5fRJy84dJOkO2fSDVHoPbQssTFSlIkIGPHIFTO2FgGykiN/fCoy0
MP9jYbrrccorkCpY9lglPJEWGwosDSlhgUtD/z3O3FU8AxuuYHHerwgfH6CjP9vmA6zxXj1LZxjm
ydFbTM7LDABQZYgOpvFtsdZ9eU4p8A6kqp+leZAjpLX4e+XIIZ35VkhF8l3IY4dQoZTK/WVrPc/Y
JV8lyNvj/8QAHR4vJfXNDLYtuEKym9eJwrDWi4fVHEPSkgkq+MwJBpyNU+N4wT25u8DR+RZMcx58
aqD+HX1ZVXEwpp5kb2ONasGVfoj0IY6MN60qJHJK0DLNpf9BXoDgFlHVSSYNcRR186Ykci0rEhxT
JXLyfbSjui9xbRxZMbANnMIRvJHQY0JkBfjgkpVLCBIZbqgQXlD9SHq+BcCRSe0k1xrIP6DMYFtm
hRpR4IjZr5RXFcVk0GQkE5bGV21+krweSU5jo+qWfjdQUdWbbxzPnQ1m/Szw6aiy2frkPN+KsszN
O4k8V8qcfAfWqLTf5zzD51s7uB0RgGpbOPcX4tYdivQWIj7lPi4UYc0fFy1gdmiPpsvXpSBZw4lg
TaAHo5EL14zSAr0W+OBQcoG2HN1+nSmMW8sktfhIErooAPFPRZH/SxJJjyi9TIteE4xUw2O2/S0p
kG4V/q4RZ+p5iZUfSUnoz+lVxhzmb+OvNcxyqg7v6TDu2Mcv9BUM4BeS8vQiIZoco1lFxzW6qH/s
n9Lgiz0WKZXhNMAWGrs4g2yk+Njs/lqeksOYgV6EDiz/NEERVk6e2nZXPAln9cummIbEhh35DTva
7C8ixC9RnHAos7zLMzqhSHYzILzmeE1qn9KmkvjTLwuomsHCdxFOLXkCChaYwvU0fhLbHW1S356m
pClHdw83PKPFTvLLVQTcJV28UKPgoC2MFHW5yF/hG2VSbmh4kTaSlPcZAD7+fHDWfKMqn8wFeP8R
Uz3q3sypzKTuJ/M2bNEQJ9Oi3rUa68IZfQzrMKxNlNydSIew35gDHdYF6nIwHIxSVeT3N++BvSV5
86BWA27dDHziBxJdiJE4SwN2J9Al605bDd0Ac3hETuGE0VrwM5HyeGG6Yd1HNCZPgonZh5gqomBX
H/LM4aQU2AD4rZg2kMPUqMFYE8jcAuqlwNHKgrtSThLFjh15IxEKCzg9KmbaqCQ81jVHyJQ9Umwx
y32xP3h2sc6uqbU/UQ37chGv2GKM287KRBAQG6tQbngzKVMWSCPWest96VcmhYcPn1m3grjuGUqZ
xIvBj0UXJ5Swr0Ce2TP6ES4Nk560EGJK69lm5W/YfSAWE7ZOwRnLRvCVDYzYHHaRUqred9LMIB4h
jXHy7q3gMTuGk2TRgBhg3fB2jb0Qlp5uI8IP5O24s6L2m5rERQPydU0KiijSVpCLPvSPQXA+ixqS
uAuR/T/xQMOhSD9q1EA5HXzDWVo9MVIuMKeIZtp+hrC6aS2wLmUE+yjx8VfKAzJd9w7xn5Y7arxS
5gJMlQ1rLE6lZ/STbKFlQ/Soynn+CmZO+mVsigTiHD/ooMkX7e1WSaVqGMeOycgGHK/eYdv4Wb7c
mXbeJ5BvZA5QqYHzxqYMRvWfFZOFSyJFam4mwRSHSqVXeyzwopK81BrOAXeRQBkKqg8z8cn/nYcL
vSYH8CIAWxqJvQ0p3+C17/Mr0bLz2iJDYp5rH1zeLBbEVbHOnV6J9VRQn6D+luo0p1x5rPPZpr/7
LAvBrD8pGvk6bjhmVzgcH7388u2OfFqytmvbg/IRB2lpjUhUqsDnnNmnrHl1u+Cu6U1nUX9Lk2kS
q5oYw0eX5CEgoLcjPao9gDXHMLvAtOLZmQKJqxpzBI4+f9w436ARw41JtwF9Vu78s1QMZASzQSI4
irwjAaFqpbHONyCHEpXG5mZNlmZa6XJNhc8Hn5uBmgkxalZjYrgz6XYAhpqBf5xd5w32+3jEbSg5
imDHEYo+lYCdud9IPdphtlAoRPl5N0A0DnMPhEwesLarjJERlTp2Pk1Tu5TvYzt6QIZzZgPUb7Yw
PvOH9dynS4XznlD5z15nQt/sHuSkaez6m1RNDZJ4aHiW273De2h7uf1eQf+5bOrFNxFHdsGvAbtQ
Fpj4Z98GcQVnIaNCRqbwOdwODrQ46clEZxzBWi7JRPdrssiLUojUSHVaizE6l5yuMWl8tWYqWOfR
9faWXu5PvLobC0Wo1wZexdNhwKsGZlHsaEWfAHZPOQAWh97D5yhKHw/U2zywGgQdez2oGdlJMjEk
iIhEV2HyZ450MY9z1xocTDmGo6noY3Qei77fURNvprX2zSPFvs6/A3OixLu1sMHD2NG28OzNVi4H
cmmUFkUQBYD75NbL0/iwWqkljgio6lMCIuzbQJ5KRyQ0ZSZOYmGucjUHP+xk9J+gcjBoH0rOJVQJ
aaD124y1TRZgT6r2I5oZmYq6UGKFXA6E4huYzWMiYcB4f4OZwu2fAHuK7bsDAnkSLpaqF8sNM/EA
487+lPwpbRdIwX4Y0e11jEAhBtHZBBTG2MYKi2UhsIzFtzDzvI3YtZ6GLkm24u2M4N7sVtsLuBwy
SIy/WDUv3TPRxp82hZTO/un1wbTwdP7CRvXjhctUhfEM2PEMMUp4d/4P7eVSDZSW2+yaWz+tl3o1
fwqtPMqi8kyD12T8NVljw+NizXfE4pTfRI1AMdS1NrFJU0I7TuNkOhaQCmLcYnFyfddcqSCaKp/C
8qSCBdFUeSblHvmzu5BI7tAqdnbw4KdB0yGixfQAyCffBvsNXeIVpr/B5IPA2N7d3geHGa6Rggwd
Ao9F9g47lDu8mJ0ULddgHMv4nfO5YvHbe/YiQvZFtL9Z8V00+eKWggBrqa5xg/Qi/kg12M51zmcm
By3NCFHZg7vbAdN5xs9M74IYNbSA/fFnXOMC9+1CTAIsW4Cy6Qq6Iw3sj/w8KhNZ9BYHMaILEjka
j91bYPnVs5r2Y2SsqneOpIEVKc664Ge/aWbRGQ/87FidowWoic1JwfOl41QYj/lZ1y3DBHiLNGak
jZK5F6EYVZOKU2xwZzaaKobxQgZlLh212AwtXGrydkREi0Us2SxU0lQASq1yjTlSH1y2BCTlsarZ
tvWMcKreimOfySn0o2bE4jVKJYPmSp8isGu5yrth0fcZmdnvE+SGl5vYIdyBst4yX42obVF++GB8
SdgCJpWbhd+xR59CXG7CddcFwnhA0n1jK8kIl2xi48RNla2zH2MKMSOJAO5zwNNlXCeS2u+DWTLs
3O4PvFFSSgfoddoaARioT1WL2I6uOHkb116Z0Vorg6BacT2N4j6IzZBcjXyBDNv1AqdM/ZRbxqI6
RPODekPAdLQcZRa/dgwphRaVjHWKBJac2xHcwV5IAC8SUlSul8WGG8XQ/pKsR5vXHsHrHomDGm+A
BBBJW0tbVh+dYeYpYshq8w5p2WNflg4SRZq/6FD+P/q8tTbDuyBHCA3BuVh/lEVeG2vG97kqNfdR
i6KlkXzV8hG6OjH6r3IuFiy9DKma5EHy1phaiFi3/4Uvg6dtfHEcsM2CzOBaNNL4GUBNISuy0w7E
43fwXN+PsgrBsiBC9JgHji/3OsOWJhp7WzxywteTjbn6M+SMuxPRvunLQOEKTfC75qq8Wwqfusid
41ZDHn1eOr9/EYqlfhuwzCFrVtQgQdMPxcP3ec1PByPtYwHbiBe+v3WGRlW9rvPsIeCPJbk3VloA
JDLYwJeO+bcGZIaU9DsfzqmdVU4uBoDUB8B26/O44Kc8cEr7YUMYL7NslP/7oKOtVb6Y9d8VxVt7
vlnV5K9DWChdErZcK1YEgN7EgLTHjyQTj9/2kor+yZsvByEdN5M764TTDcqZ7UKUoxIKUKiMq0tv
U1DfjcVBlgL34ToOdCIT8BRJmOfEukIFvXD8sxXE9RdAADEwh2HHGIIRcINPepg63mj20W3WCNMr
3k0ZEJCCPjWKwnCnL3biP7LRoFOrvxEImdGjYl99BjZZWOvp/3VDt4vh1DlK5eG9q35/RFVECJtp
3FAMd5wZb2U6HoDPwV/ZAPYe0r+Dz+P+EPS+6gQQzNdQjHHqiTXGHWNV2zEGg+0NBNyMp8udn0BX
wleKCjbZsiBXP6SSdGzxqgfp/gZXPxu/Wq/gcsmk6rYOjJkV9Zs/kJrT/XDLa/ZbyJ9MLe7zOshv
nWsMCxU7u7knWQaelAPQJWHHFx14rTyRjcbVzJA62+8lioM6ZFFsaHOwErPuqP+ZDspK6ljaCKCs
zSLxfHXO8Ar6oBp59IULf0WQerYKfj/yET/Kx7vk6I9UBWsM2ZKQ3yxwob17EJIEEUpMHtT6x4XH
uhmmtwvkwl4Bb7qgeXe9lQ9UIcDKyxTK4J46Zqm2rvICJ8P86rIbuIY/y8FPoQah14kbQF31oZ/S
UkgSqrb/bCLdTtJXIZx8GmYAmN12gPlB/GBF16/LVTexl8J/+/+Aeex1UNhjKVo68PidO+TAWk+b
gFw05hARzatZmdSBHpaqT/5xpNfjtmcv+TI7oFHyRJsbNVxC02RvahucSGm5pOsxUxGzvieHGu1J
m7N4uoVK6CKZmmPLMXPVSKdOp9v24ZtJG36Zsmhz0ozuVdpHU8aDjtasXjs7pNBpIqsfuxaGHPvA
EBvcHosQVvsI8wJDv9LYPjinJ4+18/BVl6WpTzbaIbxHDJeVAsY93AQoaUEVYYHD6Z+Gy7i1a0Hx
azb6k/61mewUAaDW29VLpbD3Qlo43NoadsUkpHSX2FX2BnOgIa5ixrKiZNrrhuj6zIJ+A05gmiof
mdXQZOrxMwdUkFxnFYYIuxgBYtj+M5CIBV8dEpf5ovz8o7R9UN466Uoflnro5bQrM5pgXtfzLaSK
nyBie9OwNFC4/37czXxE9nmu0GCmqNnL8SouaaBkZNDYpOxwZej5egqZaNXC1G7G1JW2o5IYh+hk
tK3SG8n/c3VMnxTjBckn/1wU9LCAZV9F5YwFu3SE5MEb9GgSpaMy5z0ll4fqYBwWETjEFkbPrGK7
dogkiKAg1lS7hF0VHgcEJ8qsesoOC6t67yd560qDguIBRPmR7Mhovm5GVD85/fEjhpD61laJIOe6
R5LzjHQxiYXxZqaOKuNcZqSH0N4Dywwxz3weYfIEV0DkMcV4b9WPMP+rp8zGA9bJYqv6JmY/7CZ6
cmsP5e8U/2/bnQ7gx+cpqKZVItsGAuZbif7N1+eD/gVhTb6khQYFbLIq2+OJvoZQzLEiA47OxzRt
cFRKe86URRx7/ZnJe2u92V2TfikOtqzOQHoC2YOhjY//639mqEuG0Y/xN540UvAOHSthZKM3/wjp
vEpHXO83kT/GuFPSOO/XR24xZJGFAZMXTg9RAhInokc1sVKqWc2c0jS1+a95QbnOXTzyA+LUOEEM
IEPC5dLlpGi57/rkb0uBPwIdX7ym8MhjmwgBoxgttj6GKHp7y08V3uDx7ruzjsH8ZMJzz2n1PDhd
teLNlyGCwuutqpapUNofo3o+ILk/tFkNhhwdXIEL3n5nJONEOvUEeZovIbN+tkPryB0366baGj2Z
OFxCIVg2Dz7e8hcRZHYvFalo+nTC5Kq1sbWPms3lfcc/08gdZSsGWWyEXqGOwnaaOYGYCp/BUtAh
IELCNB5TKZcNaf312bGOQFl3GUhi+VSOJ/PQ4kuNZScwH0FAp6wWiNGtnsgkkZdk1/5aHQu7t3nj
qG9b5AfBrQNXU0RiGIzgoWwIYUakN+9s3DeUY9oW3Y/olFIyDrxgxdV8FCWdPaEXVGZ5/aw2pPLm
zPECsa/EK+5oZamCIYo8V7KJOcX85/m44KyI3o5YR0JTymRkDGRh/CAXG4+M1f9OQlOt3bFp2f/E
eNxiASCNWRj6ECe/qWCneAYzxaCsSW+9ksqQ2bhER8zKxGRoqyZBIEjUFcTboagvQIkhtCfLyJ8f
w2tdZgUEi2hr9I3yu/JHJnCMAYAw05tDPZte5NmOYCc/cFf1tmS1yX94GBhT32gBQ5rSqaa6mwM3
EFUoY87LQDxwdTy84u3S21s5o/Sq2ZkPuiB0geVhtPrhmgYjMzVZJlot9Ji2eVIoXQN0YDrSwDRV
tKtr7jxmH7Jt3pSOiscopAFszaO2OmqR50z+mudNqFpZ4dShFrcVb2LvPv1xOvzqNycpvZCCms0e
EsbsdAl46S/zdFP3WNKDiBXAvtqR8PLZQ6OyxL67aPq6+Am0UbOoZ0eCIeDjUFL9wwmCgT57/KX+
ltWkv8GdTH2ZP7kSRDi9EBw7i/E/lE4FCJV6LEnmKotK6LKzWAiU4csZ6CjYZ8hwbetMtxlpnaIt
Gt6NEhCqd/TQyO5aTEAxIDr5WliNwjTA4bHbZMIBtfE32LZ5qGdMhrEnqVFUy0KeEQAZYqbcSl8R
UIYnc5aOwwBAh3F/suypAWKo3Yyl3RhBkjl+p22VsChLQmBoQGyBOnJQ+z1qkl2g6fo21RhIMMxT
p4Aam9x7YmXGjj3lyKUxEpzqu6buLkiRPv+WhpJycAl5IKxwRyIIcfZVazvhgODqt20F8q1aTleC
+vDOPmvZJuDjdj56fJoeAmARXFqvkKPLscbM1xfPdgftZiLSZjC/tICtBDVJpY0z/TgCgUcIZBX8
su9DYwVUjRWR3Cl/vu1BwBy2NzgjI2fIfbecNu5EH1lnZK7EG/bYGLKeWa8mTL+PDXqvCJ6ZMJzZ
ca6xZGrwmlwj2ZKvjnQjR4QiRmyfgtPpHJLRSSo2RFEH9u5vuRc86b4BEQxFXnYjb7E7JMOalOR/
pV+3Xn+HUC66Iko+NfLiX2E00xzM/hNyVnVgVUyKiGWhGZA0TbvPRV5fOxU34icG89r279LaKBcr
1CLEFVjsid7UxSIMi76QCqLRrkvwkxy6rYYgxSe6nYnScMAMp9dRZTIGS8qtoLhHlUrGc7pQisgB
80M2U4vutm6+vL1zUly0Dk3hGIyUdPAZhOYma22OzH6waTpDwlXDr00WABKJ88B+QoCwLIk/HKLD
Uqhv6f+wWrmb/uTGlknKcKEbATqrMPKZZkTi2RBYYhbOgpW6Ovd3V9SAKpbaLs0UAC0ppRpoWEaf
waNZZt4Q8V5SP1nJVWUQNw7IempBRExqSWFXWtOgv/FCrP0ZU+UwQojN8edsktvjCVKt6KO3H4cO
KlKtCOhhMaORIPheGTKzXMuOlgFaHPYmytWPTbkvYQsJc5bFp3szxzRm1/X2RkHPzA3NnABZCV6V
vnv40plVwggpfrhPI0jhAtEmf71TgbI/KjAMcqCafAId/igCi9GSfFWOI4bs2U5pW75NgWfYIxTd
d0b7JYmaNsLKJGX3jX2/5DuJd2xAn0x5ILBGve9DmZlV9hRJH91i0ElwAMcGq6LIXqkpG/oERGav
DTxKUFCTnmnnQHxNsEBi+HqKPXf664YlsFtwf33LmXzJFGm2QNqJIxELuCGkdwpNa7Gfsu6vrmpT
GXJWzBiWG3FCMzV0f7kMOF1ByGznKGhDHKZTXWVuyzVfkLxfNN+OdPixhJHjNZnFt/TrM1UCoeAI
AaU9iwHDIx68T7+x3g/obxua58AQAvF4moUEVFvc+VDObcpnOZRKBaIZ0zB7vJZxaNlB1JQ7ovLC
KO+51qL4iXvxCgTmOgVNMc05cDemypGVAK+z5YOwAxyajB7EB9mQjChd1u6jKv5f7ziYHgguZo2y
489KNPTEQyEh2WE+/1NqVi6IXBE8rRQkkZe3eGluyg8rvLvK0SrXrcZVpSlCXSt4/lOX1JKNKDyy
D+L5EJY+n/hyQSWS36r9Ixrc/KjJUBCHp4zdm1RQAiiMDQwlAz/USUi6HtgDw7cd3NPfijTpULNo
OQmynoalXMjAlSlMFUKT2iMK/LpXKl2LmLrZxjbX7TUOXNZapqD4EBsBxAvWm8mwmjJ9Swi/iOM3
PSXM5yW5K4m/dQqXT2x/V6ks+wgRbVq+u67A4DVYMCEe+c8rR/+4W2UL7Rb5491g6u6LoFKOyiOH
2ARKc74cfcrZnh+IACpoRkUDOzBrfa28bzSJWbIhWY+TlW9brUiOLcQ4ptI+SmipbxF9PVbutcML
JZMx4ZP3MBHRwRahpJiyEUdIhAGjitL5Kmb5y8VApnD7qkEheG6I3Exwa2Ln5+nw2ALcmvZD5D2T
mKKJgskLULzBZeYuO356tL6feBs0G1iCGe24cBpkm0Xrd0twn32fiHE/clDK8L94yDiddrenQiQc
zixJei3F8FfUcDq8d33JjP+iM+qJZVKmkMyyvEkaudBc5HP6GoHWp6j7lgMYUaFkwqwUeVI+i6CG
e8vrkMU27iaBN3MqQsQNqKMO5sY0o3ytWVTPjSrZ2d4wwN26vhugspcOGm7DWtSaeR1NPa21MMEb
AQGhlRz6pcBgiN9h0mD4GpXj/8uK0ksZS8O9qvku25K/07YAP1ag4Q3jn1QbQXDn3pmnhcxv0xAU
Ol+eZZUdthKgMKC8Yikcpysq2aGtz+wpCyOAknzsSh6rJ5jig0SsOzFmECO7Hnh8lec/gPva8uLH
Cr4K+VSI5MQ81N18dSe2zw/0iHvGLbf8NNfWZ+D3TCHZgDI5Ddvy04VSM7JS6dG4aEa8Q0BjKOZf
yuz54uIUWz2b2WPAwtyLqM4DMn8tQO2t7VMyTgdSALJfc32et2xkuyIQfqNatWRfUeaCBMK0psiS
xuMlZw/4ph1DZ3DEGfW4xlWW61QbSKaKq/DsiF7yEi5aaPSZ9yDMJZUgzsGKs5pEYEow5H7RdwP+
IlRwyKoCDkYRZ7mgiFgW4QeEEoWkXL6bkIzhQvuN950GAwI7myK98MnDWDwTtTFkAQmPXwaGPok+
0rrCRVm/dHWWKs7R6fgkt6ZZ6z09wadxN80+mUoQiI8pk66HhVO38RaxbhuW2we4VYeWxGTHZghk
CzndFdtvKNdWwn9ZNnM/+8bTi8y29XkhDcCzGnpZz+NnG/1MrJy14vctnKxQoI3tWLgwTKK6sPIT
sboZcwT4qEschdbPi1Oepz0EeVveKh4gH+gYJCj6Q/DvSUftbVMp2/Yq8uA3x2do7eiq+j7NQ5Cc
U0oN0a+87VwptKre4BlRYYyf/KNLpNNLKoMRGeo+pLdaxGmUEnHaQFGmSULz8gC+F1nM15GOnJJI
icg40VtIA02D2j4ZQvLJ/fct/czHE7b6Pdv9TX5ubvTByS9ZDnqGEgLwFLftQEAPjdTXdIGArVQu
V3F8y+4POcHEyo5L4AQbBg01mnot3iXlKUToI4bFEe3+sJK7eewncAASCQIsVgqbq/hOaS84rLxR
++0aOxolIJD6LnAdhBUHf3820Uy3HACDD9isae9iX8xOLssIAUll2TFarGVwPu0vx3N7o63a5n75
I5mWRnLAS6n41XJ2Xm2cA2u+D+kMbJskjpO+9wVBe3bUw3EWaNq760fq2FchIDXE8Ju+WpPbn0PY
Y5qKRy1lEqFzBNhcTC8D9uWbNs4U+KcdaIysWd5kXMNwXZbYjrPG9MPHDcyRa490k0NTK7qG2wh2
t+I6I2fZ1WIdHkNMBK1HW22T2DTDsX48MbIqG3S40npKj1XQLqFDws1BQ8lM6FTQ2LGDBaAUqdi0
Ne2XfwPLWcw4Jr7qsyIGQB5GOVqSPF7hEaHThlDuew6JHCgZm5LN8Fj5xt2PUcGoBaum8QFWoLK2
6qxRJPDZyc3bxRsVXpo+Yrebn6Nu0QX74hfuSobZbL+PZkcO6Pw1G/drZlf+8GDzoVbqQdq0oZvX
TJ3V+86IGj9eBwuKkII+V3UwWB2JXQhXcc6j5nLbdjYsSK3LTypVp7oQkT2zknKMGrQ6mQDQiBLJ
LDhGkjxR9wlIDoYE7ZmgLj9UwgSIw5Yd0U3BAT3NZXqg0yBWvgjlUk2IPyNSzkZMvdPDmYUVbR2m
GxzsrWlxpH9VyciEBpprxUzn4/nBNnGhXcljTzDsYWuN8REhSUrQRn3JiH7zQAgc79eoXd917/hr
ImD0nFiaYjeu8Wu3EMXvHsaRKsUHFEQV6WiO/VMoXoXE9/UE3gsE8osOTVuTWDfDLHi4Yp6QJ8iP
VJfOX9+jX/6Rd5g2h7jeqlul+Im+rwiYqa6zPxXyAO3212P+vZjbdA/krQUtQHfpr4WcxMkhoL8O
M7XYg2wViuBGbLBoCLrmNG0GBSWhGvcOYoGssB66ngDhKI+wwR02NvDfrViyx/MVpP3XQQ4oAuIs
7PGbdai69vw2DiTzQy8JiNNAf8mJcsDbr4AVm7bsXnbVN0BERMtndTEDLjreuPSJhmseWBmNu5BW
ZuepxhUYZ3hLOUF2JBam5gA8gxXK8/HDG3wkQ9hdFJ6lIXycDjgx0TzPNsl6Zh8VplwQVHH3drFf
IDoAdNFCIDJ4LOBTf2GJmbPEvaYmYtvOlxCDQaS56+TbMBvxcLeZni75HVIs0HtbAwQZwtYa0r09
/HQn1djAeVpPBST/Yhd3jyGCRXC5o4IVumR9t6IW7zZnYaBc7M2YDWgFeOXSXkQkfg9/N5xC8WPj
aPfzyzOn5LBb+p/0M4lLUMe51btOkPXGnPewa3gKuav2+tgTff6MKhvknuGb8uBXImJff71cu+9Y
IiHJecjnkFA4k9/CYAfGxD5Q8oLJMNrkOnAkDHJ1hMVQXIhQX5VGbrWdHhryOAmV97/rkgoWBjIk
y6YL460GjopIfi9AkoYTvbahkx313O8JRTJZ2OlM+XMX03jGQeHjtWinF0rMU+M6nLYTUJqjXVkO
sCKjbHN0tDyKVAU2oCiEKg4T9rbZQlQdf+/FkAAXjNbyLiqawp8IHHJTGEue+SSDIRh8JiBh2RGK
8EZ15HPmHl9BYqZvyOf4A0KdD92gMpqlEBonH90/pYWQQZFo1yclSlMXck/O9iPmpU/NzVzqT4oE
jBEiT/httYUZdnYA9XI18hKmLy+qySBiZcJYIfeBbQ2zvIY3f3Ij4pfZkCbQjuojBqpiVr9InCzj
t9Jx44KtybjMpCNpWcjfhjGBEyRN3vMqT4ZpoyQPIW/7l4x6Q1QMsYe+cGMb46oZferk04Att8t1
LO9QWxoOFj3PLhampkN9ruzAqrYgYFu9fo6H4FpLm5BmnqgBgqBR3U/u+vmmyA7tKXDUiceIHdAo
WAIcKO7DPOFWmlfvjTLRBMAEkmXgL5k8UqRAeRxcu8FdAnk234/PJYE2y0uZi1lvDf8+01bAMOr0
3wHW6leTxZg1+m4bKY42whxoj0eCcTqxCZ0b9Bt++Oayo4l3KqkzCh+tedC9Hvn1+phwV4y/0aVF
MhFCbj1vwt0guVXMI9ZqDUQGLhnX2NjG91o65sBs1z35rAc0OH9HtskWgZQbt3YLNmZy1AgPe7or
MmMdAg6AarEvtmQi89N/vMBwoSxtMEingp0tp3SaUWAg6PY3j3ddSFqjrI90+2R8pT4ov3+axRew
AIwt0pE7jqBNojaGs9kfj2tTcE7cFZq3eYZGkAmNbUirGLupptsRl66nwweof8PVDnhZtA/f8Jrx
kkIhVEpSfi8FdrC1UBO2cCKiHtG823vDihOuqmCicIdg/3rshEriNDnn+FwkiQTs1s1/pmwGrkOu
tmdTqILVSlvUddf7A5dF31xb60bUS8NrMbwCwjCLhlsUVgL7hIPWy0tkbRDo5pjNXBWypFirSuhH
JCEntTACiToDqhCC3hUg6m9ipm3ncu8YfciTMjLCb14KuZLWfTCMh6pL35x59+b0o2ZXSSaTCWim
n/Nmo2ETz8dxBnrtXlzshMITIBOcIgQA0CUzc3QJTzx4RFn+t5YQULesHtSE+gsSf6p5741ii+K4
QfZifcvdf3VONhOQsvlwHvmzOARHsVMqYd5c1f1qL/uGEFn4YYHDQmmfY9+gUwyRxrKGjgb7Ex38
LlCk8pRjh5a7+AtF6QjUzhzJByZhjtrS5FafN+akzrjfCdz9L1iz4H+f00gvnjs0YVpBRK0ZCT3o
191mcVP2H+eJplN+uJ1NAQDQYwcg2fFdt7du76aVY5wvpOGJXdc/in9fYULG+Rvl2D0/0cFywr79
urLGWrqVeRcPbXdFf0MNS/wYTVTGIx1maMi1oPZjPRNCEvC6GWxiDeqlqOSFAx5uzJVG2p/h5IUQ
WHGceRVFotlHDAADXLbH09prgnlLnE3aoB0AjXmPp6WLuim/lATd+8NCMD28PJl2/tE56xC4f0XI
cM9kRsNzzgUPImp+rKXdpIM3QkfvC/M5RInIGyrPqVQi0kW6KOW0GYdJ+EWrc7bx3WIbnN0QDXyz
Od1trglWvOtKmX93Xec6rNAqATYGw8N06adA30iFpVnqYlIAjrbTsxLNrTSR47z5ITm3RNGyXuRA
gMgHu0IDgJj08qEUGv1ZdpJ9xbbclq3n6HRJ88lATeYkgxYjEKA+B3YxxUnzNeyjTDFCp6nZR3mU
K7aQ0bqRkmropapyTIOhmtmdXdEs3S3qht90WOxIy8xGqUkMqpGcgvGpnlPi9Y/UDsPGqgdG2NMF
BHwRTLECqJkEzY8EBgiqlmZM3U7ApeUxb8w1zY1+lIpWoMiHn5gMMf2U0ygVdhw398xog+WCCvef
Fnizv4t3l5NRZJhmlaSehP/QZJk9L6LHJvsE5+QXJTVh9dX1kpt3kb4UCHBk4JUiL765ujrdO+2d
MlUw5i+DeutBgU2FZkHEMts+giLwNZy80mwwMge/3fVQFW6xHB/kWUI67k8P0v0XU/ClS2TUF/oG
b9VpZUxI9De79HslrvVTNgqz31e/LQOUE4dePV8PKKjRKKe4gtd5kr+h2vVWku5kQu6x/xMPtej2
5J5pNMTYPLCI2j+E0bH/TsT71fcyCLoT3aB8WGA18i1Y/Jq8+Tg91aBUZ+nqgP60VTIusMs5pRhi
86/g4mE4TjApMK7xk0LqZAswtLxSGxa14Lyizz7yElaLYWncCF9tUcbxVBeVfWpcrcYOoet5Q9ya
x85XZS9CFqBChgLlonOH01AeNnv06OdB4BJzlPKHO4osemf0lUdYU/Z7EwZ7HxFj4uiRsyp6sN9A
+V4VyfJrEIpDEA284QWBsDYj9uVKdJGs3l6bXP9k5raN0BCFM3SnhhKoO6O0VgDry7HXb/zmZE7U
AaOXD8W1ANpsbtll8kK+rtb9PHOEFoNTlKmSP2SGk+mB2p4LvrsgCJSd35YOxWiiA0NrbuNB5F36
w1T0G3gnXCkohfMGkXV6Y6Y03yFlJmQTo4CORBTh/oqylljxoYy2d6Qqo/egjpZ0SJuKh6xtflQD
skLxGXTS9AEYBIhhpjJf7ov9z7yLwNBh1VDHt2bTJL+Uf5snjErXqT+92a1fERXCG7+syZind3vg
+GbroL+X01WTNgb0Hbd3HzpVPBG0Hha+ykB4ggVizte93hk0KJWPiMn+u4jC1/HhSFKbC84B7pZ+
gAartbCZum55+mh3/9x/vGy4jgktEQDFYh1FB3CSc3u2CM3YAGiH3uaTYFka/q9LDr9yDTtMgGt0
hAHuY8FGxcTg3wJ5vpiCV2CC/tmwKKEv/O93+lurcflJYki3jOD03PBrBBLc6j2gV18sXyohK7zP
oPZfYB1T50vMcJ3Pd10dxuQ9Mnzq2Oqh29JzKmUiQHRhrerU90JttdUWNm4Nw/eM6d38ehDS/RSz
lp7JRFKxbg6Xf0Gmap0Zv/v5k4hWvy7+qGdI8UN8GdW1IrOC2tAW/T8KOebWnJDmCWd0svhFI0D2
x57revhbVRdM64DOVv9RIiz8ut5CFOTtUtoi98du4JaCO33KQHqqLq+seOJmStxtKIw1iW09EI8t
yRFRxOg/V1Y0agDyoGrsD56iVP7CqZbExriBP0j1Pv5WmL9O7MA3ofJ0/Z6RD63M6ZtvTj8y+uY0
NphVvyufyrwFPfu0E3bnvsmbMAKKghonehxkFPJ3+coMsDpMVTtysE73rqQk3kEEv2OF/7yx4giy
L5juvT4pZ9cck4c3Xz5h3vdIsm68qYc1WWmizabJHjdQvGxSbXsq38hFWJ+vsp03VvGe27h4lbty
n+FZOQdp8RU7zo3ESihcw0LQffAmJhMDsQvbXBtvBBBNjlKrYYfF6I8loOHLSb1IErEAZp8b9OQa
vlHllT02As+P2ZMs9nKue5SRkBT1vxS+itRaKHx3HebNKqaLscRagBFLSgli/z0GkBvinrNgyC96
Q4lf2c8Trh6cc6BWSVNw4u+3dWO0DwOkUUlNkiZ6VvyISxU3z8ZFMnSKWjlAnWzXFjyiOjw9IzQe
wcQqZL0AcjYS4q9QhquaH5ykqPiFYWn31WCra/PLFPNdHwly3d3sE3cMrZF8Gamv+6/vzk2t7Ekj
BWt1S20W3xwR9d4iQsSsS+VWHjL6rCiISZrr4ZjdM6uX1oe0zUDIn0fgPbtaQDMCeNv7KntzoPG8
3NGzA/+nEg5LUyakiRHoSnTnxCT2inUyPTEF6OyfDeir+0ysBBybHNHAICnOsF9a3ajT0YDlZ+Z4
QsNtrEGVxipepgJ6cLoDjiMsYKj4UcRDQBY5PS7kEa5BNicTVaTzdcW3fnranl8dmh8cQl7GxphD
GXWKCr8S70OeTwcSiAM3peWQw6L6tuEEGdQ2+cbrjyBBUaHlfw7aATtVpdMz1/GLBPC6Ju8RR5cw
wTnIgI7l+T0BWrNgI12lh0fmGdAUN7ySGEtTV+MAlgiivd/NprrDdhfw3yEqV0NPpRhVdQp2m9LU
7IWdLJPhm4zg8IpqL8+7cZRpcCwNY9TGQmj34m5Le7HYzy75abZyib3D+VolG6Am8Um2kxapCoII
Q3dKESu6qDOHQBoBaTfn1bR74BKUiKhtBVUU6jBN/9dVdYfyFa6XL6czOkXvbTuUpzEn1EnVUmEt
9GW/2zni25XikrT4p4AE0Hiewj+LGC/ywsxXLDdemr86ElMyhzu6LkJoGNZsW/moqsDbTiinQ3J7
VXt/AbhUTzzeId1S6L+BsepJKRNwPOLM5/UWNYgJiVqfsAADRN/Wepx2mEi7jyOgxWERICPLdzyH
E7D8IGm/HycSTEWV6eJ5B81zd0bwGiFVrxnu8UO0iewz71rsg18WPd1QV6WAu+lk/knpOEw1g0wp
C/R5XM4+QLQPmH43Cz9nekFxaw3ay0VbicvoPmNiISTgi+PCzgEWXO9hmQ0Gx28h4gTYHED2otTi
TQi09m6NHxGB9/SyHuA5CQie84k2WjsIiIBW71pphks3gvaWfyCY0DZArG1E00Cbg/0aXzhvYc8n
SStR3xFPjHAEqMeEdnrKAX0kiAPETv7qKFHQsca85Gn/ovlVycPxbWEu4eVJiIDlfG9ATC8kZcqr
8ddhlX2YOBVom7zWKbtYjBunghwE3YySfzwQVFWPMd27PUwJvZmZZiorf0YMdjU29E0eYRqLiHe1
4dXVd5XrbeX35/Czaw5IFqoCRofuKobl0b/U9p6dvLE3adtxtmpnZfUEVbwWWYing1zVapfnoqK4
ksgEy3DTX9rfm3xQxBhSwkWOwOP2TVckThqbsQ2QwQE4McDCAqnhlU2cmC9G5csUf1+rlhTQmx41
fmTznrUvPnL7YzqA7LgSAA+EskeJKzUMOuGlBdaARynE55Jj9lz/teedSPGId0V9bRgN9ysuxykF
J8G3ff13eNWEGHwwcP1caOsnX5vnkNUEufTDYFlko+WlL54ieeZCQvjrO1OjLVu5Cf2iHvq8BsRZ
oUtLrrKCpRYCbmpmhHpqS2w65HRiGqTdTz5Ft41Kjev9wd2MGDERwmYupscG8uyzDdjunv63Wth1
dJiMyuDS0Gb88V4BXRXNSufom13uiSuUdiUyViMqZTHqHQThSLu1U1hVDJTqNNmEuW/UkqYyMJWW
p4y7ngMX93sydmeDmu1kDyrmroGc8VsPlJP62bl3mmU/VRsn3jo2BiQGrsEyTPeUCkiPP7zXplLd
YUArssjiwZ5qhwRV+hhRl8tkOZzWUvt3oktIMfvGi++9HtngzHqGmLqkoL9Z5f/pjdZauJpEaHEZ
lJ1hwA4RHaSY4iuYx2BdHSXN1G4H/A3nm8XwqKyrib/Is9n+aZM/aeXubVf5uHu242Co6V0FOae1
ZwCX+fNbtncWHjKfCXooLRJIqx1ST7NY+Soi5Ch1qX4yEg4QcZWdNIGFnRZ7juj7S19UqdlRG3Rv
W5XW0qxtGeDhG1DgCKd6vSN+StqxMJ69ZoYQjj6sd2lvAocG4FR29qtCk+TqAsLmdYs2eOCuVgnj
6N8afSWNtSngjN9vDYkuBrseiFKDASW0WSAxfKFdjXEe+7AiwV8gpVeM5+mTWMmWKcdg6R8ZnGmj
B7niytwEi6B09yqgsc+vrPNJsYA1ccTCfa7ysFDA0hCxAGEOru7F3zbG9/aLG/L7Hya8gleXnZy6
HomyWkAKtgLZUPB3X4zfGc+qNaCwNifDzFaPCVSz165EJLIaacZ8a24RECDP8KZoG86p1dg5yMng
A7emTxureiOpjbTh+4GjYv+dVQmEWmGFqKFJ9/zJog74PoKjiG44FQpSBMITNZHYtKzp6CA6uPaH
LB9JufxSLXhwWgjG8lIldyflJoj2EubIrqILS4W4qfuRYn/sKSCkHUdr+GncsY3BStm5DQemiPoy
I2pGqVaTzZPaPEV+rBsyA50QcTurhze+0iJ96YkcrjKSMUpYv4VRczCU84CtZrNnBcY/LQ3OmBJ8
0RlYlSOKHvR50YXJbBtoHwnIhgl+X2M3Ebyxi112B2AxzWWb0SRHWsUlG6vsaGtyC1ng1ryF51ua
tm4eitnmNAcwPuzHU+h5S3E2kNk5B0QplN1AA92DKgh4UEn6ozJv9KL6k2TnSWmszaQAPj/7aAME
sIh506amJkOV09nIEsFwJSgGcrLaVOhbYGePBNLO2aQv5V4gKkC1D9xoObmtjaIzucGQrzJf0efx
sw27582mcIxi6UmnYfIBc3d/kef48A3CDQB/3R+gJ+MxTfO3+0alVtGDFMALKxF5U5H3jSoJTlLE
9FiO5Iavhmq17x+yAQJhlZUFLYeIsrUkHba/lL7ORcxDXIBh8IOwhBFrLLjcjFjh+2ntVijyWNGZ
ijrr5309TDqqVz6bUnRCTxQOlT//pkoxhF1kDUSkjJLZdK+ejbgezukHpI/cmp0//JNgMXFToyAd
uoP2d3fhAmWNVW1e0zvGLgefWNX+SfG3RHgRIHH5i7uXkCWOoUyPToGPgsKzW1+B5Ga7UN0qlfEW
wUEk6GYx2Z3XnY09RUBRVs3hvvO+E/V9vBhqlrSzP/lXMmUmLX5scj/zminc/dAPvhM1pC/k3ks2
GhT0qld/J6M2dtVTLaZIHzSMItQOLqyeFHAeXQyNS9/TqtDZoop07M9kuqp479eAnBq4qV9V2M9x
9jjD9lXyRmCI3zLVlxYj1692KBAnTCvVI34epbnXhnjDXHcbaIxtLHGBw5slfLxzau1CEeApet7A
RM54/Akm4hPl17nmzB12wPO03RRVUDsucvt2kzjWX/yx4Nsk/TRb4xL/r8Gf0cOXB+hqhGkGI88L
0nz70f50g1DzpfguJC7pP+YrFDFcFI7RzqxtB+D09c2wiXVjlfkHFQkhPs+sa/omO8JU4C41Sfl8
i9ZdZqt4zwgjHljSdJr4pshtL1Q6vROlhNpmgBq80Bw1x1fJEMKpfs7pGdXmQwfT0ji9c80gjnus
yrOhfkEPV6NHrFyNBAXQ7SMVwgAEnVeqgDdpX8Eph+aCOw2c5vKoz3Q6nMAPgj9lOdzyx+cRE2Kd
USjeShDO7CJ/2tbM4wbApiJ9rMi+1bDVyjUR1CyPo+YZoyreBvRysFeKhpzazUu2WlLuZbseWoff
9mV/CyoEqAh1IU6nw9yYBaD8L0dSD4rHj+ysYz/5tl6gEZhIdvmLqn6YbGOFH3L5Ovn0C9LboezR
RflUS+GGMpQrYpMysp2gXma2lJquRC1TQZ2npwX9vYBwTCUSLwAAd5eNaxQj2vg3zYNz7npCTlqk
M5ci9gSFDeuIDNWhOr4inqnbcBXeFyJ7xHLvfwRWT3nu4tXx6wcSLpiEQcwYuVIrp2ekyOnp4a8x
ok5eJgZuNTxDi2/DqVIXjn2XLfgnuHUlrEqN2/6eEMEZjT/xBgMl9Vr0RgBRBco+IauFXP/wQsru
PV2/pzDgENZK/P66G1OQgkJ4US7zi+x1sEvrrOruiY/FAvTQ/726e8y7UmMC6/giVm2Z0V0OSNYf
/FBxFss4ck8SL6Wg6nQ8o6jhJABRnhB4XCRG795VFhBRtsNMNT0eeLoizXZ+KjSwK3u4svPG7N7t
bH/0bJxQSMw0gcWf3ujNybqxpttna3qE3OKykJxVdr5733paimfr4rweymAKbH4TVjll7O24pMcD
7gcyct3vItepMRboBIzvC8QSRo3pxykBRFwnnIHDAwOaOhXtlgkRy3+53MA1q1OuEq9HBI4SD/uS
Ir8y8zipcs622xi1/hwbS1U9l9AOHWPzfVkiqOSkzGa9YzL9mc1hxICfFzVxfZrAHkipqwOs8DuD
41i1Vff44/4CppIooaqGaeVE571JtVYXKnkAIVbok4mP8/REOt7GeP0C6rN10yhDlJpzJLRUm1l7
zV/UfExqE/lAKbJhv4Rv4s7O/cxtDQUqNnUXlQsu/ehdIonWa25tIYF+dKxO4bqx+8m2pbKsyxQ8
8XpS9N7sD11hJTcgjHGFh/5VYq8avIChWLTIwjFdRcO7ne3yseXsb1eH64XJXasStB1IBD3tt4YM
+rusQleM2K+cCz514LvcGtkeCdurPZMhIZTbaYDBvi3W4gqb/D7g8Uvb64wJcgSWRgAL3qvUsanV
u5fzzoTO46T6QERZnPxEKV6uBUlFjaAWlJMM+YODM15jqZg5/tROaGWceHwe8QzNsac+CGYTk4rb
q68QQb+bKwj0uuEWiErgQp5IXjKC9STKfOMqL1P/ED4eq5OzAC8V/S9Ug60k8NVivH/1cHbezT77
2hJlYXMEbq/wtXKKHjJIE43K+pPNJCeJi8ASh1PDbLKd9pPTSqFcmH2q98IAYeCUCRbjJb19NfH4
Aa1Gj0s8oojx1j0Ehg6VVWcwDFbC81lS2zDhJDauYiJ71vDnYSjYupLJBwEXbbih5ViLjicTMAW2
RnVTWqHVS2Emtn7V89A2J0d+fN1k2blYrIwbVpo3ZXv7seEmU62SevA/wmWnhdRN1bE0OpR6WNyV
aVKYHYyFJxyr3XMFAi+7U4ci4InbleWSXkNugOeDdjkknl6KmBxAc/Ihefscix26Fxe3OupfRWUJ
iPHNAtnAfsdRQ4p5ITzT5oCySby/SuwA3cKFivKS449tSAfTUrebn8SYwAe8ddhaDQBfKV+TdUsz
/BP6Y24rspVEm3b2AqRQjtMI3g9jkeuU2smd4XT3JU6//Fd6utH1A4pgvdZGlE08V+/51hYjzReJ
Qcdj9wwh0xaJ0HWvdblhEn6/RWQNN/FdXqmIwgwzUjSUwRF++SVnIIjsnNAVt4c1POtYF9XnmFCh
MjShZAIRvGGQJwwemAsGy2Fp/QLsXXYHDiw/Sj88WTDEBsQh8vVPou9Tiimp+in56RvbRLdpB3qM
Bh+Ozyika1ahRLbCyhkv66ISFb4nCjx9OID5PolOC4BQZ5jH1HLGON1QjpiBfWEWUsJfEetbH1Jb
eWwW+Ha2sKBJJt/WQ/CHOo5pgt0w8Yg0u2ML+oJVAJPwXDK6J4OaGkrh0jRVgOnbWxoYdMCg2CWg
DQKe5wlYOVo40jIInp+QaNhngLE/v92OwJSbUeQwPhjBZojTjGw9pbuvgruKnlW9uIvcfs+LBrGA
GeVBf0ijygqEb7ZYujcS8p3gkkIFX56egTlt0NEeOrL+fJgIxkJLQqm9vnJSyV+2NDcJnUWWLr1u
LQk0hVWhaBuKM4FKzI+usqBiPT3ff2FBjtnX8e9bxBp3dN0eGvhCx9rMAFtovyY7ltiKH+zc0Hqm
u+fFitRqPZwDWgkXVDw/J8s1bGv4VUZ8c4+uQt5ejDCDIG8EJIxAE5KzXw9B4KoLkEEYL2W4PRb8
/I5aP6ZnRAjC9Jezr4xSRWWcqi1mSxyQJ8JBOeefKY3L1tvckEMAoOm26NB0D1ftLGu6a9rc9QxG
05jiPtY+zPNB8XCjzjEZuuROzU3QwHE4uTlIE6x5AQOoGRcifbE6tvAwWrYeKRRvYWRw29AhnUmY
roHTJOxXXDB9AhF+7gpX6o94Lgl5A7vrDO6CBEWhPqD0ZBgRYyhl/sAnGbkcOQm2ABQTMpwMvbrC
nh+X313gB5s2j1yNswyi86yqB0eG8//AdBD1/xE3h0AtOR6W4VnUbVGq9KJZkFkMNWbY5hk22OHH
KTS+6sGnzGlNWfKPyphb43Arg2D47TXrdeBfg9u1JTrJWi9tIS/lA7qE01FgdmMpd2D+9bHOwqaR
r37gtgZvTV0f/yb0aPS6v//eDxywuGm51nN7UO3e3G4FgSH3req2Oo4QCV0qwiwez9yY0GIm8iKQ
Q1M4AhxOiqL5vLOB5qeMegZTVO+mwlZA4o6hitB4KJ5nCRSiucelXkFhNtBHKZy8SuO9RsPocN+N
71WwGA3w3Nd8CF6ex5DPK7vJLWLlG/LvJ1CLDhXVQnCZfi+QkjvsURrdnzc9n6teRJR259naTw5Q
v252QvTQDhpkhUZ3Vcdypglvt1wQxIgn04ZBatxgDMr0t3DfRUAafVOQWB6Rq8ANlO4FerNPC617
ulJQy73ua86CIWB2ewV4YDGU/KfgS/l6D8bZJpuxSNO3lPlBt+sptHeycFZAz9vvqWpXt/KGgQBD
MZnrHSfTHgugxE3AnHhzBOkvvQ+KRNOkE2zDIFzNkOJuNZZt9jWXyBY42Q73DbUIYqurHp5LFnCN
TdHGI9oaMm81X+rCJbGrhF6lTHjMmz8D0wrpjSihkqJ810s3nx6tLm8a4Ctmkj0jdg3HYvCnNE6w
M7MGHXqYO1eovIIzwcAaaFotsJlp5gQH2qOnoDJ222wvRFPRPXkjjeOcb2lIxGj3Kck5h6uBKlcX
hIEj7GNyNUKht15Oxs4mW7OuH8YSR0FiV1/OHMFi+V2aheZzQX6G5sHuZ5+5d4Y1+myR8DxUGy5t
LKJXnYXPQn87jsBJjiUPBTsdiYcrTMBB7leucy5L6YQZJxAflrSaGNsPnAfiflJPWVP3V2J8c24K
+6ekciFWUybXJo5uLVbh64t7OFMTrg8UEm7OOcQ16eQxPQ1Nj/gcaF8Q9T9zVqHbnX0KNLoQV6K/
zG/a/QWE8zOLkCZWEK6hlRrHOg9C8sROrbQusiDjP+KC+zUIbdu0n8RXohm5p3+W616YgGVUBsw2
Z/WHKpceJsc6/RkOPWME4XAXLweB0hIzaCPVLdbNTYA+Y57QhPyo45RypnWjdYc6/5bnFeMJxGhd
aJHIb2Z6ktUod9qrot+swZf3SNsJGX+/MNAo+yqAZGfxHOyHOj2PX3yzeDbARCLiZ/y0zGoeEsjl
70lNVswk6g36A4+d/fueoET/5Y0D1jkXQtBlNe+iq/t0xVc4TlrmKgFq0hMtFHQe5L/dw2KV/3ou
Hf82YTAO8Ws5LOT6qNlQYAFrONEzIVit0cgv7eiJY9ZKC+yYgmIMIXjKlEwMGPxgedr60eNQ4pb/
xJjUq+Wn0CyLfgapf430tpDN1Hg9YZS5T2ZpYNX3lMSFVW5/Yd/TIUdVDcnuF0gXeoFZfkI/v1j2
wEkpRwL+E3bFa7i+JsbrX8x/o6ScJaT5mJpT0ZPJzCkSdlvrj+67sylVwiwEKfLDzVbunzs890c2
ihbz+TYYAiNoG25Re6uSvY7YaozlSFS95UxhRFJm0vXF3uCIR2norkaYVDmg7UnLu/NWkNL5GrNt
VA9CFnGq7CQDIxeZdpf5cyt3Q0tzTXzcP+hM1ja1dQ4Nij08lEHJj5mFVQqVpK6/SJOPvYJJFg4b
5rS3T4QZKtJRdaJFJe8jFIav0fEpJ6QJERZ5ahUnCOj5/RI6hD9e8pC85DDJa7KyZDpvt1R49Gj9
Izglo68cn1Fiv0TT20yRmE2s904meXxBAjrAeocATlwmKBaFD18eFWUvB9odXfOcQyyBuHmRO2o9
g4YW5qAL19T2nRs1B8nthFCO0snL3mEwvuHkufL3kVf5QCn5HxaLShyANIjLUz+cdHEbWh6RcLIz
Onc8WrcjJUvr5BPSUegWpPgO991U1kGCA0mt+WnbnD1KSU2SBg8iAjSyEvy3qV9SNKbGOs7VmHdb
aYO+7BNO44XvQP8/y7JO3K4Kztr0Xdw1PNf82+c+XTp21FZpylu7/pIBzbMGzoUigOt5pln6R77j
mSa5G+RQpJZo+AmV/4DD/z7xJwsyfgtQBSsni9FtqYRkQErX8jW9FRaS2FsbThQ3h+QJN/0EN0JS
/ggEFFqbs8x84g2ShZ1wAVsG5HYCP4loxkDYbIxO2njIaNArAqPB3fl26jR77xy1wOCk5lZAdeYL
ll+im3dREzifkpgsFSsh5X4/USmzywpfQXIZxLSQZcfXqI9WuIC+FRlN6uiLQE+qyFEHSmqc2tNX
rBRtB5Y0j0D8BPXyEuItG4Qi/YMhubAGqU6E9lXqGQcNCcaZovL0Wu5ZXjTqjIa136hn0DrwX7qy
LbVdsy2pwLRO4m3wLt0J1piATNQ7gHCk7tT0R+DiMUybBVfPrQ3GpocXPSIK4fUw6jmmZOdoZbgi
O18ZcCNLgDjszsHieGRoahPc+a3pf7jCrnBeLfYm/0ePAzq11zw5IBAA5+lXtLxpVbVV79Pubu3X
8v4quAziCi0N6fpjFcH8clGVLRVkw8pDgj7MyICn1GLxeYi+mS7fikn3m+TKUu+EQ2SBNNVt35/i
TGnIaOvF1ZvPsbcTg0W7VY0y+l1QR8+jvuLro5u+Conxwdq5iOVgXBxOaTTf/yfOwLFo8IsjxFGV
NjTo3XaghFzs9MAKMdnHZ3PNysH2FqxlSNeUMEJ9XipuiENzG5i8CElBR0MabZJMjEmbOi6gTlsB
ApNQJfVjILnYaMUM8G+qaQbEP/Xck0kyBS07CAi04pagS45+br06WItFe3mn1O27DzkPbkQFSLAv
oW96ppB8niW3PGaxvn04kGH/aONQYTMXfBsB2uvAw0hV+mmBQHPodbRlRFbw2aBxF5M7zgmwWmdQ
u7JbFR54cszNftwGMLbDytcne5TF8fKJinJncatEwRWztrJtaerQED1OnnL+n7Bo6mJga/cGcw05
fNXy1X1VOeB7B/SNzR18DXcLMI2PcNR2Th7j8SsIEAENVu9E+hEScZ8Xq3AbLXWSHWmg9CTXsZ6M
xaqrjH11ig/yV5E201BZIZsrkAmy1+UrilbmD+8RMgLVAGe0uvNJRX7Cpo0hes9CAJj2i4II/Rf4
iYEQ0XzIl+vlTHEt6VO92y+PcEy3FurP7NfalJgD3uzzTf6LfQQxhuKsJYYtyI/RrLdfM3qCId7E
nRZm8cj+YxG1M4vkX1rRdaxe4GIPu/y/yBHRsi7zGOsx2rclhyUxm7VUs3RBZnAyFYp+jjdB4MCh
yahXvbkfxCJTZFrJoQGJZqC0hXeslzqJNgaI8tAukJU2TVSQGlYa3k2NimVDUVJX5tvq4QS6fTxO
40lQces3IkP+c9PR+prymjRi8nLypgn2nPviE23k59U+t/gxU/QhG4UVIOq7smkSidwgkMMfrZ+h
PIBWtemWTtcNLGMoGRxylZsLAL3rsNaPdjhDxGWTF2vy/ucpssq7jcyRhbVueFSRVrI3+lSpk+hT
SGIWOBYYlFwQwZb4VLCZtKkExFylfnQ62S/T655V/LXNfQBOg+y+n0Tav2NTnkC6Y7Ybvr+cZe9j
cLCQgbZYEhSfRIkfcHf/5GJqz/zBiSgjMea7fgiyw5ArRecysUpzjjHBccOjtKHHAAHi+/U/GQb1
eXmGgC2BfTuUkGMbkeiX2Ad90HXht5dO6IX5MjMDHEGUET2+l80nzrlK7TAwz5SRVqsg38Tn2rv2
Ip5vaen1tPlva6L6dEtQufE9RhdI2J9JfsCBe8h8I3tE214hmUgRTzhSWGdHwYnVmnLZqHJqzd5w
mZnrHZNcIWEQin37WaXJS8Itd/FOMz7OSGKhq0Vt7EPPV130oQffvWteX5PtxLCG30ajtmmAQzIl
O5H8IxvNvOky6ExTYHtRkLxrJuhOa8cdAxbQp6VaP3T5iwf2UycjWvkweJcbrslgvqiTtgh8pWH2
zb+lDt4DE8DqmpgwSGpj2p/AIUCC4+tZWXQGPiefnpE6dKW4nXDuKDPxOxf764OHaOzNfHpOpbMC
M+CZzrC2ja4agZDSZZHEsu5wUu4U1CJVQ6c8YpuKdQdF6g32MaBJmCKXnhSWSiFaCmhxdBlA9MSf
AT2vbVCRrXYU11YCjVIDDw3hNxviMDLIfSU04LgYQLZmDxuBypgxVedctqiHYFt/564JiRqDPEfq
KXOxHC2oY1AqO+DbhZqdPIN+bHW1ffKyvQ2+G5tYYsYVrTtvOo3DDm0EI/0DR2yzBQMhxexSwZI/
+vSGYpU/Nc63xHvisdN5oi/JjWDoz/+lujLJOU1nB4LVvC+5LxmB9w9TORxKHKt3GQb+u4fKBnTC
V//L+6f6tCQGVlYEgXCeQRDru/4+APpKfJEhOCt77yoCfRGlOQmXv+n9EYHGbbkoGlfAcWvw7QRk
qEiZLdP9wEc9sZPd0wmLxvPgJcwp5Lwj8SyWVrn3rXR6agSvp4tOM4SvD9EazXZhQb9TgBt0Fg0f
rFp3s73Xfr0ro+Vag3CE1e6GCEsAcVvQh0STdDYdnloW2LWLvi7o3vl5LdUJE523pQ5ZRNauIgQ9
CMkH/V1s4T5apc7BaKq9QNCvu+xeXLGZXnAZ+ZnapNRIiiBeICsxJ1HZj2woIkPeuLNUvHwqzNtr
SmgCWQ4QJ08aHBHzTCEo1bn8SetVuPn6gyUSnigT11zEAPCBVNmmxy4N+AUxt3dwGO6vCzrETGAt
cCCxPHHbCxxa7uBA8t0CsuFKc+iMqrx02VCTP/aUAJU1LgIGdjGskD0TfZQkxu4nj0+DXIqpyNCd
Uy4tlpNSXCUK2XzkfXeVLYARUTdK2VJzLGHFxCvnABYJi3Ockm8o2wdKcxSIUzk4l2QdMQozMLyZ
gxlgOp5+UjwpFBo8dRM16wzczn4/BD+bcEmHv6sWryZK64ZGOJD53AKIuGRmsHV5Ig9cemxF/Tsf
ihFOnDZUVf7KDUnIfqHFWfJm7pWyOCspnC9vEZJocitlLLBpC/MC/DYXLTRqSgq9xoFMR5kbX59l
tB68x5B6cnd5Fn1CNytDbKZVDI1iPzSZ5vzx9JuqaS3CLgP3CpZlMRocOYX76L75fx+CsRvAdxLn
LKIJlAzra94yyesG208bxbFDJseB1AEcFYFYozYr2WRtoJFQakZX5P90Z7SWJkIChtB/js6aoj+G
7oQwU6xE+e+BdAL9JjXZ5eQSEuATZHyAi0W56Mgr0NQU8tqVKc2NHsystK9eKMnMZ46BjDuw9RtN
0hGlcXJrdVuVCWGy3XAuwNGIuIG1MXABpXooiW6nqFZSm6TTxQ60utdBNlyxLqKtJuGtvWnNw7Fb
RqhDWNypi3lxfvvZ72BCesCsxp3MUXMg0J5TTIAaVc2DQc6l46lCLsrNzZfRzVUl86mjjW78QPD5
0tAk7n60RFNyUl1ataVvnogVOmNclHD909vwOoqi+zvS/aCISho4trDF42qklH/q+wHK9zT9KOXr
noyyRFBcLM4b5TXsXaGJiF3etNQ5vQhw5pITf1wNA5r5hMtmrYmlG4bEzwwNeP47fZAlb5yDoBX1
+Jaj/yRtOCpidwCX+NOEJ7cGcAl/f3DXEp9sbLhFWn7Lhq0paBA94+V703oWoN0lIP/shByeYt7x
UwRca3QH73yZwJA0+QBRCZBIsWWmgMIcmMAIoY/0eghtUw+amNEqlzEm5Z7Bw1GJ4ygPUSzPYG6m
KQTOA8TlH0HX52CBGBarSxE1XsChDMoWQqIXZARBTb7ASjZd9hnGcLDYpjadtOBYEXr80JXLDjcb
UNm0NCctbI7yWfACI+Duu43l9DwVaEoAx/Rq6sjWZRNu9ze3xnP+c0JSjL4aAuvK5U/HC063JT6K
aJ9gAnrinRgtkBSxuFIzaX1E8B0vLuzWFG8IgcUtvfCh+Vzb+DFhFCVgouEvB8+mhAJR41XpD8cH
2Ni8JZtbraEr5YO7b9f7vCLJ3CjIvHY0H0/tDK5HBufMRrBk4uDiiPrKfx8zO6twtsYTK5RzqwG+
UK5wAjlGIC+Q6hyQkBEfTlw0etidu+qqYVY1u2dORn7Gse1pNeITYDhyKDSawQ1nftP3lE+ZPRol
7h6vWc7vIIcWSfDb9ksCSn6YaPVcoZ6MDIMwwahGHWV6atYyEXOcWuD9np8HFEAskG8SYctIMZ/n
8FC0EgRC5zMwwwiQQ6mFVydC1W8sVywWwN31jBa7W3WxUAg00EajLjTCHtnMYNYdDDWspPP4ueDU
JvexIOhmf+/aCtQCYFFn3Qhkk+a7YpYo0/fefpri24slEqFUizEOD9VWQEfTWzaryerWsMpm/waN
Gmro65eqC8uq/V1Bu66BA4jQxbv+ON94AhpPV6qBShbO2soHxM89B0/HNaifieXXbBPshqHnoSIK
l8Z1E+JpBzzzy/x7Hkh2xWaTxfU4Sqv0S7nChXFgXC7N4c8a6bheYwv4rtPgky/ztQ1YW2XEIAbc
92fLZXBr0ioopQF/hq91Fj6lGxG/d+YMw2GJ3NOVqzpKKpy6ndQ/22X21gAdKeTa9BuRFVkVG2TR
Eje1bFu5eMhYX5KjRdhOD1tPHsxufJwzHpmP7LEk4xfWv9hLzC32L13uMgNWsBEDOltwPXU+15/o
uW6P+J3EHX7bmplss6aGbuOfbo6qHlPLEVAMjlwS9vslRXTVJ0zY02M4zHFsgBSavTjA+HfMd4Pf
HWY0WE1HraxHjS6RTUq/ox3bxYTV34DlRpObS+W76fTziFhuhEy9xgMhhS+uM/22hE5vz1DELApf
ueTlJWiAqxewLe2tPfbXNoDtf1LlcKUMm6eOYf3y8aPkadclIBXOmZeHz/p5RP3D/RIOF0CLvEp2
ycTr+WN3pBaAVeqlhqdqyniIQk4VpAuTkhA+DwGphUd1Py9wp0vfjhR7uofyX/V+/8vlkzQyITdZ
lnUGhF7N9aYEIs7r4vqdaoHrYvPkU0W7IT07KUJtG/vPwZ9higZBqfvXJjx0qNMhN4fvTon/IxXP
LXDrnvC4xtaPt8MjMHEg+55QJQIh7jQ8LnhtbgWa7vGvZ3kWUiVBbvO44WxKAZWuNllYNGjSljzV
CBpV4H4QL+VacDj/gw/CAmyJPAhcoCsq4RZFpeI302c89J24pCqRUH18d6N1AtrwpqfqHMWZHbhh
qyqn9EEjPKAISQZAkOeemIe9XD68hdwvisAGGRkFNNY5WSyTySRC7XrU7jkXIK9OxG3PJkQt4RmQ
j31qwk4Ni8JtR2ooIv3ai7OkcqBpX7Ljmx11xsGkOpc/B+C3pWyQRWIVD3lGX2x2lXj6Jed1bsL2
BqpG7Hd3X1oXB0yWluZlmerA8bbdXUqJFkbCtM7idkYf5O+rUcBHysRh1KrqYxXObuTFOmlskG23
+xKdUoOMV4MTy1RuiQSDV3D1UOMD/45stmwW4LPcegOn45WOR66ljcLAsmlz+BmTksoSI8xu9/dz
hOF5QF4M9+3My9bvXvzAfCasqQIjIWYWfEp1yzFeXM9Lf70+4HEoso/KVOP//Xen22darWY8r5iU
DNOujlaKSOrK0BGtrRnVZ+LTJwgt/2qNuS27JF103K7sNg8XhM78BUIKISa6aHxFgisWvFeRZ135
pII8rm3TI8FbK/yZEbxPw5t6orT46kcGdaeIAr2g4aDJTyMJx4N3ivYuenMDs95COKeP0rLyQ1KM
Ec/PXmkhbOmU3NFuiVqBAKOTXslJq1E355Zqow4hMWmwjMhZ5S15+7pPbmpXGtXqBMI5i++9O36d
eHNQE7rozSfAhvplck7YA7eXYFNP4n1EiUPVwCHnS1WrcigaiJkGh3fDx5JvEMgZUeuIfz6tYCwo
QMGrOIj0xzZRON6tLMuDZsqKOCpDiXtTZ2mApjT0aguZevAqDpYfg6LAOGu9bt1EUOvdJGxq0NRb
SQ/1UicV9ha+jFfCj3PVJRzm9L2uCqE18t/hqxUsZTBwAWOJGqFhm6/SmcoBLehuDUE+L6hYAZUk
6pxMegnvXqwTkrn2Ov1khcUDh1CcMd4Gm5cM1wu4bLJhACWaCROtBItB+4FclC4gFcEokf1lsTFK
PepMENDeNfBmNRAjl4ZhbPrSmJtog5dUVUACB7tIC+CXnW5husmYezBPO79DyaRSaeN2m2WfVIPt
nYGqfMvL6gn1/o9dvf/rBfu9DbJbtMTo49e8XsHXr00xKNE5KPVDCywP3icj0oPd0OJwjtCc7U0+
XRSSCUhEL0PFX2yp9XCx4XSCHYJwoMbVEZ/ylmJOrwz0++pg80Vig1508pIAHvKzOxpy59ENuWVX
mQVUjhQvQCi2cXAkEthDHAEcV6Xqa/uZJlOFb7zDakHiD1vzqh1Z0ijZ4lqkh1XA95scCp5K+zEk
0dX93e3lHQPEbqRZOsRud5L38g1Z9MQ6FgDmHj5S8oTb/9WYP7OJej5WP3FulnM887dti6VN2qBc
s2ra3lvIlZfbGbdte+JYgd8nk7vThi8E03ENYZIJqKMNuR84vfQlh00lCfbcp0tB08lgNjwkFAEC
FZHdqCbr9EJXy4Fc014wLJ+0ExPMZ3dMwZn5Ym1TMJ2zWCWsxfFXUhDWbKAAQlQZtFe2BXbhwNxX
Dk0faXV978tGNu2sbejy/17jWUSgnaER140qj/t70b+yBsWpJ3bcCZK8+yc/vJ5Z3gw8rWPOLz0G
QpadMPLJBg2f2oI3ALaVYZkmZXuuqSoGMlo2RxzrYE90C7aVbv52fyD9IfrmOsKHLeN8hLcmoeU/
jFnHub1YTTxq83J6FCpU6tDbcwVltfh5XPN5lzK/aoIZ/W2vjyfclZplRKrjCLy5d4tGMef1wcgj
OsvomQT7npHzVWeqCsdg+YrAnkddKPdnXg3nx02e5yLBLHwxDrTP3UO2eHQwukG+ygMkzbvomeSZ
DUuCvb4It6lWlGB5HbEhGdShT+Vs23i6uS0iIJ0qvipXk9DEJlTT9ER5quzrW1uplKYuyyjL/ONx
lBTlQ9DEixh1Ea1ma+zVQiAw2Lrh9gUB+O10PW20iu+w9eLHclGpcd98XNCbW1jLr4cfWb6z65MM
rCCTPq69dA/UDed+iN4xzRRn1KcemlYnRFeMJJdS53buBbmVd1+K3Y+GCC18GWvbxpD2uIWHLooz
AGSeIWH2uXFq/+aDdGE6Xs/KljslQ43DdaCRgcS/6ZpHbDYYl9zFYnM44wv8ezlE5TURzB1/xrgl
/G0FA4eKGGDdkNAJdMXDI7lh5nDGHO3cVnNgjxhiCM40bSEG+bJM04IdVscix5zsFM4LYOmlJA+s
doYgL1M7dkqfDKj17V8gGgRbHO/RXYv1Ml61u91hd09q8hv8DICPMZATDoSbH4oRBnl3m5gj6gev
PyYHgX4mC68/MyxizpX9RkhNNHlkqzrv7BQsCjST+CMY1eBnk3x8SgBFeKVJs+WAnP/h8vMjzGY5
Iut2hmZdjB7w2IbIPuiQ8b1Zh4/vrTsHU9GIti76QU/qhTRKhBTMRxwyAsTM3x0wGwWdWBJPbSAJ
lh/BMcK8KJGedTRAp8nTlA2PPcXhEpXvauGS4AszzVyVNlJYQ0IlKmMB5kTcYO1uOsaRxgwkbIYE
W48NXeTP97n5Rf/bI01H6Y3kzmKUZDIzbPpUHpgoy8yxvfXyOuy5wFId1NNGdu63XcY/2pEHYN/x
oTeBP7eIq606T5TJcEfdMiDGMnhCky9iYhBQ73u9zID4MtyqDe8/2D+EttrcEETI+6TozgbADe8E
0zAuheYwcYIwC8KMLztonGjenBpJe02iKIHOQi5hEjAgC6xSwUeH0mtRap1h6ZfmEt7E4srkUQhb
WmKanpMOze9eSkN900OtKL+T2y5CeG/4V78jklddMOTt5qOe7efAKrTuQlbhtLMM/PeT0R0KGlEH
LmGELIRmcrO40OqiKIDIX2Oe+16K01IOUr8xzVUMIqfSgGcH3F9MeDsTeMsx2od9DywEjZLi5zs9
9kHyQVU0Miel5Sf1eisBwb3zth6s7Q4CTp2RJVZ6D+7GsKVsJ1FWAGmqC35zLDawekzxoYNY+olT
vvmSWQL8On8unBqgbBpjbv6YEDoZDJJ1G7APrkW2GsRnrYqKnZrfE03zbIEFYPmEf9Kq30caHTO0
DweIRi5Hu6QFrYJ0FU95C4kdiuEffmJfRS3NP2tHz4Ya7K0/8DLATd//JxLswopBcg4MpgFIdJrN
5IAXcuKv6xgAPAgGyku0ikg2wx7qG2P8zECq9YPmPLUv000HH8CQnb/YOycRwu3WIfReAygMETTt
46lPQZEHRnza2cQ0pjg5jWEe1fLvx7vQEOnHsPiv3voyj4DCqy/vO/S8ORs2K/ozFylWCcAWZ1Is
5dOoiPW56qe9BhydjBt3V40suSPuSxZG22l6u+R4W7KINM8dxxYMgk/6aIjoznjTIA6t+fMPcLa+
ET9m7yML0JPxK6HMw9feFPwn9lvLfbGl/bkULf6VzJrMsI5uloxudvTAq61CPrfwc52VxIoeMYd7
mPaN5hBpqp5HdBGrbuA1NBjh24FomX77Hvgxrp/KC4JP32CQ6nywULjFhcmd8gvaN0/wqoI9t68p
NdOQu0mYS4tPTvv5TZ4Lencz5W091yxKGi6zuUgPkPwJCqMCCYOGUYmxHYDVIDt6SuKx3U53Zke3
//ialEyQpreis8bd0vy2jnC3Rj6mxb+iGw7YgqO4SOi2aLgJC3mUkZI8kkEAG/HTNMGU+5z752e2
gCx56vW28Y8ocQGqisPdYJA+Lrva/Gv94iO1BlsXA4WQbciCpP00IETWb2VCd4KNZ27GKlhIxKSF
BHDv9HrKyhBd/LhoX4NawxfJaOMdBThHO2fAKZdc0hs84oHfW134J/J9TBbogvI6DmBPaDuB6WnY
FTytftiTM4tkO/bqhWZpAH5tx0MWfGQqbu2C6an6yCMMsFnEVBBQ4iDysA9iOnCDJqyXHYSInVNZ
zTZL26ZA4ionc3V4SaJOXm72wdZXmMqAaruOLCsQ/SZlI0r8+hjQfJ/Y5c+Mpsk4Ca1FnOIPBqze
F3EgItLVcR1S2YRgnQa6XfQt83w66Hw35HjRQ4E7gxWKMsk/WjhHjJNaCe1u2x05353w1xRAoAqY
Eki8CCnaUWQ7eoMl9sTOtaEoLyD4JZu+ivu9G81029YEEC3diqI25dgrkb5BNTSkzZU/+AVFHrdC
tK4JmUzQMfUg3iRrC0So7tNBPagjKtp5Ok/L4MoXLVZ7nlGRZEuTGHvv9Xr0R0u8rwbaW6dDimY0
Fg8oLVnu348At3/wXAbU2Dd7Yio8Z0QkalnVw5i5IlTST7ZWts9Kp70srZbp90PdHtU3+O2LG7+P
1fjW+hc1ZL+Cc4K+DXKoTr56uaHZqJVd54q5FcLwfPnwWAdDfxl+Nhx6Sk551ZH1gZo3YJ/2JAce
nmex+11096H8n6qQZsTrVK6k5/mBhoiZb+Iu5uHBbFF8Zx/nEG1VgTMSWC8jGgUt7+NRMSYD6vP8
YnvQkBC1J1gq5JlKfT6LpdVf0xQAx7nnECiqatSYL4JSIw8AoFxl5i8Wpdm1gr2gZvKczGK0yBs9
EmPlRueEd2cTHgg+pPKBOOqn3MXpN3Md82zCQbI0d+rHNQiz5vYcKn1SrSthLcqpsGilY70MZRjy
cqs43ynYM4GbeCJopQmeKvEhOIdtJE0gjHw7aOHWmOT9ACOO46wNn1rOgH+0JtHB/NdF+psDFfJw
e4r1yb0MKUs6ciF3J3o0t9W1a4dm1BFLj23OVZ1VNZPcwwXxuWEisyHhDIK+5lWLKAZ2doP63nLC
lUgUFFlIDnqw84lbLzjKWrCsvCu4xwAUqhe1bbzc2dteilnVApCqxKY/ne3L4dzflxBfBeSdkiRr
gTGIpv/6GW3TlSjYsMMG1CerJ6JVUpbt1ugyVPURwU+KPaDtGJVTh2uyvy1eqPVVGfHf7NiM47rn
C2RwazHKWRwNjrCi41D6STwS5OtmhnfONoBsQUq1MIFHaTEIYrjr9SV+D/508tQ5ZauNVxjY1QTQ
0S0dt9QwGzTP3Tpl+4mYFPlllsUwSl5NYtBZsDdDCuRXCB9rRr+9UXzCE/YzBMY2SHKTiaJyOy0n
zqzQ2CUNQDGmFI/ze7jdgu5/69UIIKyzG6zCuAtLAIvX6M6mzFASkBEdkJwI0VZUgpUCHx4snhY2
5zT7gKybLT2DfMvwkCdfRryVQXcPPuzHxfko/l23SCy3Ud2qSF+uIhsymg6rY6jTH5Etuj5agX8B
Iov6skZU/UWefbvZPPR/U4P//VHpq8zuwQfZ4nOapnwmmpBzIyXxbJl9OVxo8j59K2FIHf3AZyQC
rdW9UZLqZIt66j0pgiURg/11Jy16+so94+aTQyYKwJ/atAXN9UCluvxCT+opUD8HZfKCPUIW8qc/
Tezm5/ziaO61TF1IAdDebiqR6LV83DB2mjnQbAvUlRoGnA9bJvObHE4MSF36ihjB0yMgjqwfLjUx
tfv97gY4toeFMZJYxU8GdwlsLMSQ/Wm86aHpO3lNPd91VHNCgZBtkfJxITb8HebptlMFPUvNMyPq
/Yr5XNMASPEhZt2ljiekJDKL+XLnETQ6DwjmUOkFtw4QvPBspJR5OHtC0+U4EmVvghELyWlDk/Mv
+yV64V4TrUZXlP2hKtvief9RWeDYMd7BmBTbcAp9Z2F9rsfqF7DtAPLpas5Ib65qW6L/WKKgXdda
778cNY+zmJlY0AW/AUBtofLAnvB96kb8zq+qLT/qubkFZvlsUjGtOYdL4M33RM2WiXU4icG9FZK3
7D9bRkkrQjbb3ZHo/V61/TZv77EGZpWhPskHBuQb2x2LkkgElB3TpQp+oSDh/7zySLOMptv6WlE1
JpZByYNrl0BQUFG52D8Ts5lhS3wgukcuZ9AX5yhTnlMihspSg3wZdUzzuiCkcoumxCd68oDsgDrW
GbxDqli0Mlq6fCVghJV7KQ50bLnQyYDuzmaIE2O0rW3M8wKOJ3x0hjgqOykw3FYEWhc8d96XJ3DX
xZcbGvK+yYjdfwkdcK8J8wMWBrzGzBDhdMjtkJ6B06KVTERq9X5U1wFzTvK8BVdMDBRSJ5ttDCn3
N78htxj2la+UXtjWuS4X3P5cKqwav/Zk90oZXdffB+VyCmaFQqqhjK1kUDUIRDbWdxtxekz6qj8l
CX1ts+tz2WzZ9CBkNQ8OzR+v+gSNiYrOeb2wdBMPFobd2CnwDlIZ39Nq9lKoPSYjrMrQhr0RNZwr
Ol1Zj6Oqo2zqRsLBNB3PT1DKHlUIU1/nNDnEDme2PSL5aAksL9aaKQJwnDtjzcIlLX/qJrhS4bbh
k8ZDfOhX1tvxT9vc3Dh8I56lAMTDj4Ce+r6HSgWLBPL6WzCCHhCH/YNKaCg2drt0iM7LtWw5+Ues
96RI4ufXlOClhIRvJziWDxhsfqJDhEal5kgbB8Y9ojIVz6SRBYsyiS+CKfDspKRrnNc74MhP9H1E
6qm02c9bWworBdRY96ua/GhwSouce+po16Ss4GMXm8EFtoTn4NFyVpzNBRsDp1en26M0NCdFVYV0
yN04XzZ5czLxwUFMauoq9c4YbWZx5NYm4wlXqhgpq18a0rWj8nl+N83jMPeiU4EEJ0paB1oCWGSL
q5uXYzQg2rSnI0+2pWgtP/kZ/H+OBfD1DEZRejD/oOK4UNvJtKpcZkv9IMRTOTwEl2Ss/p1DAyZ/
KU7As7dfPg4/SKvQtFnhFXxcp/yk3FkXpA8OcRzMSZNzZyFq333JJHLquJAsKGkvlcwEDa1/lIPS
y1H93bjmPqeC3GpWbxrC97bJSryiMpIuQEqFBLS81L61TGG4MVBc7R0b5WZFpAdJS6nhHdC+CrS0
uim3TlVHQYvhMy/XdTSmGZC16i8Wllm+sxxSRTnWG/jS2RhPFtsV0Sk5kKjHtwnGHG6JWVOJ1ZBk
hvamUzXrZboy+Zn8fsvqUt+6t58NwhyOygY9GrUXU7/eQ5znTr10OVLa6XRuHp0aSNu1GplegZ16
Yvecnn73I5N66lXq9eE5ODpNncJYLXD5AxNkgDMdmvTyckYFncRLKdB9mENwDOXklRXI/5NKrcFw
s7wJkC/FBsUy30LnSafHEkKASgnAPEtD2ESb5e3Dgy9Qv8+HlrZ7vl+I+u0lQ6v1fVf2Hi6TGMUV
8kL9VYcNkKZPN+uEcmB0GVGppvsdO5tv7VQHMjkcG4peTPVQnEZxcP7qsjjrm5trGd1CvJ7D5usL
j1ZO4ge+0s2BPc3sACiV4PNAL9QrD5QPer8v+HHK0C4NxKrvFByZJutgGacFcm0cr+5LwnqyrR4q
yN+4sMIQe/XMXVetbj8COddbsndDLh5zZ8BccBXI23rGNKQu79K22ZxBcAMiFaTOBxO4XdmPPQ+O
3ShHrJ+oEhuaupZ8xZPt7Cr5MkRgcGpuuxICg44e1bgODhEKfOL72kJRGO6YidNn74tfO5XzRGV6
Lg4cP6AGlPAHKNCnyU0hqPH5zO7lIsxamBTMvgmnONm5MgL6hvmYNTibPM+Kc/FsJWiGZMKzp079
3w6UVIMyQjO3/CiSV8CIsGYY/gCjKNMRCCAP8DJt/q1pSxEUpmDW/R8G8ODw79Bh+kDr0NO97LsD
2+6F99VCjUiLEppgz7+2G7R9n1gY/Fqe/Snf1T/ZW20PleIdbA59z5KD9QLatRiSFoX5xtbrEvYP
OnkPuKvmkvfy040EGNkjYYQtwH/LMgXMSkr9ooyAA+zUP651LNhBSMG/ALNiv4RmdkRpx2uwdbaO
5VbNDiGnNgF8D1X6EWT1SROt2M2IvPYWiipU4ZZkpASfEsZk2M/Z4Z0C5vHoP5CwlfoUwsfUHy0/
WH2QlAjziPtduEpPUAu9x9R3Sesa2FNGPhDnJooNF8eP52rVv7x1S4rJcu86Da6m9ykYMqIjjgFm
kcjd6xUIapMyM2NUKBhrOpPV5Zxl0ZinprLtGmf3HruQraO/HD6LwprV0PJi0c7Vzc/a3QeHPaJv
PdsTA0AczX9yBqbaVfuYbnSy3y8Acs7WvuZM7GVNgfVCDNrpdejQEHL2SYmmjHHC0rADz5SmHT8N
/Sgod+kjMxhlF0wO5TXpkeh539SYY2vLQM9PzsZdh+caMWdQO13D0iSf1qke9GZPTBa/0wto6rDR
E4f9GzTt6xTFYglfw0LRSfU3eRFKPZ9b9s84TLQq/hvzGV83zasDhnZh8hmVRXbEIilw4+aKaIZ0
RD+ClX5tdu+I7K8OIJTzhSdcv2+70qsfNjQVowFrsRwHLN1VMNFGhJLOTaFi7qUZ1TFPcB+97K2T
lCBp4NLM4qN4EPGSfXqGUo8qENSRgJP2lM5nrRbsxp6nPwpU9kxvZpgZRCV583Spw1VS1azp+ZmF
cSBwk2cdS8T5O2yLjQYx+splCrZKmBUMUMQow+vcladKsuKq6iJPqTKC8/7EpKTYEe+zbzBDuXle
TMBey13Myov0BrShOSjKa7cmjHjgtHpKBCN/wNriyxlb1t76i4s49XicpGTeH6OCckwmAlZnXTca
TubdI6Fc584kSWrUUAXKFDxNYA+wizT4sxQJrF2DfOAuyJ7NcEGYkvvny4afVpgYMDo/e2NEA0+g
K/FP1RImgh5jlyWTY/2Ya2/BQuCKxg2BEjQsFHqZYPm6pUigboouAk7To+zsRkbxtdAAOvAboZis
CzGiIFNHUx7cU5aylwvFrmWfpZzGWEk+2dBQS8mt1xPKq3WCSRtUh8TdBbOdb90O2OuPpM1oIpE4
Aq67rozEd9ERZlhOM7Bl+y246mhE4MsvGcavAAQNbZHyV05k98FTROTJRo80msiGgGO44yMaBZen
7dZEipfaCVITT6M5ub/N2nyPUt/EgtN6hMDbz8tlISDToK68R4/30My+y63bp26/3+OcVVyI02xA
VzsaGd4M/qoYnRtIysvbqf5MX3Ezg6pl84KIpcCtOulGhfbwUZN7mj128z7AIa+Uge0xcWrh0iqw
mv3RKRU/wBi/sQSWGNppe+7cJUGRle4MceS1W3o2bDpSyXUQRhbTHKV0v070n7PMHxGMaOeRTSk6
jx0W3TS0g3PCtfbvHRWayU91yxTJVrFSEAJhDjtriujf22bnIsPzjfJaDOuT7b7BIzbw6ycW84Cv
D73yFzTPxS6n7FedcFtZ0JNoP7tmqRI6GaG+kQTPdwvfeTXWOGCIy7NepU/1uZCGDQBP78P/hSmO
2YB5MSupTTpC5RQ5FeMl8qmqs+s02KfdIKDGj0OTQw8I8/PDfK9WYQpnobMcvxE+3e0FMXjzNhCL
Y9tzOdgsOMwN8gLRABpcaN/l4xOxrsWCsQwrts9VoWsvRZWP6+o7jj6InVSapKKfcqA3rxQdPWya
BIsxknwHoRGUKlguHnwM0ctS7hGUwagCsGxK7+0ABzODEhMyMbWn+lrxSVvL11PgrsTAvc2MNZet
nttIdgsWByZ3rigsnkRfG8yWEFoc6gSk/HTdP3xozCa+QJlhZh00WpjRt6f3q8oNvqKht7hL5yBx
/g840YkqJ2btvWQZBcZlQhqk0INkHLrpGLoXkkWe24v9lavyQOrE5wlYEIw/z2ePACZhRQgzAzVN
6+cmwK/EuHM93pGJVY0Qa2agpSCZoPAEWeNG51Nsz5CyAq/6YB3rZKxM7CoLS6gScdTgmEAYKoiI
h3XOd3uYFMs1Uq0AliYKbI4ywFmNnpF0k+ziTJY5H/eRoc3VqOd7d1V57ZJ7Y8qC+N1QT8ALMXxy
qKDF5BqHKgZ1qbgWod3OU9uO4ccz30L7vcdSA77DJi3i11Wxx44HcwBnaBbzz909+8cJ2+T8QiIB
e5U0HfpTrI4Jg7/RtQILhHUc/PfCNjbYcTJ575Tw0C/RuEYsiS9Df3Isao962S/l1C9/7pUQU92D
IoYgQWgN+fpUeVh+ySGMr6nuc7fGecmoZ2s8xH8LL1SMKt8vFY+e9fPgVC8vXnk55z49H2VFw63x
fh1pR01+j0F01kpBoHFi2JWKbb/jRSSgtPOYnMnJOHTDqwPbwxekW7569f8t804ock/gmBGTO5Ff
K+LlKaHGJMw1hRE+2vZRMxYxPXdQ3duTiFQzfgZmYZnCVlDcgbRgekqS4Ic7fT2RpZV4dFcTwfFu
WJ5b7a448JtauhO/u8NQaVejDrq6oFwLnEDcos2R9Xl6v5rJnsLeZTzSm2U7+z6BqoNlYMX4sc5R
mA9IVxGI8ZvvSNci8ysnoebnAnSYHR7GOcwIU0UfO69UmK5SGazQxneHPeRDzH7OJA5Yhz+X0ufd
WLMZ8UTzYDm1FTLZZc/x5WyPBFTfsK+MaEA/b9OJGTEAyazbCx3kk8Ft3hFghG14TP/fVDNjiTKZ
OCRQEgPr98eDTpdH9cT3DTKnsJLAVDWcYLSta97YkvnM63I5xG2I/OSaFsibXGfDfq7pRmSoRWGG
Pt+XKEYGXUYX6ympXTInMn7q8QVm4nh9ARySKy4TKrQ9BwWzRS4UnMRp1283Az4NRLvZjuMZcQXY
45/N5+JmRrLIgJP3OqkYo8Rr3aeDSAU75t6DOtga4rAw6eYOw+Ann5zAJKSl3c3Ah86Y3JBIbV+Q
pgsNsBWjnGgXcPig3z3rWAHnqneHg5bOZzenXuey7K1JsOrm6gqlH0l0fnWegkamuTIx2ugvT9Jq
ZTGLZLFPk9/3coD/dADC2Pjh3CzfHU6l3qi2/7rtxtOcKoQfvNJRTES7Dmk6Y9VN0dWdUSUu9+0u
EJv9nt4RmNs/IGeA6s/kowaF1TItGy76+RndTojboxp2xkj1ahWnzhrZByv+4YD4kR1NuI3stbN/
WOnsSTlhZpDHaJKkf+CJt1wbIoJML8qR4t2Pz9h3ZVYIxmH3qU2XJ4HSQKycRbCAzW2whZjTsiuy
u3b5dVMXnupSL5dkehlGbqr2yiK18rtBnTaBqmh2cCSkGvtz9tcJDBp0IcvXUabHR6Nv4J7veI+u
7FDxWEOkYSLywgUHnPmK2Wly5Eat0VO5beSgD8HS+LRlirGuawGzxIBYUzzy6CDNz47sYJJ+cI15
hxcclTGS95/PI5ya+9Hq3U6p9oHeVP+1/5YXtHCGG1WCCbhwhf3lFaEuhNMuSwIitCrugyJnWhtq
s1b6neAGxqgHhlCwJ7bnnHdsDZ3kpKOBva7PndoiGQE2YGvmrmpyG5oZYt6zIruXh+GTnT535AXX
cOfgBjHepG2yLZpicKWLdOPZvK1tywYaM4y68Krk7mpd8V1OP7wQaSSlC6RFc1BIR95i+vOlTaB7
B/83CeKGDkfegCBdmgYQWU7OmqxnDTko5qJQOfSs8fb18pSBK527bJXkflQYMIdoMQkYJKdbA0pD
iXJw+k54AoZgHjIhr47mid6MmGejiU8BjJWm+NNceDDT0+YawxVlUPSIqQqvl2HHQicG8p6klqhk
qFgMgsVyrTwO6KRcXRjWBv1ruHflUbfFdGnq7LUQeRAQBZnFn0O+hNBrPUH+qYKHF8A2IoQqxXyB
q+lnsHEklrzhg0YOrbVojM02sjwYIO4e0Y/MhZBpup8MN3b/Gd8PchVdK6rsFjL4zKh8pm5lZcCt
YtuP9v/bm0gxK+PU8aaHY6qBaboVbgbRcjFNNWV0RVfARSxYtm6vtoLJDuIj4jygD0bvF0KpmYmi
JT19fBCYurZnOPp3f8CT9gdElLR/WC4SiBQpeBx3+ycN+h5H6xSmL6OhoCr9ER31/meJbeOjDI4w
LJQ/tyuGi6cc12eBC+cjle5BWDoBn93c2TzkLLCS/KkLdDHUEHVE8GDdIU6Ul4XZ1uz/mljjS3d9
tC71t+7rVtBE7trxj1NcRyg6ESuIePsqlZcEE3gxdH6fJ3kNPVZtTDG41fOxerDenleYJfzR0JlM
qw327QAwxCNq9OO7w3pTKirF55DxoVYLIBShMCe/OYl8vvrV8HzTotI0o1EnEAsf0Be2olwvI6Hr
BnAyhkw0yC3+GRxYPykD7jI++EDL4yHaYSXZKrHUl69PfbsdgicrFzTSY5i7GKDrYAPEPiVE7TJ+
X8YnteSKFseerruQg1yAnV0HXgWDQzJvtHcEMBZXdBrhffehMjThSxLZyv4jTQ9N5DfBxweJDhg8
yt/zjytG7Av/l7q3labNUUOH5P2+N3RiUiFjHXvMeeH9AZsqs56k2lAPwTRIhD6q09h5HJ9n5RAU
8gluG+ZjkP9rjADQcO3xAjXd2KZ/ZQY4itSdN3rUjWRYqrJARw+mIKuKkGpXcxOl3vHbjS3HYQ3C
gc9K7gIU+QgnH/z8roA/IjC0+AQ8izxZjvcWo4CCIGA7ECmfJgwFI1TVdaAH4WB+nmQdXHCNhQtS
GkQbCIC3K5/47gAl7LTuE8Y2vN6ZZ3gYR5CTycePE9w4+v5eYi8kMNVUlxYsdfyrKaocRDBWs7Wa
TEAuxbUJ/HOl1UQs6aL8cKuFTT5he2ncfPaMvOFCmDVrfU8a7c8CS+vtwxVovoJBjoMzHXB4aYcx
r33ZNjMRG5a150/Duo5vhw2IGsWJucXahNgC5N//yFevKjQasDkJwOq/Dd4yWlvQau8Z1ofAX8sV
MU7Qey72Uw2yUfUlaO7xGAScDRBFPlZ47Zx53x32kSS5WJbrGjJKppTChl5bqwPtS0xMqGyORuq3
3T23FJWkiNrvYshdW2Tw0TeuD4zxL43bhcmuZDGnixPBmvxTJT6UhOB7tQSD0U7zMPZlWcc9672c
0Rp6bjGR72x6y32d4raYgEdLdXu0n4aLgWTMWYmYcjsLoDWSSxH8YH1RXgvptOHqdW/W8arpSOrz
ms/QZ0DNmLOcpMwtABOlU7142trCmnzJEYHQRy+K1KO7tkMlnrL6MsHhcjx8fYwGUI6nO5C2MDo4
XSjl9z4ABsMoFbowZz3kIwpDl46ZCY9+cwaknS+aDlPFheJRIyK+MniNSK+ahm8YJI7Wc28QT303
3RLgcebVuH+ZG5o+D7BA3tV319m71PM7OB+iVI5An+guB+59SNyDT6ynrLMRUpd5JuYgxj6wFDIw
KoxFtQ79J3ap0MQpYBvEQ0KNRqs9nb6T77lQdl39Ta2V3oqd64+P3KYl8IXZm7nZi4RFuHV3RKcv
cPbzVsBjVBiEnHjM98oKjePA/RM/d3SZeaDh0qqOJm863uuOKm6lPKZojBUNC5ZNSIKBax/YS63f
5J/brbFlzk4ssmuAd6E+mkzqFRfXHj2bMAWZGgX0k0Zqyl8ZBzTry0GkyVi3Q0xEoVMpXVX/leae
Hwadt65ww3VywKqSA0cbexmfwgsqAMJ49m73dqQ+kfBB0CUE3qJnEsnYz8Z6IKFcs18VqrYxTfkq
PaYGYPVJmV6Djf1vbqAirY4oHnBDF8yG5y/rfguUNS0733YH4ZOC0t8U0GgO05cJBl/lm3ORrVda
Zmb8R3BZ/R2eUpJBLSOCWF80GOCYJxcvQ/YZVpUsHi2NevE7sfGD0+qEO2uEjHIEnu84h1NePmxf
QgHp40EN/oKI2epycSEkC+AJxFSVWM3CpBVEZsZNAni6vRg9/fkHZloGJqZ7WZHMDQAD2L2PpVQF
914230HDCp069Wc1In4zaeVgg/jqF4WkNuzNOk1jdte/LiKgvi3Nd5QZYuU/cxNppVaTofDOh8bN
lPAoGIXspent83HVnbzWUBQvjQ7PqIRkJyswtUdnBhdDOitvn7f35AN3yzvR9E5WZDztzPHNDMDE
WXY17CLtQwAF/Eya1fQBZ4fmVskE4JkWPNczbHP8g9A/7xlNwSI7MG6d6XGgCTacIGvBbO3gLYJM
U8Mn6hce/cv681ifXPxoOdMAwqOgXYZLeQgzYQc1SIf4021yTTIrPIIhMMMgEoUVxoeuejKrPGQ6
5b3I+R2d03Zmn7ZiG/wHtkSrNG68aT4Sg0Q1bMQuQrXjugDhluXzY+uMajocDUOvy5MIXKAGS5v7
fXlfu5pn7KyciJqVfeUg5pW9Ecsi+cK1kdKrK+6TYd9Gb+Zd7JxXTEr3VV+A7PW/THPB1RzBWDym
HVhVJfenoS0ONrXikT3FdLKtBnMNUV+OAviC2P+aFFEMT1DZ9mlGLTeomIMnEsM1PLVdN9ZxxUsO
QgZueAVQLAG9+OI5+yTR+KSbkB5xkOvxrMPWG5tSA2OFDQ6wwhmsVw0h5WB6u9+BwfYnctSYMxPa
G63V+azy/j1FfAN4/nbCwcetG2W3Aen2QAM9LCsV1KnW42JA78BOPxtuHgWtNNu61D87Fvww6a+Q
3/dSqTMQjX1osOftUa3JOeaArkcQORqcY2DNvgtHq5Zl1ZnTxEd3una4NID3StcUuCYFm6en84ib
Qs61qX+uaC5gqowhrRUxhSpiBKB2y6tmh3oVG/BBPri2vtA5WoZOvXNf2KOsvzJi/g6Rlmb7Xcxw
m8ohg/M9dq8NVtwPjfBC2n5MZdGOrvAHYtaB1eu1QwLRc7FIZpqoQ40aN+TVyUSz+/88v0RrKT+2
piKhGA30M+6fJws3Wl6ediTmioqSUcepR6449wejoY64LTQfEq6oYhcH+EXiKY07nkkoDmRIKhNy
/NO2B2eZoN0lXncfxSoJX882lQntjFJM0T7z1VaxxyNJL7IYFRGcdTgiCYqb6iiaMTAiorDpnSZp
olX6xK0tCYdJVlVjKKcaxNPcF3G5LEoG+lp/tg4T69XzECkJrL9qRGZiLWDoyoRzoqwC38ZpxWrj
XMSapwH24mdOLcgw1+ULNO+dI/w0ZGxiuSmtYIvcN9vWGLcdl4v47E3z59B7PDeLuqWN1FBuNsR5
ufybE8SmfuHdKIeBhTiBLQ+UCexL4hjfAmLADWxvj0yQU3OBoDx1mHRnZMBUUO1mmfT8M+IwoJ+1
xMOB5SOSTolyM831wMmt6I6acqkAn2idXlk1KI7Fnq4ixOpVTPoPcq/f2AT2jCeKCApRsxZNUron
N521qifrX9z+savx9Um3BoNo0XgbXZR0fj4ETq9QazPXhRfMK7WSU5AruX8bzbyv6ZkvRJVifmDC
SRv51x92cwcGzGa2tSQiWqFLUdyuJxgt6bHluoYKMku6UKOy+YrqgdKaT+6lP3n6txMW2sfWGg3o
jOa/jxtAwumn3PMxSwCh5ZSlHsWqrghwIjKS2zhthKzKFiiryfSkAWxH0huBBaUaSYgK0V0erVbt
xcc99gnzcChtf6vZcS6UiNMLT7QQVFz01atv1Kx4hI/1q9CbvSXgz6DOH+Iy65VMoa+CdZn0SjdR
kPbPSdCzibaUp6L2ydb+lS6cgB7l1KrWlhrLIU26k3Nfsfaf+xQqepCl3/00dHWt2GdShkKNZ9yP
3YeSQeCp22y3uVMvb7aBPTvDI56zIROuZGD2DQNHtcXZc/2YrOc8eDH+8JY3FZGHM7MSczfSQy2j
KCdMOd069lMBhFS8A4/E8BSae4VCshUSXBA6KDmr9pIFlH9NObxJVK++hzcNNVUhCPVEQkg1Oom9
Q67MLK7utp0VSBibRH9yUqOfK93M4SNFilbEwP49gUuaJ3scAXvtlQYBujcVBikDxmF3Nl7v2h8M
1KtFTda5ImfDtMiE6/94nypnCDyYkGPQ7ma+uF/uMua3cclPaXT2vvb2+KBPFVsWlGkCwYNKVg6K
9jBG8qEqmX7nscbAXMMbjRBjfmkV0G2dXHMCDyn34BztHeol3R9CAfbVJcxJKPq/xd19DIf2QJU+
G4MZW2u/b0Ho1pCnsIVa+AxQA8Dz2FxeNLqFwcl15CO2QbvUpHYSawBzjlFrEjHfslnbyMVwNcAn
VFk1X0TSFC1aKIX+vNdRwXGm0j9GA16alpda/F6/Boc2R/Qa4Ic0YttxSruRCzEeCfHaTlJrQVB0
atrRLNv9oY3eSYSxqwJWQrOeHdL9zx5IJMohJno6AryQBrEvA7lYF1nl5Ug7QvEs+mzyg/q52Gqg
tmSHy9tKd6QsWUC/Kah4qnQr2lbGXyUsVrcuLqn5i6kTgaLZc+Ty5XEdueXOfaMSSbCbkDO1uYEb
npO66k1BRlkUsd++BI3DrpaLKFT1Ij53LKDZQJ3mYtQcgzG/VEcitLsGiCKe/luw1+7o4X5CO3Dp
X3rHUTgZbg939UHQzjGiWo5UCWy95svWv78I4RtAYfntfOyh2iPZPasgQub1miaNmRn8Vk5JnZXD
vIl8/cxoW0MiXLT07a+HBaCuGkj2NSZ3wi4aIGEBsEJn9gCDV+HGWREmHV6rAugjNLgLI+Lw3Bad
ImQfoFg8Fa8OA1W94Sevorz+proMse4Ky+bnDKX4GWFu/GIwRolbj5TLmD6FfzGQqbOTeSNaOOD8
gg59FHsnjCBMTnZfVGeEReS1OxbBobSWbzujKOhDx9p058R4dTqE8A42g5G2CF/hGneQcJskoyFT
hpqy7vya0JNCSNHPAfjmNLhOlVpUrJfJXtK7h/YHDYQuUznJ0HEyPn/ipAbTVShNS8c2Rr8Yc8LE
cru6YOXXnmFg1DNGN4OjyIitGrNLktIIHFBJzFeZ6dQZl3qMB1BQyJ3u2aXCQgUWo3W+yLUjy4qG
a4B5rN8eL/LBnSVY7ZpBMZiOFMKiBTB82KwqrErl6mk5ypKop+Q73KrJPJuFyQ4JzrCBeFHeTu3X
R7m5A0IcN7LY2n98XL0M9Ee1/ax1TCifpJnmcNLyGMKWPpuWUffCb5mAzPB3FtRUD/PTDIhK7bON
WkPKX78DrAzzNu4S92yFuQSnPD+LunG7d1aY+7K8gQky9e3XfMZ/VxnX00XbVGJ304kWQdDH8sTO
KNaEWlcWXH72IJjtIjqvJ/tFJ0mUYCsSHS9Yf23uTjZI5CjVfuDr3jGNPY3ChF63F75ZS5TDnz7u
nUnCzOpYJ8zgeWK7EA/adfFKdYx5eystiPoOs/eSgE/H/mDE5kflIaAj6bhGrDemvia9yLoC03jJ
m0ZlOlFFkLDY72GvuMH3YSoyOHHFhylWZm+m9qgb+d+/9GWfPqO5FOCH3bB+//0/HmGfsug6qpPH
jD5oOvw9h7iaA5lGlCottIL4pVro1fq2XVlQZoJaqZYx0btY3wp1wg+Wh9u3RiGXpBUzedUueKfH
PHD8NPP9iSbYRDgR/AStd61DNlRiM1bdYHMA2K7tsmxA4tucUkzhZGeSeQARan4NC7lTSiqyq5BD
jjZBgrJbzgxT4EbHWzjK5Zn4DzTk5/bFc+eXdL9DB9a1ZI4oFXB10KoZQrwq6povS5RIxnnm2n46
DPPRdHUFRh9CqmQLL1qlIJiKQcss8D/c7i4OLs5Dr+UvvcMxIoWnyBLALBN79oWX3HJ94Ck/xus0
liNG8w7i5ljdgTfx0MPhwxCRJknW63rHZLm0bqoxgpoBKG3YKnwG05Gyqj5FlqAzX7BPoOo9/e/f
t3uA/FPrqj7FSAwe4RyJ0D0ZFGOIq18SvA6PucvI9WC6jCb8HWeXaOXlaZnX7esABFJq+raxRZY2
d8S/W7lHoA86qvKyGpcVMYgve/A4BwQDKWj20PoYrmo+RTcZALUlxugErgg6AZr4TmzECR1wtrI2
qo90wnYjuxEjBWF/yP4uoMxL063oyQ3OPxXrxQ4JthC2ScNt1FifYeOqKQ3n4S3JLJV6XDzkDI/v
NqIS327pojNACEy33jkA1HSinsYwzF38tWUCLj5kFpxQ4vwTFq9Y1jaRFYoQKKzzwuANzAA5Ssjk
sbGWYYy+Va9Oxl0M0vtBxvLlW/kXLP6TFOePaRWgi86PUdGQ9grzBDbVAF9ho9N4iJZMEWhIWtSA
Q4T+HBrR2Ahw05oHhAG3x/WI5c3RKw8GVSzZHRKG9kax9HfnjVv3MOevSMi5aYk/iq/g9kUrYQoJ
LgTFEC1z53KTKqKJ1PjrNmthwpQlNHUWZ8/q54higQB5D4ZCdbk/EaXgu2TGOUDbPVXzYPMWA9AV
2TnqdyC+M03MCuDx9mXi4xSHcQ4sfSo1D0ZHqqFVYH6t2Z2pLJVQccFfADlE54phh1yZng/KAavb
unEDH6FtuWc3y7t7idvxF2ATAnn8oVDc3uh7uyDfsGPZ+JuPiv/71qoZ5nlHzvXg03jVP5Uzkh3o
3YmRbMt7DKx0ZmqNMVwQ1imTmXz+Zl7xLGfkq4udATIX4nWCHD9nx+X68uCG0sRio6ZNYMw+m/42
gE4Cpk1afwrnD5MKoeSKK1eZU2p7RfJshmtzHnP4ROccBQBDVSSKcWKkzKd0dLlM6p5jG3+xHS72
OlWL8PFMNtvPMB7esxlT0tSVJjs2/nX96IJ/lGYk5J9L5xHzPyKXXYkJl1pauZK68pAhIxVYmIeK
PfZxpNYSFqM/wSDWx5wMN4Sjq/syY6bWIZ66GTAKXbhzhPXNsSjd2uwhUP4RO5/SzmDexwphfBUz
o4tE+ju5i428aI9HsKcP92DziOOgeKFF/ORrFoLcoNKEnvoFt7er+LuQYzEFGmbw6nH7iiQki2B2
FiSysBmOBfyAmfQGpFflAz7PNDzJhXBnpfjNR0cwgHZaNS9uKPbnhxk5kJTIKBtvJfB9nMDJ2Tuu
JMhiRuPTizUxPTKRYX42s3JzuOr3vRxedMOSSg/UPROYkTw6irpHm6Kc6K97NeUcP13J6Q36sd8+
+CuKjVqieQTmw6q4RID51UyCxeM8ajvyOtQBnlGVPNFoY/PtmOSJe/kq6ezex8HMZspRsOG4hVJ5
nov810n68WHJr0G8Cbu0fw+EXxQmzpW1SKDRFRiuWRHjPU50il48qtEcuBc8R04aTKYZxyzPwN/T
tfckG6sHCR0N939gAfkCIZF1NwDP6Uic9+XVuI5Tm3N5hanul1HX1WEvdcVdcwxMH9GjhmcjH9V9
tT+xsyw5Yqr02MUunKPj8cXeHmlgT7LMxgEGTD/y8tqACqX0DHED/VXu7qSgC94dSV2zTd1smf6Y
3ChV1yXDdoHAV1eLHF4vbpBOz9wMcIPlN6zmwmACVyAWusSzaQHreLGE0a+nwzfQD0YtjebdrgQS
EDAPT6IzHnyLbEUrALoc+nRR/UmsoN1diu1GWn+zeFZQm0gZmYaf2d7jxYd2QCQ9um3WqMR+Xeel
khKUlA/x7DePcra6tJTyq0gnXKbl1GTNcVVdU7J235Hwql567b6G2z3fHxjNAmK8uSbBgF3yzyED
6/GIWZPtCkyVGAjyrDXKrp2HwA+yjHRYHL24ZLDo8N/xNTQgd2xPoAd56J549wXtUBqJDmgKAklg
obRkBVdjCSYXQExBqlddN8wGmayLvs4d30bYGUSy4UqugDsAjpBlqQpfPa2di/Hg5TQaIk3I85yk
mkt8FpXONxa0KsInOmSRsF+TD3/Pb2680ozufDm//xjeGp3F9u3igCLyvKKllAwDUvkvDrx/OnkL
b5gQ8O/QsDy8fG31N7b27eii16x3aSHwpa0KtAT+SDVaoH3iC/DuHVi//5dWVVoiHLcSA/0PvMeO
BN7MC52H3OX1G+eIfZ5K5kCPoVx2x+BgrdW9EEAto1LvOsFKWHqQb8JP16m+1e87bmez5a2W+Eau
vZ0BELsabaaqEauVKmyzdICKwTL2wltUXkSSyptLy1ajPA3zHMELzKikXE936LUt8T0n+6nHc1Ec
3r+Srgt/LLdxsW76dDzW7dTg0Cm2dkBSv/y/okox4M5e+Oitn7hnet25xXdFq8mIqS4GNuAuXEjg
SFmoGwZx8rF3AkqdSSFP6n+BgM9h8HTh5ZrkOHWXf5+m8rNzMdPdfOlcXUi/HLuBYrGLmGpqN44m
KSbjF4WMl8sUjh4etkrcnPt6U1M3r+TxbETa9F3lWSMyoNq3DgdiAE9XvGokIs9prSi1R+LkQPH8
O70GKOzUWDWtZLP9rcKMnf85yCh4L2IgGyDoWnEl+l77o3oJCRdBZfONst0CsUlM1kObHvo/7zG6
Ll5QPIbn2L7LmR60kiIlBJ8DPHhtWCn80lVwrsEKXJGM/hCMAojm1eB2qV96QxQnXF5wo4edA5I2
30yfQ79MJWxKptDlQ/9CoFxJzgV68tTJnJBNCviipzok8f3Ukd4BqBJOw1OhHBYkP+hB93Xjk9qe
ePbZ3Ewz47BC+uRl/xhAOrwv9rSjPHHWF2I6zHdJGiIp1ZGv1d/Hg2nbnDY/ZpaY7TtxmkP5ZZF7
Mln/BsQ7HkEDsNjp9hG59x/V1JpaZAYmag3xsBf4FfxXa/Clf/ZVzcTV9+r6EznlKNXZerTNlsXb
cb0HkBsAl8rPFNBaYbkb4GiSqUsIncGhP+YFdIfjUCTXsD5C8v3PDJicRnBd0qYKBTz55RN071vo
mqHuTfTMaacJDnIH8jslXGtwNAyQaPVcIQDCzP5GXgXysdvTXVdU+FESdDcL9onE4iMhl+m+ZbPP
llg3qGSlE0LfPZn96ii721gU2BSljnHESIpXjjnLkwsrjicnBCVKFgZvE1Yj/sxxPI8rZQwywrIA
+G9SqW7gQBYExbfoA/5OOgYSV2KBQ/8lVIkwgUVcllhRvjEtE70KUG87tt76iFj36JSLGewIyKVg
nFWvl3+jzJYieT0A/uOgvZ7spEHJbtuKs6NGIhEZsDaBuPQzC+811eho/8JtT9GXjNOogZS4VhMn
CbxhA6qz2Y+v/najdMqvNDdIe7nzEUEd+GKBiCGeGwAqGKryurLPUZXgxNXXnUYoqQ9AdKf+P9y/
I3gTywTp6gaj0vrU/bcMwWLkhWtLwQXSQ2TYVF2yj/ooD2ma7otd07MHLS3+jaDBiLBU7vHALxBK
MTa1bCbDCGQsijlVsg9Yk2koExKA67GaAgrVOoWPafiFYejlBUxWD4OwFOxWIr4++8RITlYhfFkC
sGY00m7lN7gqmw1PFlHgLOECBV/74ouu6TSFW8nT9APo2CXJlPjFbrkF8ApmInnKpCYt6a+3QLzT
Gqgn/j1KuhkzneBHQySqlw5I43vvv00/7cmD446asYwzhJxSKh6+jNECjCd3m1CzY2D3JOAvxEyt
LwjSEimVEBnYu06YtYPxjExsWh6YduJGihd1kOv1xlwRavg7jOvp0jB5X0K+P3yXj1dCMN2cj8EJ
yFofNQD8CjqF2eUA/ue3s58zpuHA90hxdNLTvyjrqZsaSngBPmAK4uH1fsElLrbeLeDpMMBfk3si
64uw8IvHdSxVylu3PJ6YrDUImNTAFN5W0IzWri25YJk0duB0TkDz7MekUw8PgQKYBRXuzXEdRRTH
Cby7VfCJal4R6F93/t+mBhi2ml7T4lwMujGnZhXh86JUr0MksmOWUDFBIf0L16pnI58PIBXelwJz
WAh0FhRth7lNHYVnzF2O68aC851QYEFC/qfF9pH4Qa0PJJMqfqXt7vmwVU451kcIOmoV3mQly+C3
+BTxAI1yhZT0Sjq1PzZUIMX0uowxWcPAYS8VN5od7LI0+57wDuoKPWCpq1bfC2bSzUG/wKs4LBxK
SsCYkkZl14QaaZt9JPsxzuWgvIuwKiWL4+4gXELqgOJgbh2GLxBXbFvvgke0PpzC+gLdVSPzr4AT
pVZRzAgP6tCWgyfrC0XsCciJeV+lOiQkUXQY0hSQeLbqHFdF8BU5fNSpzZ+vXoEAc7x2jkjPBpT2
yLYqkwxOFLYOCJeXbDD8gVakyB0ezXJ8MUEB6ETUe5yOo63us/7j2mxojzVzEGqbGN0YrQlF24hc
ZsPM5LTv7gwwxEATXPuZWKHwtt75ZOgDHINxcu//oAHrQavALdYp35+Gqg+T4GnBnpsumMERcBGY
V2/yEAyj5B1R39fsQS+Fb2r75X46upt1XBcs4JoGrpDL8jOm9/o7arIQzZ/hTZbZw5QGNvplNae+
U6EEGhWfViRt02lCcjiPatlLlAYQVyQu9nRw4kfPRowJwQlXug4LczFX1KlTSkjiRzZpADFdL53R
BACNve1hnRxeACifMle5SMeW372pD3KkWpSFkC4RcJ9mupdRixbAUf1bg9ru0issccptO+u6Wu5s
nCWoQFiETs34Yv+4WREud19wBQlnfBusPv/18vL+1To49HVc4RiTsBIF7JriFfXxIMYbfAEWzxqx
JdfSiWdL75bk0fpCIq60TCshDJ3Cs8qpwZvSRB4kRoYbvpU5dYIV2Fq4mVEDPDRdttRJZ0C+aSp2
3PQIFwu5M1lYS6WwHTzDVCZLL370TNub3amuQM2J8L6w1b6MrGxnr3FfLoLvw1yJmYjlbdv/mMBf
X4RbtvpsTNGtWgiaL3h5fhb9tM0EAM2bhWJ8MJivarci8egvGqCKsCwx2KNcPXWlFjZ181pkM6rr
szBeNjZ+mIt4raRPtNiUffaoBPsYNAhZl8NlWoK+q3ASRjgizUS6MMlG3akIYR2enDA54W6myqem
fZ3AKF4oNaaPk/vheF/t+Xh4DfGPJqOxkDJDqI/Ak3yNiPslV4/kL83wGO4frspfEbYvJnRQozTd
KDJLNcNJasGYYVwV1lKBVWjpajcmJr8OTGe+FCf8PcIOgMOdsWE7+CpBNpNhPdtG6Z74UWo0pgrm
oOkYP+pmX8S1sYbsExEwSegm6E0zRXzCwDgIR2SlfDQQs9wUmIVp2rj7RnUhVePfGQA7NXraZ4cL
vn2CY5gjt8+f7yguz0F8AEP662qMlQ7hUM+cH+RTxidlrcWer3wQZICBsDHszQrCSG7T9JACtD1V
mGyQZ7Lbe9bT2z2LSc5f52ifPuHjQJRhrM/6nrgt+rbLCV8JkcXd4drBsIlECOCMDrGqk+UKcA2p
Fy58GWrwwAN41pSZNUYJZwffQRAsKFuLk8rXmodFaNTf8yN0kvQEdmDyssDZQ2twD/CnUXLA59a1
+G8HNAPuolM1Wh6pV3vjCajvpKQhS4DpM1UqeWM94Zt2hrvF7OexcySgnmxO0cryU9/fVEiuBCiS
pmR71u3Ib48tVaMJU97ywTNgDL9tejYuGGdC2cgyIw91bSgM4JkQjxkk7WoUB8VXT+rUbvk8RxTz
LEtZuNgqZ2uVSDwjfWKyF/rzmJdB5MVtVmd8u0ubFgzO8KEkY8qnHpACmZJQeBP0S8L7fZv3pIOs
46tzvXOR4nbL5g9mE7FzKZmcJhRZDefDbSZlhE/7nBOLR7yQ2eujwdCJdU9gzH5IkVGIubr+t7cz
FsMyahh9MZ0qjPWKk5z9OjY5o2D77T3zhUISSD/699VDJzjk1f3KSA4SVs8Wj7hCFQI+I/7eA/Js
vVI4nWpl03QEjzmjO25/KuaSuTlRgRVw+df9HSFGIq0hs5M3wMbKZusB1ihN3sUOE2asq04r31Ol
eUVXlNwj3tsdBfPin54BP19i7Z/XSlyGV4E2kKhLzM1QpIg3SseDEttBA3VyldFEJs5BTgV7ycQa
ZNNE1hRmV3ayxvSbOE67dgwxytvmNU6TdCG/EGPrvQsMjdauwalnnlrWbF1UHwYMphBwBfjpFHNH
NF5ZXSqId+DNflbjET4GTz2HQCGMctd9hPbZbFdIS+9uXuR3vK9OgoyeE05+8QP/sfB4OrjkQ5ci
/YV+HB+LWRNS0oXnYe8FiRNXAt1Z8KAP1MOOVmP0ZLs4xHXqWqAOIlOmSpOc8A/7QWyub/YgR5hQ
lsGL80HeQF8y6LktPIblnpxkaVddXh8h3govSS1QqQGBCWMGPRgASdF6npKmEJt52xfO9zVearZW
cyMDyRTeu7XIUwJipP8x6u12NpyF++MvfO2dpWfrxxYM/NItVICpsNL1fELth04us2iyYy6CBCMI
9GN+Q4JZVCCU1LWebuOFg9c9FL+tqFNuVcTL+CszlecM0dt901wbabqsgr7gQyRGm9fPTGfbGMBi
JlNcrYYIc2CmdK8VQM7don5qEmgqPSz6+QSTJZ3u/DOfTOUwdCaXMj4Mq/qCDNblYq1gNnqi3CpO
DtKRaHMM81J+I3KcgVps5ev/V0rDLOPk7c3FCNPYMw0fN8iWdVfx1Gz/SavdlqUB0cUfVeKFe9xK
O90XPwdw+76A9aM1qTTAIY596kaVixsxU9flOO5zOkV1yOYh1Vk5ux9mF7M0DZC0QUGwi7KC0HM8
ywSkDhHk8B+KUP9UlwWwJ6oYZFTfLT//7w5DmH8N6fBu68c+C1YvsY3MWrhVYi/JhN3AtA+KcWXx
M11bic5dKQVE/VNb5s+Ouaz/1N3kI+wUiOIZ3QHzAEcAvEHYyBafg8lf+TIj5wxCeA3y+cmix56p
NA426L+sp9PPa1WIzkrGexndN3FmTszSIaeFM6aUqznL2lStKdR4s83aLlGJSY0iOD/X1jz5BxVb
2+iHDzEkkyww9TnA4FvvzUd4aNBxC7iouUePSv7HdbQ5R5PC3LO3qgPLEFcbxiSKaEXQwj62kN7b
EVrpsv2Dd485GiyHCqjx03Uast0DBFQ5t+tgmlkVyIlnMCyn/f4RbRB/7M8fXRKs0Dkcy2NmQ5Rm
uYZ0ylz6g5PZOhP45WXB8lfNJ8WiuCnt80XjP6+DU3w7hcQCzaDeBj5+m1+5XmEEPnFEqfMxh3aI
ZvwnmrVZPSQrXHmZZH4kfABuEHrbwzHDiC0unr4nxXE30jexNjbG5wcNrMq3+9QEgz0btLy6Takg
4P4uTbUUO8Mh786WzG1gnlw2xf36QrEIyzt+KonRVYXx5rat8b6zYXNToMrE0AC4NeZeju4+ettU
pEThRrr9GTLkAASq2x0xfZkOAgNm00Nh8oqLr8ymo2Y4D9IZVADPfsxu8RTEN/yvQcA5ySmXmHlg
SPbynVctg8ZfF7Y/vQ4f65TN0dbQu4VXTBMHDjqdAg4lCpo2bHakyrA57NjQ9jrFvIfmlqGcT/DB
s6fhu3grMdssib2ehMEHNY5t7es7EIQOLNJaPo59EgW+3nFAK0kBdJZtB7wWg/vIM8Dea9k0i8jZ
TL+w5NpgwJvLtyGCvhhXGoGadrz6YEfroMtuTBQg7ZyAr6Tu52I9bM1VF8LJ8ZPlbvEiODQeUHAQ
AcSsvkaIAnese8ZqZ1Bn7lZNE4qfAEroc854W5g2onrKXoctsSTHhlro43/BLeY4BhmE8CHOJTel
KORX4I6mb1An9ToHZQiubi8r+RsEA45ZzNyAmmhOLoB5HJhz9IGZGFSMxjbI3MnJqBN8Vwr2TTsx
NOt/dyHT8XyBC4E0CU7X7wwKYw3AzX4agUJDB2Cz3dnAKi744RCvjh6+TOtdF8vsJ+tT9BDoA9yi
mHIXzlAFSkVYnDdDisRTlGLX6nsa93dG7PLzNK3Qk1X9OTuaIc+H67ddWqymGkNhgfu87hjVjxHc
hG28gFV0b4Wvuox13PjJARJv4Dp0NnY8oESqwl2kGGS4St6ZJkWiILJF69m/2RLTV/+wUc3G5Ua6
272VQ7XIaCs/4MLdc1U9T5Etf3moymehtrYV3JmC4/ZE1aq2m5nGslkkGQ8aSpvIiDMH4wtTQGTf
7qtqjTSGUPFPh/fGw8E5ggSPu0OkLl4EYqNUF/f7CdZwM8Gqv4yYsdOeIxDpvSwvUu/fUsp8QRKd
mEiyTnnvUMd8vQHWhFRH+Of3isZVsoFDMgKeZ9w8Nkp68reIWC/0bo4vYva2qbb74JJw3kRCxk81
TorTA270UdjYoRlx8DPjVwSfxB202RHy7AqfPMJqylvopecaV7n6ip3VvRwQuEWndovyBPxXK6Cb
xg97+fzJHdQVfUUqFNo8joVn2JWJXM6sygCKt0ehwkpqPUIg2ixavO5Yn9Dhqmb0DS7BuA9S4mI+
8jPPSjim1bffJBik4qKFjRS5SGmLw611zNbwm3QuCHaFe12kJSK+znoOn/HltS8skQIp9Y5jQdXe
n866kA/tzU+M6OICEiWoe7jpIwjgqqdBP5NkDN2zVmgtMD2J99KtllhhNhTfYqFwgDQ06NzuMOeU
+kzDuET8xHQtzixXBpk1PuTaAxb9lai7bHkWCGx00zaJ94jM4+nW4p63OD+WZ41KJRtJP6EWgQMh
NnxpAXqYx7SGu9iFXpbd5pIwGGtFDpAbz6mSeEEfa9CB7PQ3LdRLba2KEuEjY/6fI1mTyCa5Kr3J
n4MB9WY5+Gosqmy9xST66rdPviGvCuJG46hw/IOkBerxT0OSP6VMR0XL3LGV3XBxfZsWtaiipDZN
3sHcnYu26gRmCD3TM1AtLr9V7WGgW578Y4FjQ10gJ0dOyWzdETY/GGMMXz1uQZCGbhMrfwgARrBu
enmeM2hVxfueNSWFrK0AjEQF7fnAvPd0p9Oedp6CWjHTgQKBZ61YEc6u3Tsxlfqy4napxqr1xtnV
4gz1ZPHSsMFFO4ke9Ptiyo0e+TbRj+4gKbsJ2WIU1ldfOklcor3PsBOzyou8nXqI59X/u36OeJIA
Bt9NGzayBPWcCY1bDfPuilGL9pG9n7+uF1SHzgpUsw/+a59fMqk9HCEY/qAiAepLv1IiNA/Y/m4w
XRwjmegts7z51l7STz87m2qYRRpLQ29vs1jbW29sKY0+AkJdwXegOFc5taCloJX+CjLbBT+FFcnW
gMtINmTod5dcwCkvPQ/pEp6HTLIGLRXfKZ0KujElktiGJdPiiNeyhcT62A5U1Sh0saQ/ks6hrgPD
k5bzoBVfFgR3gPzsAFhKe7qLfHizyB/e6eOT3mtMAaTZTwFp2mPeu/HSCR+E/2WllSmxobnsGPsM
jC45zPeo4F9uspOcuVNvSDQFwnwiRZqGjQ+PisHtXknuwZQbuJJdmWNLropvbsFTuQsmUc2aHpTr
ielkQMiz1VdyITDeLN/oXp4hTWpKqb76nTrg7zvzN0lG4jFQyjQkAK6bgHAjcBMyQf1Z+dzmy2/4
pOUFwkr/XAGYI1pPTZ2lgLUUFhhbYNqw0dJmHPMIcDwO79PiSRmFx0I0yCNh8bbk9jZKvBhsh6qf
3nrUP7aWZPJkg5LVEZTgJ4zK3BS5bYv8GB7QeBBGNSceH7JWb8calPI4Dn1ap51btJEuAxfuyIyz
wTesurT9itTGZrLu7Rlaqbu1bTaR+ztywlLN9KKjvQdwi77wUrhaWorjd2Uq5tCz3t2n6ruuQw63
g0FmgQyTWfP1y1r9XfvX/cC/Zg4TU5SsvkhxAvVHgovp0pPZrkGlqYcu+mc/F34v/HLN3efXyjfi
1N6p/2aMlwHPYq3qeJrLLBTHetlr/9sF1AiJEWF7QB0SapAc3yWbMWkAQxkWZnq5NmJ+tR+lwmkz
jwWO7/lO/lrdKiXDDFATy9hFCrT2vr2QSyH0AIMQ6c5i1l3p90O2/+7OSAuCjaaMPcRTS/jLTLj+
N+knCWhUvG+OcmXIpfMl3U0uor2FVlEgDt1vceddLIncC0fkH6vCbp7TOx5mztnIBo5/vDWgaRtm
WnYn2fNXi7OsRsBuRHObLuusrfeNlpwyEl1borcGMO09m7reB7Ykye/FKggRQGUgFaSQ+qOn8qHz
rvfx3vKNeR4ovr2jBaWIkkm2bU4GbvwCrumr873AbRlBXTrzlSdcV5oxCTLIVELIm/hd7e3rl5tm
ZDa3fWlfT9b+vXjldkSNH29R9ozL5wMihQmA+IKdrWZXXHFDInjBM7en2bGvBL+kHMuDFWJJokM+
gcnPn/DTcCiSl9VGscJ86QGl1H9wM0lMSKhgC6nkTruKykhOSaDQNRBD0CVpvVPmCPGlKgZ79L0y
glgft9v/OFlblz22zFJ+A9+egdyPsEFJ/ZhkZkH0GPzXsXYSYJNGxZbiHuVKBTzu95tWaSshN13h
3Ti7M+gR5EfcUPwq8NWfKTyokKc8i5u+O9n/3kYfcbF1lLubwwej3d+kLdz7It0BuC5oI/5w/Ik/
+QdF7ahLtaNCSv6cREkLM7Vu4JkMvzm6EtYCJBSyeXDl6yq0eWgErboXffGkhKjPs8uiLOwo6HsF
eFB+BXiyPQA+UVBsxJoqVfyUY8lznuUZygqQ/wPG6vfvPM2VLWDD+803rs8tPC3OmPeJtUGVbfHw
X6tFwR1+tJw1J3V6sZhz3TriqdL5WVwbvhr3gGS8N3SRwYUbfCeIC5ueqU2aGRGjabbndDqxnXQx
ededEsz73ssozkItA+7zQiIBSaV/SubtM2v8nHG67AqEWlWVhxSRQ+Uhsyd1Otcci4KbZK6kklHI
8/XTj8hDlpIogKaVpDsUTqCwDlXY3r9Pt7OTIg1vQBZCORJ2yICXDOrhHbA21Th0dHyidVjM76N6
9KG5XddUTUvo5OqzVh5KyuO8CuTeEpquJKpHWgM9rHZV3D57dmklgdcg9x+EnTmylgN+I0lSFkQI
ZFW/hjd0NLFHbzMqKzkdotdafhn3ZiDkkCYt6jxsS6iPJgkhnG06pJ/mMtrKSfvpjdT+kV5LrQ3Z
VSBMah8L1YBmrzFu2f5DBsLuK1rdfHj/Oa5FvmBStloZulUB3YDz8tt3JzblBdiVezWqYOcYiqfY
OABnI6g9RGbd8zb9hAKD+ky/2cE5q1STn5pg9cnoztViYOWkrkkGirxeok5Xb/HzIV+wNZXM8QXQ
d+9PY7BNWjP9t5p8ymvprVsLHlqG9Ernme7gah9As65XLUJB6Ps263Cda92thYnbCYOO6W8vfVTw
lNUdNBNFIqAF8xt0EbhJvJTFeDLhhZcDQAasxPHxMD9Tdc5HDHya9Zls7ku1ofsHDYdXZ+qiMLuN
3u1VmXn5o8tyEGs2W7Y59AMT5EAbn+dMDR6bByu8ENlReKof8yqzjsAP2y6k8E9q+eVaLNE3huuR
VkyJ4YNmLXM3/iInIlfL6b4TymFqYRbKZKeTMd+kFtH3YC3FmR+THKhvToLI3Mh0TYxu7KdoCSLN
5fjaCgNxU2lhwcTSy3duwev0UZJuBd5pjaxHnHPdoh7ruBlBm/q4cttc/rcLub28b8NDEmAvFKuG
nzm/aZVwibh857j+LW8Tv77ITqRIoSuKbD5lqguW110CjdFHrmVPhVvsqJiOe/bj+AMrKATRyutj
N/vGTg8ipbmJ8l+T0eMwbuokoumbEkp2wLOtmy+Wf0Mn2BBIW4yxFbXrZknAanOoIA2QXRhDySOG
QPpv62IG4aq4qTb3dy+OoxY+p7YL+Pmp7yfLMNF2ILE8vtceZ40WwMejHy5zWm+Fa8vkkS/t9oVd
LnhfQ2mCB4K/lGZBn8y8llzlS4fmoLsFhAyzahlVz9B/RPc7Ke7D9/lxsJxAzQ0mJfYG1X6gFSHo
afngI9STYKQIfbc5e6bFSi/cURbPW/XiOKpRggSYkwZyj4XO67ekoj4oUE/3SaV/PD26zgj6Rkro
RmQw/f51I443KhwauViXHuU23K9uA4fr8xG/bafsQ4C7ZDl20Cp67lEvFA0Qqs0bGMNNh8tbjG+G
g1x/w9s/8O338gnRGfeJTBMaOpvAII4ZcAkho1TDDJ7tGB96YumhOSu4YQQlR6zGmpS/lfl/E3nb
a8VGMe7Y5bljOLBqaLPGlYN6gY6CPdFRDfbLJeILTxKkFA/rKarn/VlWrsKb2ZNo9ihWcK+a28FJ
KJaVWG7X0bw/8KJSCXfge8LvBKToQNvmQCPYhFrtyWIqg3NnktDtouk0GcS7ZziB6tbIYmKBGDQf
PcHvv85Op6bAKf6xdlwA4NSE1ZPqDw41NTpHyMjTlJHPebb7aDuGvf3eYJAHRX/E8L0+RraUaY+e
qbPvjbTA4Mb43THi9oJOE5LWcP/jqMQUFjWvx9eRV335H+X9QL0RdpkN86f3tPRxUZ8ibcyUf5iM
yLoYclEGeXEbVIaJ4E1f39mHUrgVaG6cQV15nij8dRnKe80o/UYiuBhX19mZQpLpGF9RC1izO0VQ
PV2HVmQzgEB+p8Y29MbL3KTBuU013c+nFMKMsBuoVQdWjxHkHCMtYU+k3eIPbEjw6YOiMJsfIoCZ
cXs/A5Lq2BFsHxsDk3Z9vk0TFIiKPZIGtlsg8mcz0JegD17e+zawSOR9uDhv7nkEAXr05xlhO97X
BrRMdrmyTOuAgSIuxcgJ4Z34f1diEsMaKV+mvZbJMJu8AgFKyLcRP4d/LinWpSeuMwijkMAVpcRh
iX/N+pngBeRtb3MjNXSuU8LH7LotNPLGt/0F4jVejXS8YuTGIg4/hxkJpTnw/6PDS35dXyecnIfW
51SLBNx/khj5DPNfHOxG5F8crL2qFKkgNwQFy2dWRPTKi4VILxCU/dK+FJq3tj9gbjPS3IQApt+c
bY0v7IdvsP4J//qgbJYcK4F4KrAwYaRwU6voJTBL0JA5ecYauUMU++3owmfEg4joMAlRMlbPB2k+
BJycLjvLFivCddiJtWZAo6MV12lhuC4nXqitXUgb4ceV0dK9R9hpxO8mISgCPtKtK54e3brZJi9C
7Q7/WkBk/WTHmLdQGXk7RfENS3LkW5TQI0zjdUUXPe8aSbE5oJOF4hsWAZxFGp1+b7GadUXzjaCV
jymYQNO2gtiUUXVydKOyzi5C8KD4hF4aV1VVTkLZ/O7GCRs4UprM9p+pjRirmrwgFN1oIAK9AV6v
XlIyKWyC4FFo9gJKsvD6+RtQnNhKiE5rdDQECTTiMYOw3i2Bj2iOYHOWqdT3E4Hdwc1Mc6vGrCKn
Oh08y+x2j+OKGChqctPhEKrNBgehJcHuo6GqX99ar9WQPIqX/8zZVQLvDpMgTb1a4tGkUt6kSWWh
+e5sEu7k1ciuEKlasxiB1Y9yWb9aLSZYVkms06Z6Mpy+3bLKztQifM5boxqBRY3mN8GQARVR48J5
8ZM86rNaBy6i4uhp07ReSvz3XUTvrwnUQ0CrZgZdDzToPo+7a8n6IplWJ11HAP43FAEJicMzWQyV
6/MOg2a2Yn5t7A1e7O51JZeA5pfd5ZoZhCX6U1a5Em9wzRl50PLC4B/fUaHtmAKnKs9wGhf992/v
ZzXCt3ugwvRM3sxmTMrFKsgIpWXHiHZk6d7D6tMdPvwKWlEOBXs9cmi+B1Ft5bpinyRhe3zY7X0v
VjAKB89OQkBiMtye0DJtzYMLAEkR9QYKaqAP7gyezewXV+3SOpS/dpLEbS/lznig3fxtWe4/WmLU
Sk9Cp+ef4C+LduvyQyWS/rrWOBtc3ryfSMemmAAGPCmCPryaLDUnFlfGQ5Yo2z/aM4yeaeaoAMtb
itKcE53jvWkdqahPIs39Jm9APoCHRjc7oe0McGCAJYhC3uF+5o+6zz2J3W0fgILduJ/m0+pcwooV
XuX1WLK3CIbCl5bIozxLHZGGJxv+J7ne2Ty7H6PYdvigiKZy0Iy1D7132vLoVI9lxt7b/A7QIxH7
aG8jMQf4EQrKq/3pit+4ZpvDBTqVTkGXJad7BIEthUQV2uNXehS1rC1ravTP0kBLFzOJWZYrrar9
XvMOzv1pfnIJ+73KbfqoYJ0ePu74ldaaAbARdoiQ9hXKS7aKdhuAO830TJqhs7xwsoYl8Yx0PgV8
TG/jJxlzSoai1wGgx3oHVGvDZsWOu4q1vMk3GUDnimtGOD9z5XUvmrO31VG1ukOwedqYs3UNFNz6
ElYEXDDeLaeJJEl0+TYZxRT3gSwVvsgtsDUrt7LhsfZExss9Bu/6D34yH9cWDnIs/UPDXCsIcZD0
h+lXIR1ElaDSNL/Kv7q6n5y9TGJ4jw2oR3CjPVtMK8MGmF7m0473Q918Pf6T5Id2IMWEb+Y4hTAA
UM4N8KLdz72+hvIjmEmFighOlenH5P+oi0pBnALvcADpfSSiqr/EoDTtO6iDN6RZebj2Qp1PtEjF
cLW6osrjrFJ0JTTqG+kSLF38MJGjevOQcjjXhZwp2qsJl3dEJXqS+gxCboZnCYLrjeOl14Ou2G0j
wwTiXZk7PaldsUd/a0W4JwHWmABiT24Dsi8F+7rw59EiGAbN1ZlhbvIZqwa9n3rCOS2BBqrVkueI
oeFVOPkKQ9n1bVQC9NYyU/5Mtdr+48mmRKQr/+8dEBwvIzbXh5V8JagM97QFMGus5NNSmE+U8mQ3
oVSGiE7EyaM/0ve26whMVjyEfcNxjNwHlQta8FtGZivkpWU18Q1blMXnKPHZeeyVKWdZNSfcn5iS
cgKXUkQZxnOw/rSqF5SiD5aCzyLXzJrgBmL0Cn4eM3fb/NrgK5MW6THCYYw9nLUw8yhIm36Df6YW
S5u+tGwVtI9NrlZuTXSMiPAZJ47eLh4IlNOQsXtVzD8x3fM9K0V1CkSSIfmd9nupEtlZTCPIc2pb
tTA7mqyfXQZn5HONWwGlpicGhdJnyVPgYhHFN7bm7SG+9+JPxit5DjMuCLAVvpET4yiFzXqokETi
oC3ct6qcdEkS+BoPeNg1sa8ekww3NZuchQCoVGQhPptXaXpfA+EWIyh0n2QbXlbvS5zjrIUL9d1k
ixg40SSrvwzDJMMmX2mEhIs4vsS6+miPERl2b7PTU9Lw4KDn4vheSouApeQNNR2fWpccV6fbmpLU
+//avYy1e8lFWXkVXmmpwOqau35EL8eF82GsV+f2X0akrsvbxH+LybNUVzH6Pfue/0eMouQ5jt5e
XywyHo3esTcZyYSIa6fHDAlpck2myfyMMPOSRXOUBX2u+aNgKs25ifdQvGsjwz7z95UeIk6JW2HL
TtVyihT4wZZsQOQTqcpla8trTAcxwGX1+zaYHxLHDEMEV+J8uzXLkCuq9Ry+OHEin4Ph0an0EBCB
nqqRbEaY5SyYdD6MJ7/F5Bdki52wctskSaXv7+n8ZOqvCkSZsEnAa8/3GEvhcccV9wn+nPsCKtAr
TacSIhvi7PUVXzTlT86JyZuNVk4Or8nocgF/VjUCG7Ftx9uCkSgy4xy7RhRZmWwBekrubZAQmiYD
wqmTFy043G01McqhqbTMBZpCWkFTxdL9hEodtyMOKr1fJTs/JNpYSMPWTtHZ0z9ewjW20rTxVcNm
zOcm9wwyhhhukuryjMFs4ZQeBy2NGSh0iccN9VY1zLdf3J5HfiUPkiUui11Yj0SOBjh9UyMuKTHu
4jyMUCsumpJnmPCJAv7ugowe9VOCgZZEs0x6pZdsNt2VDARdn1fDI+T4YCH2RtUkU1J0ZOcjRI1h
9YEXhnop0Jhn97PeHW8jTY8U1gQJMT5IFAcepfLijF2CnhLSlTpiDZvSFHs2+ifxasPeaQ7sShuX
GXXSk5p7GisHKDk5kQ/Gg86ug8C5y0ixnHyGVprYBpS8v5CCxq2MMwUml54pAyk9CXb7PGoB/5S/
fq1hq6TzDneLa+ASLsCbkrrASUOy8C44hrFMFYlz0XLqigphogDy1H3KLzbi704bCyl4P5eKqkQe
U8qeTunfBEtd6t/QnatvrHQy02Zyra0P7jtkBDsePAfNnOjyqlvVjoR67PsRJFfQX+CJpXuGZ3TW
y5txaCM0NnkbFrIo8lT+hyt7/3Ay5xpWvAP5KAh3BTb3cW4eDWlXQFwpXsYxpcRQW2mMeWatX9Ny
xEiSEGOtVEBOJKPaGgy44QIp/TsAs1k9Eh6JxGfWiHQA8R7uomVLiC8mgiVjFoyQGICcvZPBWqmX
zyR3o/l968r7PQXIWRjkvwQJH9+oiPZIiTYhUfg8OoUhVndo/pzH7U6Epsj3VF9sjbK+j67IiJJX
nKMLemp3i8wXU3Of9D9jot6Acy4fDesYqwZHX5gcxtGmJFG+MYboR5zxROxmy5nJ4NgeylbzTMyQ
SRPdXZquILAA3vkPiBcJsAg+0lNYXQ7YRfp1Xj22inKPfXbA02GnNCa3aqaqBaQEt44/bBYoNs2K
8WO+wlqS2ioFKLjzcwGHu6+A6EyKurgrmDWfUImyZzhzAph021I9EhIR6zEbZ0WoZSmciUHT52DK
6P3sgfIrNhy1Yh6bvIonkWPsksc0Xswz4ZSpbd0kSIz/02Rqi6/zL2fxSdkNW4r9FQOKVyVfrIMw
LLV3JxM0UH6+OJbIbUPd9/VAcoKJ+URuoTPJcosjaXRCow3KYVKKFUDsDj1RiywUOCJZ71vOyxGL
5MXH5ciJxUjUWZ9PbxQQALVMQNFaYO8+O24vSw5w61YYTsx3aXGIvPbaPdHLhWDMAbJ7E0yWs6k+
JnDkXJfSCZcAxKh6W4hROPYenRry2abfzdoJaH/cGU97PCICUS/7QUITwpmJeTXKzhACVfbs0Fob
DvBlini39oGE38UU94lKINAYsn7qVwdmSeKb5Fw5eCfhViIJXJbLmPww1qr7BuY9SlRDJ4dtpE4t
Sh9KLg7iC1pTUMhFpmDmZRU8jLuil7+feZE1bXkIOQCmXosGcva/7JHrD/mwrzjuYiCmLm50WIh2
90ohHS/jcWmF0SnfWpvTziCfliCLPC4ZWdgLeNOQYXeZbA1dAt41ah64G9m0VmQU7YnOmDvLtp5K
vvpT8qpBfxn8hsgkXPM8N7HxrUhUiM4Vot5e8vAVZQdw7KCAFWGxmkTpEfPAS6UIx3NqC4XEb+P5
YdgCjfVTtlLndU8YJSk4VTmc9TPoJ8mrLxblK/VwZDPBVe4VubjK/drGdyiHIGGLVrKySMvLcJ7Z
dlUuvb1iFI9H8w2aL0My2W0EmpNQqyce8HglzYfoBQyxiEeDRJaNouyZUpXI4K8MI4SN5Ojf23VP
hWUiBzjDdCMLxjyTzfJLzqRL8YkqCpkp1/HAR3apgqx3ly/ZnSkZIo6nnut66IAR2plPBmikdyY1
IpmU+hrT4hj276CscNjNse/KaxpZlHWXtPECDIf5aytRmHOAHQ3gjWpiC2EYKgL9r2T5FHWUtmkJ
tAOw1M+ZQ4qBqd9YQoQtJnuvF/XHp6Bxet3sAAGOFJ3gP00qOiLYhV+Ccp6ENtifMgtcf+7XbzTu
Igw0q4gMz3cyM9TmDLvAIzs3gjRdajrDoU9DT5ExEeWtVdkPsPdS1QzXi7iOhXjI4GIT+D+TjMp5
eDrexR4YZfOrlGLRDO63LDrHNUovBfYUXtJ8rZQ+MX/NMVuPWuzXoCN1WsnvdU78YQy6soDduNXr
IKBYpKNACswULgzkdydTYVWXXikNnwFMhyMljavd07KadavXHLYu8DyVvudMxgJy9N9XOVOPCJKg
zBX29HxYYwMpjudKSBqlVKUWZl/lg2lJDgMAckfpls55CAJGA8LaL0ICXXoZGTp5Qkmfy58vhpcS
C7VKCKRn0UHmzYRQqWXF81Dk6KoyItHcMzWoSwpwxbMTm9nhwsgAzhvZ/iyENpp6NWoHgBMZAIbJ
9FHqlYS9ZSHd9q93lPHnE32/B5ty24JbMFOaGiTD6QjVbvwF5t/Z0cmneWsM+vnIBUkc8UXb96ek
/izDlGhH4UgeN0FvBxuL1WXqTF15IvzvJjya0AbuPw/RdzNSnPKfJkO7dE4qV2dUzIwTaEAc8TEo
8+6/P9O8rIinq14zINSfl7NdB0A4dgPSckLEi1RzzzlRybrlGt0xI9tJe860S7UnwR78598LonmX
NdJ86RDEKXEwQf/zovjUCrU/TGbSEQkV9UJAYqSFMb+XCY5siVCUNOyNvN8yElNwiiHthg2aU6CN
noii+rsQUrkMxzy6hqLSGNKIIfMqHkPHjFNnBXLQitdcl5Cen2/t7OFEQ8uLq6DQBjCMqNJewjTT
vSOGYtJjodgPu1HwugpV7qbcaOvs0GgmAp61TGr5HD2vZydwyXP0mElOOGL6kw3+Qhw6GD1VPMma
C4j+37BgVX0QYzh69is7FeCXCKQAZrj4Ofy1RadqrtunmYLNDlUZ05qxly+g3uvytT3eHslP5D+3
u0IkNOAwv7ZkpG0W3RSnfB+l1vd4foUVKHPC6NKz6fg3T/cWPWMf9g5S10jaYorPk4EQI5iYLKUY
W0ld5KjB0o1bL3POE/LyT0ERAqyCQmLZt5DznxGBcYTI56qC2e4Ujwn0GXKYbQjG/s7eezzMWaIV
t/9m197YzvUIWuvA4BZAy7SDQDPNjIYm+6d2yLo3d7yKXK0jpL/gweIvdac6YMFLAvnQPwog3XQs
gKGrD6X7wyoNKkwPvN3cmv88uMZ6FnYrawKuBmwpiilsUPoMHEsTAOmWNB6QlbYzy20cpS+Vq1hy
r617ZF+jJErkQsUrZEZbnETlyB/t+jV2lsKcnjQBwP04hr0CkY+l4IIkDo4La4DwSkBifQmY4CY3
FHjPaav5cLnw1pihsnA8SbdVC4Ae3QU0D8Ydw0WbUp6PrwkcSw08fv/hYMsc+Z5V5PMnSU9nd41v
Da/LgOzzh4iRjApbaNvRigV1LNzA4hr+bIs88xXZiV1f8PxFG/sxAErQFrWSBPE5KRouxHNiDbhr
IC6YHJeeexXEDEj4hQYT/6mgHRuWBwcqsT4Sucae+a4v+YdLJDPjSNAgh7GbV7/xyv/E2tfwbc6p
uDRtQmVNIxC7IeSJ9MF0KQ8m9toHD63FF9rFid9BDXNQlYAdqmotBIW2Nhr0rQ2GXeoRS1ZoPbES
ktsmEbi1AxfmRtzHQXMAHyEza/zWGPS0Q57GizyAFiqdpSDw329SvuphDBt3zfzdgpLFnNuU0yzi
XXKQjSmMn8/18L8em4HtYicUNrCrTmS4ZV7nTyDtSX+L0ScVghVIlC+U0MJgHsi5tKfyHJNl9Iuc
1pPpXyJuASEV3YkP3e+qFdZ7uTH+oa83Pl+C0ByGwiqDRERYUQv9ff3pMi5/LPqSgowVyyS53tah
Yc0didzMmobk9fCPESFcQrA1QPtKK3kgmhcPWNiIZ38iCIwTQsBy9tXol+WA0PFZUGnwSh1xp2wi
Nbw5H3oIMT0t4ZkF3WK1Zk3nMd9bCVJMuA70BJZHSYqClHvxg4OH8kPm/Gl6S7Ve3jaY0X9bnfzj
WjFvmax6M+a7gz/rz0eZylx+binDyjs0k4npZQ4taf36bsuHWC9Xjqj9WoOc0tT53qs2lRVd410f
gfSHYLcnxvk+G55KHt/v3MQUDQLPI7GVF8cSCGMibJo3Jv30E5szZcTlDooXYeO1pJilXR+bw6II
5240qK6RoVzu9kHOhUD9w/+ADRziPW6Dq5o1ndg8084hNi85L543FFbiakOqInT3YmLRgseqzewI
hL48sQNovo1hNxYBfSi5tX8NmsDKYUhlATFVsj0mrWlN+Uu0wLAtAzKp8qfN8/6+N/IP+uzKpgAq
jQWgTj1ORBMhnz6TqWgLVkEHMdLMdJ+kpluXr5b3t9Oyqv2xFy8fuwNC3WBXe2L5sDw6x5tJulvT
GxCdraMmA0jng33Oc2We3+jNIbTBY4r/ELLzVAdv0K0FbWPuGm8IDXxVF9N40Wa3ysyk/lneXD3Y
s0CVHd8H9qWDlhqfdvo8v64veO0lySZFlCZ86uUwuWl/bZH2K2DuuLgE9QAClOUy3q3I4kCygiVn
Kvg1LLQz355UDWiUmQcZK+EptcGDajZzxFKI/Q4T6OeW+SGaNQAsYbEJyDwPQqqo2F6KctHqXSpZ
KMblUmZlIoL8jfXxeOVijjHqY2obnpMY4YWMX+TTDs+mP6l1kOSc66reMM2zPaeEuTgFR8KBLsYn
a3TW3BZtd0nLl72SbkIRESMQ+Rl61or92JnvM2fsgBb4mJzhaZvizMH6U89PfvSV0zpGTzojHpxz
2W0lUR3wde/dOQEHtyEIB8e7PiF0HFFCclOsFGwuDp8KSotakQILR72xOynYmM6OJhGvW+3v6ThI
kWiYBbpYjNduK/mxjACchP2MAd12Tx1eZYI/GQlimMNXFU6Ird+MfgqRtr+9zlKqFBMwoRBjrIyL
PELDP87Sm51C4iu/btdr4wzYh7UHzFi9YfXNmaInCMfGJE2XvO4YZwNN5fKzuEwVb1bzXbBrKczy
bV6qJapxZgwkklMtXMMethCZF1UpJ6WrDHyISl5yX8jbHm6DX9evuOMNKz038WG1hgfiIeZsFlq6
/hhAqvTytsOvtVEwnyipcIOR97CP9VebWjlfZlYuzQ1nwZ0EBLoVnUvjPqgXuUFrobYG3HkUjrkf
oU7LWX7f64Xfdw7JhPShSyPq6bEdXCjOXGwZdbWXyPPfMhR5L2AItiCNsl2K3ukkdB8l38jGjhxM
MnQL6FVi0wtUjYVrQ9q4yHF0LWa5PtN1VUROm5j8L7oitv7bZnF1zbY6RbovpV9vtPmINvdXzff9
ENznynPnaCa7rb7mBNKFJOM/eIjqwhLlwoOfB4JlaTAGrErX9GwKiuO/qtfsIMaeUn1ly89ldbJe
yEvYGlQTmI+3afcFIitGuQT5iIhJ0nB8ucETGWFwjbqgcEANgpexJTEfU17pxTqgwvIyc0ZH+4CT
rIKtuMb/zvBd1SxHdz3rDRWASe+CENP4LB2pf3BwhPyTRJwrIpE113xEaNm69YIJ+tPCt5jBn8k5
gqM3+GaJdPgOKJPEUUVRwPWaaYby1rRBqkkwDFmSZMkFF3vkTdWaX3ZPjJ+Z2Qx6A71CUj9i/lPz
8xzF0l0Y5+GcR3NZNCt/+7rAU+s0XqtZt268G/eb3k5Gbd3kf9c3IqM9mJxoPip7H9KL7/APrstn
vVpOmuEHtncwPlvMblLvgdAtvaMmj1QcFiPWLq1lTV0MGFp6zkknb87F9TSZcUj6vIJCE1vl/xdk
ug27KZyTKHdsPy3+nW/wkMnfxv2taaK0I3982fD4EQQL320A1fdM7q5pdBSUeRVai1dWkKWV4hWV
bu2CYUuEKSSbsqr6s5aAz7gstxvSDStXBucQKvefk6ZaG9GmQiq0yhybD79pnDPfulKWNfJYit74
sdirNTQjVU+mLAhvDYxK2YQgd1cVdzkt2zWKOyjqbb/9n2rsYf3agoFOkyJQ6789oTwO/0WTJUP9
GpwNdOWMmiUzOWIhIBWmEYbmDNnUfIhzVRsNEmEsph9Px19oCpFa5GaEViDoYwtjftB+7452j3Y0
5FbkumylMDEbVOmaaebUG3e/6Xuqoo6oI40bGG1htoPihS9yWAOcgiIQuna3CkLxBy1fXoQYdurM
7SgbvuaODtUDYmG4+RvsYHKybMJN6kAJ/2nxx/NDvfuBnevKRG8sxi9Smng2AJ7bsuD+rxLr8UJT
yykN86+vnshZsHg6KNOWMJhB/VHDiedSeKBkNptQvDa2jlLajHqdDOh0g0b8mdQvFh5SlQRWvXyM
Kz5pvNPvdO+5APAjBb8vND9YSXLFZO4ZxtQB+ELBytIStyfleHZHvKFJAc2VI3VFYdjvj3A2luiP
44uMw5mG5kF8u2GwgMeyBsx2P9n/NxwgTQ5a8LyKIOoBr4hp/u0jBZmPlfpDmIv+ud0+Ktmws7d5
fEkBsOQPUSWXZ8ZhyKweDprypg0NlOEXvBNFVMmWuDbx4wQZaC060yOnwZK8Py5fC6MjlFuK0/yg
gCakZFWaal5QBVK1BD5CWXTRKzVhzGqPhpuLPd6oVpFe+9UBQMvOyWwJFU774LN0S7SgVL/TnSDo
AK2wkPmIJ7RsoiCdBrA+VP98B3sZm8dDIu5ykigijoMurcJ6yOQZuLozalRJksH1fjpq0Tfuyinm
S6cNRUdqbjOWKlNABMB1QqaO/3I9/19grqswkKLNN22ELDyGJv7RjV0mHWyj6cl6hwdP1Wx7kNKU
CtuaQhjxiR41myIS3wuOTGKC64Q9dhTm2VRGG80Rk4Aal3OvCZxv7N0C2K8S64AuBObBqaGxFTgS
jMhqOScLxU2XeavXLEwvPCVag+UUCrZpGwASj7yCexruFbxQO+RyYuPwryVDM2bv2qT5Y9cM+wzz
a2g1SJ0eq3qaOrG6KRqGD91ImvdpoAS2RPK/lRwQVAq5xoDv+Jo2tIN7htBaJxEHnhvew4bO5Go9
O3YScMVMRjma4S7TwaK0+ndZWcW0zZWlqGTzdD7atI/fO7k3WmRSCJhcGHTzjopumG6+9kGsJ5Wr
32glvF90YFlfXBM/y44aRnRH8ZDVimCnYUWCJ38vZo8R2oaO6m9ha9tN9RdIbLaNYE/3pOMn48Jw
d0xbJrXzByjg3tuuSOfsHtzpUMT4wYyHCONk+ts0F+RrbnUjQG9EuTeLuLT3bW9yB2T72GBTAoGg
pV7bBYldM9oCsHkHcoZZL03hzseBKIijmy9fhDUJb+QtpDOWTJKJBtqaXU2i6NCCSV5gw65jBg2Q
7g+uMm6hYdM718kN42lpyGfu8NgIzJtZq4xmF2nVQCI1HK7Q2qZthwMyKPSKiwG1aXZ6OAgFoC5d
WvhW6aA5NA6eVDHoZYx2S9CvJWg5HJl/V0p9g9au7qZh8dS9ONQLX2vGh6BuFK9To/lJmzOc8rjX
SRQIlFD3SQa6VQtsC8Ws5FqKAAFAgUDye8P8+h7tYZ+/VDQm4QLzZCPTyDMpehnOF5EiIDfF+XHf
fn29beJnM7zsCQsfq3sRCHczcbaev3YRbwZvKKtIn8PzREKi3hcFx+JXozgDeEkQlJRIH+tUiTTe
Gur5+uNz97TFtcg/CL3gxRJ8tApG9smKFxl6Zf5IROy0x3WaX3MjIZeZRxbJ2SCCAW0TVxq1kKod
VGCDueZsbADWNNqrpNTjCLBOmRlt3/aqNEkds1z/lNc6PpdWAMM6z+MJ4o0X1OSmWtJNlYWApHCX
lj0Z2VU15HSo0fN4235/Qz+MYAoViq/wrl5zkB3BJLM8IXDTLIizIq5Yz8ViAkOrk8289wdZSnDL
Ozd3X8RhqY6O1QpmIySjuP++lBru1bD8wfYE1lJol5qbuLgvawPD/UZhCCq9Fuj+08VWOuQL4Cwx
j8dbqmzg6AzuOla2NZDR3v9D4ifkLVCY2n6UDSH+K1igfqTwynuMHRwnAXyh7qo6k9Dz4WHLgMbc
o4e26IYh26UHBbn/DU+0I3J4VnGbg5Qp7YFAi8a+NgU9FRCHspm3T/DFWXYRG/MmliQa4HcLJNcr
QZJp7+toJnN+xFW4zfVEkFdi+Naf7Ed3CaLjNlfJd1wwUph/VziaiXyvFlJBnvCvhIu/75hnux/p
nDEEhTHztRzGRHqfqx3hICX/baKzaixs2ztn5/rrmyMnqErO/Cax0G+2fGzrFhnUf0t9QhzCewZP
h6ntsn0+vCMGvmt5XcbUBBhIVHKhx+QJOUwGPfjtTqcBzS7NZDbfVNicYXHDvupZg9Pv8nPhWGDm
jasTJZr5j+JKzAB8mqUFFfY/5qlBXZHM+6CPGpEZT5VZFREtVzXziBG3aUxGc49wznrz1wzti+NO
+dkEVtf08cYUVonQbBg8f6LECWReu8wEOpmTNTo8aZ4qfQRd3ueknWxszUjQZYGshqMIyWAGUI3t
YwkxjzTx9JVdDhcMSg4cbiaxMSB9elZqIBdaw2HSiO5J6C5KD/JOkMnbs6/oBodmn0kVywRqGUw6
YQYwaotxnweCxIosRv3ENCKeHhhwU2S8wVzZmaGiW0jBvZcu8aI3s/D8JdXl7obS6m+XpbM1Sd0W
0jgpdCnm4Gir2Dm1yFagJfkClngi8wA/8tl7KtzuoONueVGiC618IAH4hVhxBRoIeYIulyVuoQLD
s7h6aelCjjRPWzhSlTVSyTOox3VlQpxrO7V2cs5E1uMP0foAJLe8VsK+yHb6esxcTCloLYDTDahQ
5txFmtliPK/ojzw5IeM89sGn8rJsi0VGgoYTOoN3Em2rM/YNHKFOlubsSPiYDQhyus/voxA0kKzw
FySBhe2hYgdQeePHwEb8rKigK5+MMDShldUh60HiDk6ecyEKfksAKjkFbNx93alYCb7lWg896yv4
Yqwd+1/aGtydLiM8QC5n7Sa3depoAlzj7Z7havDctRg3dd4UAgd37ilhVbzFFyXq6fJvmPihGygX
pHG6H7B1dZC457uJ3WRogbrMjAFhjuVPKsPlhxAeZZYOrod7ZaPU707Gamfqfo7ac6/Nggf0oCln
Jya2r7U2vKq80stIecTVP3BmRMXLq1pcZIaq7ffOYX02IGGQuTVHKtf19mgGnLYcJm5I33/tfxqI
9PorWRESDU3G0paQRQEmhpPJqqZHBNY35Tt7U+7jiDQLbu0A1Hhu8unecGfYFuGYmDP+kLFB8+pZ
PEaEj32JRtEqJO186KBSU3GL5bFht2H0HXcEpdUAxzszl8JpSR8DFjpxMO7Us6lIKewVVYsGx7pL
Mr7uYyUXYJQQ3+gAzzhFN0SzBcHPijbv+eD2EOjtPdglK4wQ6APvi6fPnyU7APcrlbUNcKG6fz8R
semL4kPh1U0+BTIjjDEX0tyrSwDjLGcJjb5ojKhAX4Js+vCNpP+KNU0wfqExgWhdtAs5cBzVEuGt
SfPXPgRZg+qcPIzqcbuu8cXE4Sft+mLrLBW80/MExpuNdyM9IISU3S+zSSq9yl+CmIrl7Qq9h/+G
vNoRxLEsgsCYpJmSiTMK4gjvFwOYSR2GkD1d8yzE0Mxmzh71ava6CmC6MNYuXUEXKYcKI5evmPee
eB1OPRue8D4uNJFSRF0cVVbZ38rGGFM+YfxOYh+QGfZu/q9i1ZYPfMr0cRN2y+08dScDAkepxerA
18aASYSfvtfsayYfagfMbA0xjSh4M7+UZFUrNIRsaKkQ6lQrpxzGLZjhg3zP2bFI4JGyenvza84b
0KWsPUXXnA5rpjXSvQMb4+aIlgJmBeMBigpzmNg9jUIXWhl/sxLdGzSORv2XyaluKHgohEwBSDP8
8jMuHlV8X7Kc4c9YMpNqrWFNW5nRj9S9CQBUSL0SvbABMXlYHYGtAQ0OJQGwN7WDpNxDquQETIRW
6qUA4vXZwYwoZe9RuVDfetiMP5ywNf4rBp4zzDgJV6UBHka4fJqteGpd7gwYOju6hY22Sw1DLrp4
WsSm/ZhBAMjPXpaD5PhmoTXRIkHxBa067FHzAlwGw41wyH1hzmF2nwv4y1iZnJ/c6EgOzSXN9Ryt
oC74AL4wWUcW9oJXEgnDFQt639H/Cl/IIEVDOlyZOBUmkBv5RwAzeIe9EfNe6Cg+7IK4M80Ak4TV
adSB2/ORIya0+VVS463cqO8umklSD6T157jNTI4J8DNXMoUxax9/svaKSQ/4qlfnIi1cfSNFskUP
oT4vKZ5lFPaujsFDnvV0xjFQhBFb9vHD6kSeLJItDzNt9JIbuJOOmfC/7ZTjgd9C2aoKSAen6a0Y
+NZLbo/dBPY+5s7GvsZVDCra+7kv7eGsmOdTy472+ZLggHXJfVQbSfb74VduO/qtgSg8XDVYQV/9
CfPqF2ThEKLDKVbgZUGedQjZRoiblXQLvhQAdNzXfWQZMIjoXoh5LQdz8Fm4Nv5/y5v3Vd5g0NO4
zILqAdOqufC+nsCFC9J+ilUJUg02shb1tKgBjCmxIU1/5fuHXojQug7ZdV1GH+ew4LqMrW+skaC3
8Ukx8APRhgcgpeNCn/my23XQRgXXLHzKA+35IoNsNVQ4cOHmleWXufs78quEbA+p5CfWXpXO8lAX
b60uNm6+Dg8ju69Wv3/ZHPmoOhLC7j1Oado0UBwW7UZPmYI6KvslFF3U2E5QtLuql99i2nfpny/l
23/NNSPtnbaZElYbXhJimMLU+nbNt/1WqXvE0kt6AWkNyFAl91yp4pcpO7d6QA4YMvuVpI7zot7H
EZJLjgWpH8zAsJn8EdX70/e0z1FTK5zJlStYE3Y1TzZxJLtsEkm/yjv4tldHLtOWRvMkmz7/LUkP
6Ykmu8xRxuf9VW8lIbTvHuwMRrXeMgowGMwlPO+80sHti5WHoP8KAb6SWa/p9Wke+c6yK5fjzo/M
KUYdilmsKUp3BEYepFuFMvhcEPREbVOuc5ZmXoVeC7jhEjT0cBeF1n4jyZ/uSVxfWuFdgLrooIBr
s7ceaE+6bxVZFKvnmsoD61CKAg/a9UZI771tOvwI4CNwKJURndWdoKaQT3+2XNYlEArnXzyjbqOZ
kI6cxRP5Q9uZosGdk3dh4TM57b+L6FemFmXEKw5UHXiLywQVOYehsW1eJkLymVpxZH1h7rRymAZv
APMcCJlJ1PSb9aydys0zoCmyUPxPqv3+BUkIXaQ+/kSPTgfNwyD8PTijqaVrugUgEqhTwqr/uyes
uZoG+EYmVaEwpuIlPn0SVvgfeuGniKsqFr0rDPi4E9dxBC3q6WnvyYgSZnJv4fpREhhipSPA/7Rf
Eki0JeXHPEw7tE7vN36VMCopU49JbLCnTXJtIiejpoUNgdhSz2/bK6FhePtlA8Th/ipGhfMfTEst
MPq8gAVbzv3O+0h6qlIUlpa/hVUBMbxy3TVlaTn/7c/0fTiTQoDa8hUHO6nXYdWFsfJ9sw+02Ay5
S2do8pEx9hdxGUVNzuTBOC00NE8gFya+A+3rOZ0jwtjOYxvPWUn+Gpcd/VIN87o8rkmvGjodPYHA
It9iH01H94bB3TRejMuoZlj30E2TpJqh7zj3kDypTGwK9c7xo8fhi8TCVMSpVUKF/LLiXQO2rA4K
B7DkQ1mHNz4xhUbxg47hENI4LFd+J2j7X/ETJ555oNFlS1imFosGv236tfOeUKSjX+ssFmSHSqP0
iWh63MfCqthfC2P3/LiayLsBSE95/+RIEdhmQjLiIVYOL64rQnX5+P98McBQdXB7buIC8DMtBWkO
nXXMuzXxd+bwDq1FQBmooM2tl19FCryOJzRb9eBlSoiM3OScR2m35J2R9FdCQLOr4FRvcdaDScSF
NHSn3LxBucQcxYjCU01ZHqZqTTlYait4nHT8Jbs9UgBgHxvn+7A4ZunaZZRjP4SLVg/cMBrlQTZC
j169EZEMToGV+RPPAy4PEM5BHLnX4vs4fNr8wGEjkm5QoygVYPdc/o/YQxX2e7VluHfUHHcspYv5
3hFF/oSTFLdTqw9m8vpnbfEzIii6+FSZ8wRV57JsEw8ZUoagusvbX4+8jxWAIx4RQJPBos+7nP3R
xO4OEVOQjaCBwQbSnIXwtJhdK8EYtwsEcRE5oW2UjA8+rIevsLNrHztkxA3rb8osSgo37Shhc45V
/BOwas6IFtxKb02FPRj+dw6DdZyzLVlrHE/QO6EcBB2vWKaRfeeJKsP5VyUDVk5TFtkkRmRkgjur
wGH0+jiRa3HUCUnnwJCZmIOho39CueS2IkQ8FkA6le3vH/3MCT0/ONOqJcWzZFoR9bRCrntCtTlj
Q9mAHhhaSKxlX32QnM9jBayA+Pj/KUI5EZKZr3Hy4Ow0pl21niJJza3zq1FL9lu+4ai6FCrPfVz3
LOxxR/enuVakqPMIzx2xAv1FefsU0BaLS+J6d2joPl0kiRf7aS2zNymcbzji//7AgOg4xsk/BPOx
KQx0/eNsgdbstEmLLL1umvFlcXX5hhbWQ7fhW4eU2syFvviKFFJ8DWe0byHdu/dqEfKtTFT4YIxa
9TP7LFZh5zcD3hvLBdYYv29wVaEsMJFHf9gXuII69zBKakbLF6zXw5UU5qAjusy40AO4hNnUF+1D
WknQ/dJiCObAQlbnUoO4YXXaxWARjtztR+cVItyw9EpXr+6PW30nLajmldL1Djao6ZGoM6KzmpbI
GTo28hxzAsHBKHUMbLdjS7mzfdwUBu3kDqC0MkB6mdQl5PRYpq1oP4Vklp/ERBlZEhBP5CQ/V1PH
7sJ+RbQhv0OrKqHhyXV6Peoi0CiPFPkNyPXuqrCGg17B3if7ioY9iNIFxzFW+T2lXYStEXFXd8hp
eAl38B8o7OcCUm9wSAmngwaU7D+j+IHK9rxLWuIJU7RbpLzENn8m3L3GHv5w8lsMYi2Nrn45Fodf
7fBxXRAfYF0tQdSRlmEmrrmgDBiGjw2iW4JoCB9jMId25oMOQgbJIWqsHO8p3DHjg7CdA79BhJhy
8GXSeZVMgU+3+TJ/e3ZorgHVw+wA3n8HekXv3eczXy8b8MM6NJYSmh5IyqwebIxPSiTed1Z8o0xB
+nKPmwkCWGBTpESytndfFsbphU/yT79giDbMWjtuflffs7bZ2Xi+BAvqTW5XjD1F3mlNu+SML4qa
k7uupmSv+u8Jhq7NsElBSVkP1E6f8Ii4MNfbmZNFV4URMDNixJqI0Td0ayAyvbGHNnpTsk7JgqJq
0qOOuxV2xAbOyDXOoE57xf1wAfDP1vMLhhY3IUwXBBoGZjvsD8Fs4+TdRMUe5VyTM2RRKtC30tOw
UXYurps1itLJ9mtILEVvsh1+FIw1ViaRnT6UULmgmqtdYDk87dwuVYtNLjXJrSYDfqhdBx7TKzX7
8mpRQSgro14X0E+q1+Qu0mAEugTSriAfnbxEffvbv0igfVb7hkkfU6uLSrzutVz+u5kWxDsGFPYL
uijnNRBukCM2CRdfRpoRZb74YS4bFXKmgB+LdBCS6q/ge77C/N/svZRT1dQJPHIhnB9Oc2b3Otq8
Ld8xgcCmC9Vj2y04jjWwaPa2xvyyDox03jIp+PrKBq3yEEo5Rtn/UggQuLxa51doeBfdJSChfLxL
7uksWO7qrh1/CnhQ+rObxNQBPWlHdzS85UM2ZcgCJciib1/FRRKLnLfszajW4N/XSzhFHJuRqpkN
DC2Psn4zU0RXxc04Jz+7BlspDvOq0gV5u6DQWMWEBCaaMHdcbz3cnr0gQ6HNQZwA1SLI0oGHrPsO
x2yhXuxr+SAEmt4WXFzhcA/tEy3r8dWmdelsx6wtE0uD0G65NFccgCT1XyofG29WamDKM12b6HYm
PQLucsfo4i1rn7Ys6K66gigH78BYVpEAjfLy6iSMYAiz6rdoQvhd61x72uGcG1sBh2gqaLRybQS0
Hg3ItetM25o7zZ0cdGCmuWvulTeEUvoAd6kEZMJjHMrU/b5KaRDvlkFkXTQVVubdErTnOQ+9J8uW
lSfDidvX51komNjKl6E66D/VyodFUC1O9bkNrlgWsruVuQD4tHUybEpS6vXqwnTYw6yqAAz9Zbdr
CveHd2ajbbDf7gOMTzTdSkrGJVI3gCw8I1Of/FJUJaJe+csug2f9eSHe/rnVsem8A8gI19WD6sgT
qMyDKEU4ltSKm6dakt2ioJ87dLOFzrE+M+CQGTeqkClgd7NrL3sO1yVxJegwRYLIPcO0HWL++UU0
Ct3soUy+Hnpw/5j/0WSx5d/5S0tM0Sy7cY5/7fWUZKDXJvaCVACbIoF5Bp5ueABdCKtBzOGLOpxl
ZcCBIZ8nXuBF8wrrHrrEPeKTH39swR8RAkzDfyjY4YvF5LHxisFBkylpf1EDpcx4mlKa+EmwQBTz
S4XWo80z3xd9sPh2Hfs3B4Od6oo/36MxGghRnfsM2ex2ztjLU97aZnCvm0xfqojKyi1vyL4qDKnw
il/iVS4ndyD9jLnl/JiyOu+gu2WFHOeobgZk+7z674XM9fSTu5spBzL1rR8OKqd+/DJmg83KLNQf
MiFkzPR1KAKg/yqFJR7EybDJxoRSbZ5cW8xdKfJxqP4nN7gi5fTTG0Tam9HVFd1pXq7jOT4THrdb
wPz6awIoHo9Icn1EQRarHOkELzdtLQPSUoPoJkNv/IGZK+ka2cXpqhXPYYAMl6s9N/IP8jg/4p7o
F2K+mMXs9EiBVqCer4wdijzSVAXEvhtksqb2fk+Nt08UbwRt9IVLFswhD+ocxEAJAU7jQrq09jzP
yaBoRKrhe1UD9e9fVSHSsbTZyL60Z43q+lUkYnbpYekFKgbgjjnPgzeo4nYWBMl2AysNMZkeIfPU
CJeh1895km9ppL1YJyoWMTnlMi+jIqPs4hz/D7EnjBL+tOyxbw5yKzVFpqAmaOdML+hqI5nzvKk8
11IHUtB6MUYN9ahSCYYJkeyHMJw24YSijiGPrZaIUGmYzKR7dMTlKXEpcliSSHXQ802+u/Isu1Fv
HY5qRJJjkc8Ag18FMkXTPBDfNkLJu42zB0UhhlFmQ3BYyEGp4gUDzrMNMUGnvICgUQKIS0A8b2HA
tG9QiRaig2YJCwTUfgXntwQIrrbQ3nR59z8yxXYdzG4BCF274QmxYs9Dj2IOVm5ZEw6FF45XDhGx
xP79JxsWMl/Q5WF8Ov3EQd1WNbn3T3q/jiTIEGA9bVbLyUpEIFWvaeRGfB870dSnAACH/NgJWoT0
p3Djltj5GRIO0svwDmj85LSR4mftA/+GEoQmILhRbUfnO0uJuuFDAbZVz0VhdoAV6eApkECEEY1B
tHLRQlGvB4QmoT8Z0tIkRLOOzgeStt04WFz3kETQwRl9lxLLn7X7SbFjTrIYOS8Oz8NR6OlAy2vf
JjsGgpP+MNgTg49a8YixLniXGVrLDuMPLWjh44UeDWiFkW4ZMt3+yGvtZTdc4OlnYQCXufXfv4O/
QYhWtie5mVqRVE3LXSypznPE9xDZlcwqwVcdJyqYcZSbs5tdnEc0ObBKj7FOudUeducOggl3gwX0
fU9WnfkOIufRzjmQOx4P3z3V4h+aj/wpOZulwFOoY+etBeoKAs6eFLWyJ8TPsXoKGha/4q8KWlKI
OddiYHnRN15LUinzNeQBcECt/GejEfUu7mpkh2Am+WXvF7MlI5NZ9QMJfIisaBBMaNKqr0yvKpuK
ZsE8fAZ1GiTjqI5vRtMDNY1Z8o/AUXiAf9JM4S1x6G74MRbalu+k25ATZxpKTxT88U0PwCdSFXRF
U2fS15BJqV+Zv7Yo9XBWXuqMYQhY1dHpXh1cnn53XskUNIh7buGE6012TisJx06K1BmyVz8i4jkP
qp+p6iFIJKDtqBQPA9zjPWYoSXaHqwDt4iCRHLUv+iMgJAGS8nQQueLO+LTlPMJM1migSjGFuK9/
kh2E+xn4Q9E16zJgmhnlHMk86bz6jpKLGQ5Um7D/rtyfVLPlOGYXVhZ5Kex9466FOVqNpOY4LtP5
7x7sZQW9ti/mGV7/N8O4dvm2VOZvIgocCq123ezsr7OBzpTZldi+NtxVT0dOXZVdSWQS7KuciU+g
GgU+VqAeBpJlchR3KNEKbCdvD4A8vlDDOCYs9bS4UpDRmOHhHd35D7ftUTeKF12ONFKtoq4tMFQj
0O2uTHa3YRfDRKCoflPn0GekpX55GdKoeWPu2EDhlBgk6AALc2OmXXhXOVp2TKb18BBFhEaDsBCk
nDD4T91YIOudKdNcJ+Jd9vg05y/ZNGBhX4LPlX6FMhGQxwot6eFy8fylp4+LWskWhVk1RETPKZta
PjgWBvR2bZ7XIPk6KKDdyzIk4hm4Z6lkif6IOQGhb4BIkuQCUD/IBo01pydkGAX4WOdwiuG8Q0Ey
PWVwG/8oQjI4hiPh52xsBup5SP2gDRlBV5LAeg1vTulW7RyQYb5cWxpq7lsWNdPwDs90umla0Ln6
L60HCnFpOVl48aPOEMR20wvzNehBjMEzxLzofutkmLo1bvbuDCxttzvszdB0CNEJHZPEzdQvKHB1
mrxa4+WyYLIRg8tLxBmUJQq3voPb5IPbt+MSaNOBOfcGdf+jrBe584qV9QPNFBjG7EBdf1WcYxvo
mwScwpA4FhBTDuc6UdRuCX8tcgdIIyqICfqKwhZII43tBK/xNbu4RHFukNPatBtylZZJ09LxT3nF
w23oCWvbA/eMs3yECuO5CpM7Lpn/OFINpcZWUjZMWk0PlvGUOMFzQL46ZgijBosjjpNwZvjhlfre
WRzuZNsBgpnrOKTankuvNyhJ3nGDY9KujV/6vMSx4l80WR14cCGIIkEbt8Rx6sWEWWaTm1D0puJP
opaHex+aPtHLmI2rTen/ELMbCM/nY1ukWp3JqJPCj+sU3mPTHU1AEXEkqOEfvRHCLZxR3UXkcrH1
e0T91APYew/WK4DBF+X+FHxDUijebrxQucuyfgrvnBAoNECComcTV3h7GLAQW94OuHefZz91sPBs
KruayLQtJF+RXwvFZPPmLusU16yJwob+5ks4/OtwRdbyWdM9f0bvJ/RfVTA/KMTpgGFOOAOhXK2b
C+mI5jhAZaIidBybmOLDMSEbYKI938BhI+8S2RJZ2z9RSwvIYWi3NCaxndIx2Js73TS4L4ITRscy
7Es8StAo16IgRjJcKXZKjz74VjlcpgVWCge5PzD9IUVprV20wyp8SMf1gIQOdZC7qhpZLPj3QbAL
HlIu3A1UN7m3uXJZ7/edyx44Wx+7+VtdhVA56x3rgAJpt2SMOD7mxDr+PU5Tfdbiwfw2UlLXBAfg
Pjr9gXsaBNqlQcNDdvWPdnIC4vTfJ73ptEp3YQWcc4dJ9bHRQ78b3nZzGKDMc6bUm+3sghoi5gz0
kV9HsgzZxCJ+cGFk7ZDEwx2Ph704t5ve3gO7Wwtje+WvKcPQUOY9YOR/bhU3rJFefX/DeLEX1DKf
+dANFIgFWbfT9PTJ95tNdHAogZ+awP9qfuvEoUJTxGd1FjMnzNnIHUW7ZjlO4TNSDQsPJj0nClX2
Fl1ayiT3kXxsvyUlpphMOdbuYFVuY/gpC2dSVhtuviombNWXuFJz6RUqu034hxwJXzf5OeBIuWi+
y3IN2g7LDos/Ca0e+qVt0h64tjoAu1/PO3G63nhY8tN63i2oiBt+XZ3YvlnQYXcmjM2IGL7Kuxr2
158tj9pk5E96YE9csF+UN+kWDvMT2IBFVThO90Z1arKvLt3KPsLxkLkmheiEEHAozHeK2cs+TUI2
9t4s+Goj1BEEeQPGW+tKPdqmpafqmgRNY9+4p3+ANlTMcm3THMSflH1xuxXOHFYgSUWO2QdNYK/x
TtbYy27Zg0sdtOofQXR8sP1voswOapAkhgSaK+kO9CVV3/yFVVpmsGAfs8Ukz6xicA66bL/94F8T
XEtJA44X+jd/Y9svS+o0NdNjISCaSSJmRkVRBTaNnbzI2ZLXVfnT8dZfyjulSKOTN4K6d6PzYeFw
pY1bWwvnGDlWV6wgoVQvqA1DrNnQby6Eccd3mpIXvMlcKOhMKYroef8Niwh5yZo9uHMgCmyOmC3Q
DlHJbeLOV/9in18B/2CT19zjE0GHEZmN8HA6U5mFxKYcpC90OEzgiZ5FgLIdAUHSDxrRr9CMXGTK
XrzId2QX+02JyAYy5UPl9+IzQhv+GrR7uiSwk/RzXUQ2vPtiebCcV0FAKGgGcULm1Uuc9k8v/LRC
6udfxtgr+lvau4043Y/qP8SNctTDCXHoXvy3JhoJ6W+R/AqNG43/d5SBjp7O9IYoIoKAd2qTxlwL
nRqdbxaFp0HTSenX++Bt8yXJwTUjBnUMslDSX6Kh2rqrJHb+ax8qFsCeZKaXD9J1vpAkbx1Oaw0k
TNKYXEGvoGa2FRlDPOKpqABVBV+PQ4dEKGXpocDGx7Zok590nmLc1Cl9t4dRzbx5HwA8unvJlCPG
GLK92ELEXXWqQSllpyitcYnE7ftEm7gHzEjwi2paMaxCtSpofqRCjcRr4YN+yf0aMBNLHLwAVAS2
rSJu4WwiOB0lUpyyG/h+lUVx5ESLCsTq9oYu/rU6nBoJMNiiwVPpl3tOL6S6Tu5m5qNf1oKdj6At
Y4ksXmijex32OQSmXSnCF0Ei+zyIFVi6iEujpWZf0PPVT6wSNs4Dh8GY7QM4MmdCS6+Ol6Oyw/Bo
phzLXQKx2aAP4RppclohG9+8xiSIrtsFhcnP5Of6WV5huxtVLkE9nYxXCUkTb/bxenOzQfKD8b1g
6jWQcE2hywXEnPPxip1mqW6PC8Ax1Tao7jHoOoN3oBujRMVxDa45QibX6UlEtvGr1+y3LFHfUByY
8IVFtn58KbFHLWxiIEAgzqO538S8VQCdRe1D5mOrLLFLx5xpCJABK+CAdTmKdy6gL1RKUupht7tH
sQwQACy3itf42blqGbDWZ9jgd/mSKJNOElwQvB+DXJswScDashGFXLIi2APs8Edh33uD8/EMuc8o
Ydv0D9kS/h9XqSCBHD422QDn2Y+rdBF9kGxcKwnBEQxgGseTzlG30Se7pX05rkQG1o1nvQQGuY6l
XCqJemcUtZwdHN4OXbtsjHUSlzBuAjgg3tyZ78tqU1QlbHbcgwf4qrkXl6D8wcyeEeNw9uKnoMvr
3136fkLM7Wky+lR/NPxWi6xYyy3AIRqRIg6wjw4+V8EoS5oKpNB4Gxxp7XWHPy78clrj/uZYroYF
6bDfCFWcZP3rFS8POPXv97WSv4vAf1ymg3YiCryh9KDzd565jZ4eNv31XSvH+QuFQPKXlD4qAuAh
jxmnLPJL/zbMXRCANkQwSecMr5WWJfP2LYbYMdZLavcHC5aflAr9jezXcQIeZQJEaJDQJPN55o0g
5QE/8QwJ2+uyNeUBGceqDSs5EqfJI3Ky255rpHbstIIWlP5FyLX/3Uc5sUrxIkJV0mVxPiS5qa7f
+xpBzxbhjFICmFFxmJdwtOhl7+8RW3iXelEQNiB2HQMn+A2LKrqJkI9nDkIyF6C4KE1Tgl1Ico+u
TJ3RTYC1T3to/AoCE7z6h28mMdggXMoT/ksZFTnCRT1FWd0Ia9FsgrtD7YihxJ9h7MMpLjSY5Eoo
XcLepPTqoguBzdE01CwUbb6kQSz02OKWeDguLRJRsCr3WvRFpaQYeQwLcxoCgdu/rE+arN6j3R8c
tfIiv2WpBdbS1dJIRgIg6AhYkvIB4bUfBAPjM2ocQ2Q5cjl1BOtZ9i2DIDehljdXIkOTJDK26VXz
p5Xv5jxPM06o5tAnUkD3vyHEGW0WBaDUVAgEHJkhLG7TOOfxYcIIzm+OjDCifWmcK/URnZYse/kR
uBGoDa+7FMqOzOyMwJB03QXbh1AZ4HmLF3BC2APcp6cQDVYReh9D7CyCgMCsa6wx3f31wN8uZA1F
CuXjFLcFYH7lDheHUMkQb5ef6f8NCxp2i/j72eCi/acJmLZ3McPK5bb6NpyckXnqEMeqvdmbpVXe
IQ3WYTSb0BI0fsxq9IUfBJIiFjZGxWxpLAQYSovG7n1z5nz5gIuyrfzHBC2d6O2nLEaT1hhzvHzj
bcDr3H/rC+1OwULQNHDi0qcokbPGJbhPU//eJhhDH3+Dt8G7LiINrwfRq0qSrGT3a2Q/yBtRTTw+
jfRD2FYH51sRelFGYPJoiC6v+vw9CV3TObVZ75Id60sT1pnrds6DEjEB9EK/IGTs0+gaEjSIyrja
tnoFfFylj/yc+XsXSvgnjYzPDCRXsKTWOqeZKXVT6pPAQmTE3iivYnv6pqG03LxkqD2yCbREQxWo
kIL3EMAllhk7XQBQ526LGV08zVKr8HOr3r7i1bvaYRsNXojm7Aet1LG15sIkPKQP01pk6zx+9oiE
IyUxTXIid5qpNft+fUAXCO4YOozQFoMHS2oCNbTP/J30j1ZACZ7dzTCb8EmT7eEL0MvzDoE2sUuE
X71b0ZBHUxGMll0fvSXUCk27loc3N0jn8WhI3B0thsRHguhXn4ASl0rvmcDDBiW1uLAYPntkvLD1
R40iCaTkA9X0sAGJquxcveM5ds4hlTSS20kqdjSlUXhem4NTU7PZP6p6KSNBHESeJ1b2ZRHlaqiY
kBrqowar6snaoWw0yFKKgVXwdFq/Scm8+YK18wvbn8V5pIdp/isQXgraZTW9cqIjpEBLqKRe86zR
wVEVfxZVkHpL8aL5f7mjydVHs04JIpOEH/MV/y4yKzsb1uJxQG2N5819M0CDh1kUsZYQtfb4XLtW
oG7nKrqpQQ20+jjggsnofpJ8VzvhHxBV+o/xGw+hUmbnB+7h0Y79kbr56Q6fZsRkuHFzjW351FzN
gMzV7MUmKsf3K2+vTd9YlhwelMCJB4oDZ//A2V7qryTpKap45zzuvPGkTAnM04tjtaQp2ZWw9Znc
p7XVqdCWFURWXxusNDEJF0jkLVDWJAIz1TvWumvBwSDfseP25a4yOx7b9ddHu2wrBjiIkpfHzdJJ
xncPENGYqvS2V/lcYIxb+9uQ3allwXzE6O27P7e9nZa0v8mVGPTsc5GjAFroEO5NT8rG7846dEbM
NGj6Np9K0Ed0ITYOnk+w199f1cQ9L0x1YAfQrPyYV17enDT8twOufh1ZARX3GWNjKVYmur4WVV81
aZWWWQDYifbYiPdCZX2ZSd78TFjpeNjjPrHfx2PxP15PfqaLkiDtf9y2K9kKyepBoKmeonsasW9H
W4uaR2DnlQYvFjKHp8gynnC9lVpGS916UG3/MCsNmc5/8rq0VZtO5BJpygVRfzoGyAyEQmGHiT98
e9WCK8L2MEuH/FqS1w9q4IP02Z9TRPJ18QzyLOkoIL8YSrMFjywHK4ytss1F6MQESNYfAsnC6FO3
Lpu223JRvNYA2KB3QmSzeIrnovXV+L2qTV7K3/WIq8kKEp6ncVUzh4jznqKSbAJ+CUJ31EptYngk
pw34RvJKPXwe+rSRIZ6Ex6aF7sbivQ+fTlbAzm1rXd4gzUt7buU513XAjBvJFxu4R/RexNd9d9me
JuV7Xp6j1Jb+6Uv8H33g9K/Kx8Xm4JSIgCGmRJqHW87JikzZD2/vD4SSkbjp7x53YavAmK0nNwlQ
Ro5uKwMVzei3zV2rCIaWGW8+Mg7W9lgzjmalOQuXHjgV+OlqheZ6KugQS7DK9vpE63zLB9F6csNa
DgoxWXEVi245OkAQcR+2m2trAw9Qy45G0hjI9Gz82YGPGM2CfXzK46CvGnMW4ifgS4BQu4Cl3a2B
v+IHGsMxb31WvI7l/CIK1R3Ko9zMe5OkRVaFc7jatQ6zoijqTWlJHTcEaC65N3ahpQFXy7PwADQ4
LeDWGSnn5BPBtgEZ4Dw6dF7HadLZ+DRJgZEC75slnMRM1ZnzOA9KT4gq8JBmYC7UACC6kn87ji9u
lToML8R2AOoXIGAENLZVyqhZkT8RJxLFcTVhgexHX2KJ/ThKOP1y8RSTyWALosb94D4F1atAgwGG
hqm7mGSKX4JGP6WXzx7481RCZYdDipp4Z/lL5NhTQpCmWB7OLvZCyfDIR88P99P6kmXRpJSqc7Ol
nHJS8etuZdI6zSTWsIyNCD3zxsVJVzHmqhxKd0bnfZUpCretnK7ppd5QNnAYjqfW0mo3gXBy1sXB
28Kw1pYhv1lsh4IdUYxa8rrsJiamEBkYYmBsDfZi6sJkoQebgExKI6e+8k1x0KN/+1iKYXPoiYfu
IJlVIFGXfKt/sC/QA2IrPYi0uBbCgetxD+ELvr6EO6pA4+R6OH4oLlYl74yhbQDPv3KRoVfFrlUb
LA8WFC/CfoEWApCIdmB8NQtX68LQ7NCjqcXEtb0ENXD6AgtXZRQDQeZXsDCjCuTx+6qTl63oCN3X
VAJYSR45MFe6rmBBPtaC/FZT0qU/EUMg4PQ9LIeXBszT5YY1iYkEfMKur6T41Dq67HrsR/b92gHc
qBg8CGA1JEELzln6hBBPeCGdiEoj3MAALcL7XQuWbUBAzbjHUlu3Y5BcC0QhP7hlRrzUwcY8UCms
vMD/l38lWzEZnS5n/PnTNoJgoyc41piq7ovpY7CSf+STaemxAGpOTPcdUlilvGdOIvxscSh2tKAA
aesh9HhnN3tBjNEpw2eMFVC7EPIWC+tDrli/uLne04LuTEGBC7ef6/dw60a6KNy9A2zwDK1kyN9Q
A6OYnXwHpnuTJNTJt9e65D0V3sRuJNudupn0KhwrFtJVsQp6QS9fJWysu3Fkib4876i7c65cBqNh
aNWFrlaTpLztbH2FDuqrcVXMowpkfnB5LKcXlzIrcdYMd7p/k6BelkYet8jIIZhyP4fOxSJhj3CH
FOMXH15vWfhep+HpDm4n/4eMhKAqXMqoF4q31vkI3gFV+7017PtAtdahd0m+MYZjARbvxu1VXdkU
jdQlOQ+jbkE/XUJ7FeS0aGdIpMpnB54yiiS6Fq1UV29JwLZBnZillyqb1+DzGubHFg3VGnQOTRk4
PBJK8m6PXHOclh0C8jPuFn33IFu8aZQhltskrZKl3ihKAi21Y742hQhSo9E7gzg+hYUwlUOAUpQz
Ky9SyUIqXJS2t/kKUSiKh9Kpxrpnnqjxz4U3EGYUCI8Y7PYAcJyDt8T/TqM3ROO1fVnD/EmlZ9mY
yaoNjftIxACMD8rGMnGIhUbQlv2JoWxm7ppM70vCrIdOFV7lj0+PVU1JPPNRgVgQBtt7RAd/hJkg
eIGK7f0YqqnFBQZFKBoYMo17e5uZtg87EHkzPEu6ERYWevhoA/PY3KdIrTS2JshNKo+9+Eep27jd
7TQ3E7ePwjwzKtZ3COcBs8NS0r5nu4I2bVGM16DTQnfBdX6FoxlTiGWPWv0+o3uw3fUXsRLO+0Uk
AT/4eQGTGxkTo3lq3i9yX8GUdC3egscZztB5YBArNu1p6Pz7XK+im8AuO9UEF05QYBMxPB8ta7DH
swPtwVB1SMNGSaIREvSN2O+3XBf8UpKea06hg4kZpPqT9r1/C86QHNz7x3JkMJiHiZGUtF6HDE7i
GwBK6YZtOhAyX00+ozS6Imu+1FviQAVGUyFb5dqYJw5J1Wk+CYa5u8DSHqutY+dHdd9sVBLZJlOl
FirHAaG5qZHi6wFO0qecLADyPtziRblk9d/qltyg7eZs5WuT7/VFKEDZCG42ChrJ84IS8JfCKen/
pmANJ4szaDBDEv12RInuXhSIjpUL/vdSINfH/E/JwLq2dD338WleFuIIE82BsWw4ZQ+j9mMgPU78
ObKGBY0C15SWJtCfDtE4QGnNx1V8/6YrqZeXf/BIv9INwv1D6nnZy4i0aNCLQByBvYS+GONASnhy
0/UpRsJJcIn2k/gkXd7avasKz56VZIlNANKHe9wIOYgpa5xTum6QWtO8sk9m1EjpoJeLnXRpqZeh
HI5COFpJplK2zs1gUUHDceIWt4TiiXcJaLW4e/Xghuy00VGXS/5v4pHJ2yvPiiazj20tn9VhkC9z
kfxCWuSNXCSRpLPtaf4GCU2EgeZzOEnrOlj0M+VIiP+sgK2Iez2H2BEn07Pnm0RIl0xRIgXlAXo6
Zk4Jd4+CAYt/aLjj990tcgeMeAoQZBQ49edZjrT1ZZVgDJ3JB5ikuvO0DXwdrTCPfkzSMNFyLCBN
D+W9Bymyxg7bttHinPXfwUSVMSBS01QGHx0x7p3VIru/aKmPCSfCu6POi7wNpAyVwKiZDdh60kn7
fE6gS7iESwfnJTKX9Ivq08tTyBv8lTyA4cSA8WKtYBNnx/ut2dmI9iYZfVMC6kvy3cMd+e7uVHte
T0Z6Ie8jasqfOnRGymhVKtdI8kFJ2SxsVz30B66It2WyhwAxoYeIlXh/24CUWO7VfyjYvxN7/URS
FZfYPQzWsOj5cHbmOmfqRzDMSblPXpxjwTdV+6/3i6WQlHAXwCixEo60zQx8jKKLrPiVuJ0xmCcC
WStOKwLys782X/vKYvUW0mMDlncMqr8PaLPj98gZic08H2f8Ax5tCR8W/zPc/W41ly4hlgrhTnfd
Hnoq+dXGt6YApEcd4mKgRlpucvwLm5z1S0vAsC/hc5GeATZsUkidHepy28JGETZJzQYYa5KIqFiT
BW6HJIH5aKFcN0nvxYekCNG5v1jAnYdeBI5SFBiC7Cxy5Wr8h+O1blKBFtmJamwPH9FROTOq489V
s6RW/NWGxfIrgUd87NGiwL/CziOgPPU2NKX7tDee+SvEpNd4rhR+N2mHsIP+Q3Q9t4Uhs0hL9Mmz
eRnFDhY+RwQ3QURjS7YrikaimQkyEhLujrzsxd9dhZJoIBtTrHKYJcGkGUR8y8fNRKiMXDtgSOUy
/YEiVNfNoPbyGLcl4yoM+awuSQMD9ZCXKmGmla+2YiUjSf1s4fwEaJfu/dWCkVMRxZxYi2hxlwp4
+Md3uwD2P5G0FJutv648HAopDHMlguOoptUvywOi8u4agk4ZI/dEEsznnPdnVdIHXxq7Gemaz1+s
VukEbGvoig2/E8nr4JxuBF7yX7DkENvRTiqXsixqoDWUKT8R9bVjNCM4QHXz3wZlbCeA+qSA9Kyt
C7P3H/YDdcv+I7titobA2NF1P5tab7qg+nnpinulkZlt+UVc+cCf8cEWWtihiY4TK++XJZDbUv72
cBnlJe9ootu5b/wL6auzyKwotnSYrjHkCQD4pu3Ms0hd67Lvgx5daBX1Mq1pjJklfT4pUdkJ04Gk
A6UDszmaVOpkKUrxOBF14xIOuSB8d1dCaZuFx6+0Jjr+KoalWztFVPRbIK+TMI6YgJEXynTyxxB1
1dxyTJ/YbVMFxo1ktnG0gHbSncczfK8/bvpXkpScp8QU2dmcXK/dehqKPhBuUq9kJPAy95opezyg
MKQD4Prz2Sq5Jx/hz2gH57VndsPe96ZKW3B66kz254cTFkiFxJHCjEqR6K7DXiFFynIZFQvGqJdp
ompCAi9GzbACHMEBAqYcBgMNa9lKecdGFMpDjV4ObL4Ww6xKHeD0wGOyXdzepTf5prWHC0kIzrb1
WYA637xLalbr8WEcp3OVx9wuqvQ2D0KB/FJCAuBcKqEnff2ZYdHLIPRR3K8ZB8sN1rv5Ec4CrJW9
PPSZI24HcDgUNnyGimYsnDVhT27CIonGT5nmlUh8/OCAWF/Yvz6aQnc7dbLcygoNj3uxNPNErWfC
wxZK/I6S9xyJufZBuVScqL8YTPuT1nhs9AHpig55H6VC4055bS7i0P7djTPEkkYPEX0cnROd8ITv
e98GnNBciSskNR44BJqLm1PFkANk17XZv+QovrEhGBMUhEUVkh3//4giHMy4KYRtLHkjh3YjdpXe
LCNbaQvPAwYy2KCGqkZdGu1wJBGHfd3MVEfRKvq3LCMLeLhskCdM2ry16HBDnZEBUrOvVs5u1MLj
cNiNfLMcecDLOtUVgWha9UgZt2OX7fAqA+rY+aqC6/C9rZtjzZuHeLaB4Pk9zU3r/tf015K02dsi
oaFZ9xDa4AJoIk+mfOpI1pHOJys5o2piJRZvxW44ETWUMGd2azO9h8uAPaB+rGJkLLbgjBsW0rf3
4S6H6QdRSEm+y4W0q2ycguE6tsQ79sqPrK8RYRct5s/kN3GSdeg1YmPS9JdmF6hpbr5yik0zWjja
rizzyCPGdQOi+HWem7N5aH4zyzJD40XH1xe8HVSLWnXrWiMhZ32UA+z07wi40a0mFhzgV+/t31c/
QTgvU+HoYrQqPcF+HGJ1CRK0CRWrcm1Gm6sekNUQYizJ5H1CNjyykM4HfvpMFTqwYE6eBhsu3sGm
Qf0wsGiP1eZNPZBJ1cELx7LTobag4NKa7fkUDY/LXzMy8QUe/9/aTv4kxgSEokB4XT47G5T3TmOm
L0Z2/n28DiQKDrzw1jXVhD6/XJQH6vOo162n5NDOnp1Woys2eoWI3tF4LawNeyIgXqpjPWUWXtOP
xoKo2uc202+0rmdTYN/FFDxv1pA6SgkcI7UWojtFOtID8KEppv/qWm+5fJ2oUd8v8c8RFHeIQeYS
62wafA0ugoZCn6ORy+dcpQH5WjtXz5krTDSqtR34CHhZF1rdaINs5pYMkJGDDkRq9iMdm8EMz/Zt
/K68j0fNBvarXjKzi4MARfwBmV6eT9SFH167Qy8rM8tJdsSu8HtDKObdlCNSx8586hbclF+Pjr2D
+ur5YiIxJDyYHjkmg3v+kIxpLdN/8XArrV0RHxttPfR+tXV/cNJLEs7dFrdx1oIIhXnYvONrLhus
IDNUwb9NYvv9vp2gTC7OqHgCtpLA3Hfo4++RUzsPn9RoP4Atjr+6UhLa0A+79lkHqpSd3f6a7UNm
1h+2u0t+GAvCqINjIX9uNa0k35y61wo3kDz/9NqYihOXxiC0u3Ag1ehRQ5cgfgP3mNSN9opiSVbH
Y7quxUL31mx8JsLYu37C1E4EK03qEC7Jgf+aXvSxIhVwptkYaCLSMub4u7CwcqkbjsFustkFjICY
h3bxk1f+ysaknzlK5o+OFASdrH8pXJegUEwgZWGglnQavaR+6x13QAYtWMTgDIiaA4R1v3nNZa5+
OdcXSBsSo3bIq9d2C9ncX/f2aQwtF/v/x/ICoSC5y4RRkzJ8WZpzAwKt+Bosqcx0cXw1Y/n1ro64
965q2L7kg9wXlWGcM2/iVrx2YzDLuaDWJB8pCfj/rwPyWGBoyvg4OYon+J2Qp2a+RhxC4YGmMf98
sfbNcxfOPMCiqWhMkYzcpVYPtkmFN+M0mxne9FII7jElTzNF1UtGmPXNQZ6YmhMz257hunx27XfL
vEey5vgpDrc83QOAvyO6Xtkq3g9OvXlSHigIpHEZClVx2oyYK31Lehprg3L41yEHZoYo1Y9ZgASY
vT2Ggr7gyDIgrKMHAmr+tojXcTVbBRr9gkl6pO333ZEyRF3HKE7JQHcoifrgyWlJyhu+UYVUlpI/
CmetcuFAdB9iZXiZiwZWa7ke9KCqYRfz5ZQ5wK3GwWbzN9L2Xi1Df5XjdQY16c9kVY1nGsQ1Z4KN
7Gd4+2Fvp7tuTGbAGBGuoggnmao8PTeh1IMbYLcEiFiTimmkKTuKRUvrgLgOJixM6grBHNHrpi1/
pBQBAQszg5hRR2cbjG+1+y+W8feyRai6J8oWqdttoSDIaTixMI+/VY3qEGJYHLlTKHwY74fv0x+S
S7MOfe+P3/D29c8Rc3tNrnqXEkYPDIuPzj5aCsoIglc19l+wbTXDQOH1UYZ7mV2zlBO7JZ0S7wM/
CFtlAnlXGVRaXHv5GEvCHsglFP0nDLFgmZHtHp47jziVmHCpvnYBPYYt3hXoTFhcUrnEGgPmsLyy
LwcIpQ4UZVLYcWzPKiNuEfHMK0kHC1NlkYJrXwfyZVCkeFWTayfEiEBlMQl1O9N8VIGh9YxhNuyt
PowsvpSZ1uNYc/FwdH2R+bkjIWOEuZtKWFBtpWvy7cOAKK3v2bk+TWOr9mgJQ2uqaVqqNeUYQAh8
EqmAYeUCtPcBpGSUeUT+fL9F/IQMOiw+QuT31ggahY84N1zGMFNJKKDd1BWiUQRLNZ+pd4bk05jV
SYjPm/JafqZug/rAB0BCYmda9OzjHWud0HpBd/YVdQshlrWc+CUUOvRmFzWXEAfyV67d449YzGDJ
AgDHL7YVY3RY2IpOJIjPrJ//UvvLGV26cA4XK61w0pEPkq4UX8wyOVtBHYuYGVf+aCmx05k5huZk
iYicW4u+fIpegSGtX5bm2YGt3QQMAtXmFNUa5LMZGOe9w3u9d9wysO2cEfOccZX/kfffbH5dgvri
BnVdOuhgZSliW6uWI+LZdMex+rXJYno9s98EVMOgKDKWR0SQ7SYW0LrL727RTbzPs2xw0XVpTvQP
iFupAEx9NP0vnDUaFl/r9Fs4+PIJ1i93Ts3s9fEr82sFg4birJROmGzxLzaKJprY2c/N6/I0OUoL
KuGErUAjwiViLokJCzaEGuZsnNDO8hMAVgwyvxii/kyHzS9frEmhAoYQkua6nuuyBAxtbUCyFUf/
FIphjO6mYicegE9nKrHKKmBeGzsMfT2UmrHgWI7/MtDj+A+MkFYDgyfdRiG98DxizM6LU1uwvkta
McHJklU8gO0+i4al0uHy6kEmiNJGNna1pjgvtVGDTWPCLtsvA+PZnGAk8ETonXvgfrXsv3ChbeFw
HzKr97EFp+JuD0Rvb5Zn/iYgWR+Y1LOs2CXoxOAOQBKoJZ1RHwLO+e6WJPyKIqe3JMbDLdoxccW8
EKfu1zDhuHg1JUBcL4LunaSGtqhRnTvDMp97NfQXxqM1pW0JUMje4DV8UWZV1oB8CzHxWRD66sdP
l+PNtxtmx/cgzpwGsIg+p2ZtjJiwtS7Jlbb7MGMmUkSMETzuTrp3u18WkBtYrWA+14Fw+2CE1E3v
j94jWLniVYqcmt+uL5UTclTNGTbzdxdqDpTo84B54AymnFkfC0KzlvVrxl+HCmaZJ4bgce0Acbxm
+1FpmKoX5/8xjwzNnVyZrS+dUgjMkz4ITJtBZfDmNZIUyRtk6MeJWHJiTmFrXNZftPNREmQ3vEFR
Ekp3emhzc6Gh0b8R1KTLRWrbsSxBl2E0HlFLWKA2PchRC/5rFK4B1LAuXFjPyDC9cEr2Oh3ZpZXQ
0sEIEVnOdASdLxzde0FvK3uXOpIHNXlifNGJFLoxBDaYge3eFxmmnYlz7e6m/vwdmnKqfGscVNPc
5RZxt4D3kqgmZ3aEYtVhlpfKG/DA7RLhER//EW+6t6NfLLma8I0n4YJu4SqdjEzcXO+tdLLM3jlx
2XG411Mfr7u2X9sU3V6UDUXjYIXFIDahfDrJrwt76wPqr9SGq08DH2lIRi3pbCiZnM2y7uArnPfZ
6I3DQrBzW1glyaUEn29C57Z79mV37Adt5D0YNdTpON7o9yZZwbG9DRAPRJgYJDHH08B1lLQUJON9
T+SqcAecGGQA80MGIlNsvvdJlqZjRYHPj+YL98G3m3j65fdS3CFCwE13c5sBimiqQGOEXtlX4b8O
JZMwAPvfQzMGbBgb2x4udlQx7ZkAwCX3ZxvAP2xzN+O8CB2EQUbtLeWfRwqiuW0poQvgL04gmqQX
dFfJhyiZShbjldaZ81y2RLef82j0k+975b9mOhWtQOv0lMUH70xXaVI/x/kXB8E8uHM2/VgDr/VU
Ev/AyfFl8zT7Ob1UbTaukSL0IlT3eJw0rCqoq06Q99eW0PLjF58XHk6o9N2vhtRMNYqVpQtAjJLb
pf5+ZQ3w8tWhrCyHW3DUveDjpwY9imPqrDmB567Tgnstznb1kaJM4/JlI2WPh3o7U/AH8eIZqcNN
yhMU+QyHf/GNJIsFDroUaGQtO7KsmnqcN1htetpcRlKz+DaxEyyRDs0qGKJEA8zCHq3Yr4GQqK5A
M1I+IIW9fM+C/5dOlnTXKFuCXkGGULM81dMrkiZIQ+gJO/lqEALzU9EzokZsLD6tXtBZNCVrpTnv
TR9Z1hgZ+ZDrx7acIo1JPWUZT0sDqqwOrgDqHdxDT3d61S4E2G7PH8lHJLcV++rDnk12BtOtdvmS
MfeeKVtReENQrB61J9r3+xUQAfcJq0C9Cy55+iXMpyDLrUi4DdcRMcqSB4Zmy2OiyrKz1W2B++CV
1YjETbB7z4wyuIsWQ+2Cj7wFRXOwIox9FIfO1gdHaVZvyWxb2nqwZZ3Wtop7OImjBiimVDjgNXnH
8P07ZhAMxHhRcDbx/8b0RW8jZjIAQ7nnwpVvFYP2LA9im9w+n3qVFe3ciUyFCTn3fmL5ZZaRZ0Fu
zuT0IJArioS2GiSWiMv6br6Ir9M0XPWagS21g6cYyEFX1v5/QIzmDgrCSpG8psVgMyUV2ERiLPdU
p2Q2ErZYNNEdcaXCobKZT77RqPl39q+8A9kt2mMeP1Xm+/HST/8SvG3+0wP1RmTSzxYN6D99fIhs
O/5p4KZDsZOGc4drgTlOMh4a7x/5UcMFBAKJhUQXLr47Tqh15PWCWKuW5jZ8o5uzBvlcFQpHUXXO
6A9sMFQz8+rweed+u4pBXM2Oc9sPBs3nlPR4ejkUjHimrgG3Ry6x6EwhV8N1bU9jR7vL74EYSO7A
cBaRZQwzxuV8hRz4dWCl1BC/O28f3+k7ePERTzaD27kLYsZmW6fY7jjs+U3RoO4YAT5jECDZwcZl
baKT03N6isQfu+Z6//U+wRYGm2q381uy0z4jjCLdJCLbEQmcPPvcWmRxfFHnns94HS2k4HR5gNny
adR5C+rIP8A8d7RaOxp+1VBj0rey9Euj4vNRof1l3qsJJBUHfMNtil02U9/NJfbS/gn3H0tInmoa
r7Wl8iPQSrcw3lJtx2Rv5b7/V9wrKYO02LB2i95yUhEd5izRg4vJY026jdgOZjSgCntDTig6B+Gs
bAaZzK5H/hivuTl9TYH2v1R/h128V2DJtZuyyUvG2W6xPKiVzYC76bdGCv1MO/2HsKigWpO7r6eJ
GXuXq1ne8Rv6dvefY7vXPDs0wnAE4mok1tIssrxVP/m1W5WFmWMO98wXDlrYTCKE+0vKHzJbe7Qw
CfBEvqElh/4qY6tKmxYOPkN7/IwA8NW8FmM5sHGoXemLLG3qlRPRcBekrEyvJOPO/58w0BT117KH
NFL7QcQ8YsQfOlCYZaJIcnRuv4dFsCF5DVjQGxH/1ppNaH/vJe/o57hjgQBLYV3TEUkHZ/lC7+qg
OQBvzzJoLsJ3NdtLKYheYr4N8CIVlUF6a+pgHN+uFzSnc1F/a0fZzUz9PTxMBmAi52hZQmBGi1d0
mTtd1ewzb6dSImTEiyr5TWSyx2zLao+Jg6LeCbqiaM9KzRYDmtT7pCjWll05QhBMxm+GlwCGMnx5
MGzM9aLGw/3SBMHA2pB1f25oAepsTTK3bGUSJC0tyj35zesneBRpCzVEvulrBjr3jgrhucVnhxBr
dlggq83QFw1UvjSSEXrYqquoNI4Shrdgh/TLPpyzCnR6EI8BlkCihWBdynNWzTdWVRpgRo+WYjf2
Rag+K90Qooa95xnUN07KqNfCLgmb8b5iM+PuyDqqblJObDzz3ie+Hm5g5/+K00Ej+N6goY+KNoPU
RoVK5dDTc9qqRgXtgkRgeQiX+CJEjVjDmzGsonXdGsCmPhyM5rIvTcy8TBOaQhEyjBrk3ZRJMDiO
Ixnk8cb9fw+nsMi8R9tpWy51NWw6JhIdv6rAKJ3Xu4KRdRTENc3ZjAkp2OoX9lwSKWsG4M0sePy9
LTvtIECTUfSvJD8EuCiAVUfR5KDHX9wTC7qGoipaMOowJRH0qBJQDECbT4JwOGeRZ32Pq27jFP+K
uJGcfmvzYXWi72FNEHxINMbugPZGQVmGiE88beJf1vx6bEQzNqLul4jMKklWvsCT61NdB745x4qs
9PEy9lY+aRJxMK3QPGzO37dLBkvVpgrdrQUCL4gg+8I5Y7QZxEM2rZGgLgegQFhnFTbMLdY+u8OP
TlhoNRBLVC1jc7xlRRqEY5M5hLPEwb7gUymAvGY0alc94HKLgrCTSfO+xXrgRevWYwHPNZgHQ345
71G4kouztAjRjymCqOIPCJX2H7eNjymWue9JfWzADPd+fkXMw/9kEwtEF8U81JTQsN4si0eEogJ8
R0ORsGuPeWwR4MtUIol05/cv3Q5Rr61xbeUC5IEacgJTLUePyWpMZWnZw5L4KCKLAqHbiqkf0pwu
QChbiAEx7+Adv1ovxi4AsJm88ZVZ2vRl5OZhAraJQtvNbZpizlg1mCoFNlhvdGoATIa6WDgLIqpy
16TyLY5iwmu+SSDHznWNF9z/nnzsGsLvAlQ71z0DSF/uMFx0/CEV2WdMgzkQebklmTmEzWHJHB1H
FJ7FJ+oLjXNGfPPoFXs5msx2tyj/dk34LBAumZJ0gKB9VC71ppiqVBZQRiDJNTfbUNvj45qUlFZZ
gKoD8Vbm0RTtXCRRaWNz3pm6VJ31Q1Lq7Ff/zeqYOGe28/3Ju/ETGJ+q8nylLwcmU9Un3wPzYnhY
7whGEgamUrREruDGwQzKQk4ULopT0skj0p9DbGxw/+FK/ZR2rNysl9MvkLEDDoOMgnjTIknJqZjd
MiM9g5m45ydLma0bEBFihQXyJismLjb/cKIGR/eaPeypDMDuZ5FsqjNWxC8J7INYO8WfZunl6mtm
s1se5y7lFQ65PTExKIU2Nk/vqaF4u1HV6aYGabJJCdROFg8KEXZXNbYOfDZsk1cxfVziN76X96GL
sCy5CZJJZKA9hf3pJPffckxoYfYx1HUXqTT2bIMrIQNeBkux/UJybKdaKxGDWmFnvjRXulg0EnsN
7jthMrT5oPiNNslRXiNkwTsEKCXLyyXtU1aL1pmj00jPZaniFg3dEWjZeOfHm64lb+R9bdDcWi6c
19q+J7/35mqtxQqDH3l+gn7yDZ0b9wxPTZ7eER63RQBmFinvu3bIBczEpgWZu7ITbYyhms0mUzMZ
fZO9eNE/dWaah8IsKKIBjZSBzAlJHVAD/EVHm8xaE6LCpEly9MFQs8+XC2hZu23gluXtJ4nrms4t
kuFgSKbhho7uKXr8pXpz5hJYdebkwZLgAlaiTsBHE+tkVI6IY0/JrYcSd/E0UGx5XF7PbjsXoNmv
N7pUh/0T5wrjo1+NzZOXhj723kKQfGcT/mwSO8S2R/Ozc8/7Ly5UaDvG0BJDdGn9d83HWgl6p/KE
qrhF8vfJQV5AjjeNpCgx9bf3cMPwyQBDdEYifl2DkZdGCV1snr0O55Q5AkE9yGzFJ8yRdoFS8TmA
nHYWMPJw3+y7bX/D0D/GWatMbLuE+H1IPFg1YUcyWY32hD0/cEysH1sJy9QurInanzSOJcTr0RXT
RnY+2DbvtE/xPjwmrrcELCUjzFxhyC/sfPnx6yYn+lBQG73CM9aL6GbvOBzbQNlnx3ZtiMzMg8HN
I+yU8ZJHOM+JclimKlEYxUJbr1pB6GPCV6oB5qeauzNihPaj3rc4dzB+L7iat1bdwgNIdVv7V4Nu
OfDmkdPRLIz4OSwm4zCqcMD9Iw44siNz/d/cn5Tp9i7cChvYALlLzGsbt5Nzoc8CpLD18j+jKrp1
Ie6M1dgZYIpjJHbGMIe9GYUS4NCekKaT9cKTBu+PRQ0T9H6vJsNLmlKoXqUCIqDMC5CCPFwrf6zS
poEVePCX+h47I55t2wFcAUV8hUD29vsf/r69aVvClYH4Rskc4GViTcP4dAN7JLMJNLfdcBSqQGcc
yy+fQS0ecpvhurOJOEjSo1tlFPOx8vp89OghTMd81Lb+//0yEIriSn3z/xwgGr4lhHrRxGlZrg4Q
e86wzhqXndOYmsY/67iFo9WvrKD1+6fJucKw8Di+5adQG8tDlfGrKiijGVFwXPpmzkezo9dUgcXy
grmh8GlfugFZxri7g1QySBIXSpOuesYYQgCnOoEjBRS75vKSnBFGiXp+oVrXyH5ceJn7I8iYNm7c
E/ixrFH+eCAu4jogMwJiKgBgb2V4TELTt8IInJf2LDnymNuu34FLRCyCH1YK3J+Pfb1M1uAXjlRZ
qxqvf/33CcwLIhbKlbA4zTYNEIbmRFP6qLIw9aVFsD2FgUZIz/tGoDlgxBJGIWwoOzxiOs2i7wds
10pR2RvbuxuQXV6LKLDCAdq+T9HFXzRRT1OKwDvBW+rxxBxb74ZLDROOYNWA8zar07e29LFhDg0S
kIwuZdyJgv5qp33HVbuw3st46SaodML/ZqEqHjqDOVME+/qltoSgjwzbLDHnZ1fzepmF1EAEoy29
qG09UaooHsVYCS0LZeepzhpcmXeSFGXNM06TBStGh0+IiSnS8rV+TmiY1T5m5KXg739y2sG4X5jG
1n5Qt3/XWt00+Fwf09wNQ66tWbB/dp18p4nKjT7bb3q4U8iS/vHM50gljW1FjXGx0hVmPSZreQ4e
JOMSmmnwPDcGMHw6tB5z33j603Jm56x1IURxlaYYDOrBnpUH59Sq1pZOf1SAX61ZlaDaTadnZAfM
r7MoTc9aYnoYYzRs4bpiBjSiX5YZq9bR7UPUkaMBvObiYMPFSm+U6FCRh6jCD2vGSCpsSLB2iS70
uZdHs3TnLYGxsuaWC2XZlGoGzfsU8+UWsp2mnOOIFpaDdDnQlP7tNJh12wsdVUpYT2lvI0F56IEX
3v934OzW3x6W2zi0gbki3ZJHbbS5L3ER/vUmNTWMlFlRJULwlKP1qOwqiUm2Mz29TnBN2h85yVM0
hVSzB8YkRJ6IuxBlkM9hHNKxDd2n7CRHczylDHCPbyGMJ6GggA4jT8r/s3jFXtGApnROktsel/59
cnrhckvyAP+ZQqcKq/0+9T/aq25QrB2AN57u8hiPWw5oTGP7ODcIxoQXF6vlZ52JxDmrN/QxtpZJ
dxmzzl5QEIY67g0A4Kds/Me8VwfeHCnBn5ZkyxqnobxIaFkjLse8yvROc+y26BYdpEBMoLLuKDBQ
CmbwwReB9PlTYwuFywW1lSx67S2R8W17NRVKCn9+oKMYjXMfvKm3ORq4j+8wgO4mY/Sh2dji1AXL
Wh/ijC79rXi+R7s403/12O38bdATEmxmI4MpJjnQQDmDIcELqLr9Haaw8kY/WwSb/+K4Jj6bUd5J
/kIIPlJoUupajUwdvcngthsEh3LbpD8CyJUOf7pePVRMwW4zLveI7gVT1t8Sdh7Tg/GnYQTMl584
ZsKxp2VKBvdomeMUJGe+3YpF+ChleoeGxAr/S027Kra0vGixUMWTmtAROkX++/3qYJ7zFfamZnuY
sGaKeqJMAwQooQlTqZbO7kcpSVHhj/sB3t0CgGKRig6fF9/bWBtiHC1Npw1XebKWtQKtHUrelC5Y
1LSETI4Jn43vuY03hxd/OMOzE036DV/BRIXV2vsMLHHBnou+RWsxCjvDVq3Sxta4uJCKO52q+XoO
aBIesARW+dZfez9FqGKl58VUsO6/UU4tz1AB8CMvm/ObD9q8Ny8qmR7VLIK7Zlva26N20NvTzkWn
4utGAM1GNDcYsAX7HKN3GwhvvfcjZGkZxSmzTUEmudJvsyXksEppd+MlzGSVD5Et+ot1sSvwE4be
xxaxqwdeXPE/LzvbrF76MB+XJPFQ6JdX5ORn7xY90nrsyZYU4gerKx+UXS8cqiaqq2qq5hfOV3fa
uX7y8ipoAiSJNgEL7MO6Nm/akXPCUIPjLDc63hq37tCD9L9j+CrrZEpPsZd3HeduJtGtEgrSTTNf
uMgmAbWRxzTtgXWh8662QyrhassFil//u2nibdrmLd8KziM862xvwr3c3fx4LWXYj63tOy+2d+mS
GSu327/F5ZAPz40RewuoCrmF/RZmIdmWBHrbvPgUTV3dVhjWd6yssUUM6SijpxAD6mpZzL2uKRht
jIgdbhqwnzXjpZ3cLSMBB0VByRBj/5iGzxkf1yl/b4j0E6AUIrXkY7C2psC7m1gpThLXZDbhmsyh
LSL3f9MTFWRvhlgRFa5wiN8MX/ierrTb1FubdxE7I+qYgci8XZEpDlPZ9JSEvtoPPbZsrLCvxnw/
MEFJ86CyEkFHqI0YiVDjn+1G4CYleft5GARDmQHbWdlftcToisFaihANCNJK7PqphO3iLOVnBXs7
HmAYdDC0My0/dcO58mv2fLc/5suMpKtCxuT32nQlZxRZXNOru+LD1hI8XadgZ+LURQ39DR1Mu3sj
I1wpZ1GiYRK84zxKgR0BZWj6bwndQ9r7ZJ26uz6xi43LOW4kDQl6LsN3IMxFHGzftuct4i5eQ0Fu
P6heJyn7pAL1YK5XJ6UT4blDAHA/HW5t+JoB+7tVxf3EUCVAIFY2P60DzcBKNmdU2GXxQQ93XQdb
Pbdk4aTbdkfjPljfp4cTGGFJejnPIpdYO7VExKY+kR+ILALJNGHviOsgulPtU3ZZvLNvg5+zbGAx
yHqi6daiPx0dfCFtsfAHgsZddkrtgcQmQYksNED6I+lnAei94/sUPn1jIVw5hIsXKlAEWTZvwuHF
5uV0zAYSUomgTYTtYwJCpyQ65TgQBFBlDn/UUJpPg6SYbWiGDEV5tmJNk5JxdamCBiMlJTw1huR4
+TzQB1ALGLuJ7X5v36EpXLF9sejkBLd/p5xGU6nLWwJTA+dyX6sC04qJVwLluMZA7Eyx++hoE4yo
f6ZkCdpxcTVOSMRRtw4Shj5TFuHvfcps3Mg95edPf520qjJuyv9MKrOFR59qf382wbB7izX5x4tN
XYV5S85+AVnT2sEJLZc3B4qA1oaXY2v+HWRhUT0WRtTanmL+dXaM/x+3EMDkffPhE9+ToC610xsP
Qe4SqU1lNBUJMZKgamo7MiO7CDhKjaGnRNetUzn+vdWfMJk2iAjjd+iLHB4psCZDpcBlogIaZGm/
XvkYAr3y/Steq2lx8tedW2Wp+lwVSxmpr4sMRuRLdUMLBQzsDyYDndDo01ILnz5tu3ovUPFTfDzf
l5sDVVdUHJD6Q1+c2raN3pogkn6mlzBk/A2agNA5HhiBqr9fiUeIAz5eJbE+a+TqMoLr5ZkFATRH
IdAliHtHiOY43+48h958y9Z0Vc0GZUtHwb+dtfcA/nq406PHKmXmh69hmnjuEjPsNwMWf0BuWw4O
JBcTypeAsOCr31QYWAQQ2iyDuuHPgz+BFcdznoNgXJtxFwbr48eXue1mRcJi3iGk40VJ2higeF5v
UTvU8PEXpm47ln2NzhDLbvGWtNXb+EvrZ9MjvmSJORyS1mDngSFGrQLDcEFf7UfzWMNWNAT8fcYG
CStQrX9mFA9vvhMOsXknHi6wUNIyATzlC6yCk10v7xvBq73UVle+DaQMcCwhX3blledC37tViNwv
0x3uRRapWRJsTuqMH4t6jJT7sYfVdsD7Tc2+vrWx+G8pR0F/N46hDrSoonaukfwUrVbikpH3BBwg
XnQm7eub7vJ+un6t86R5y4PN1qTbYu7yP2GYMn8ShdSM1iWqifvVtb9fEIcsswDzEz6zoDoEnoiI
Fd62n3GamBtVPgDzFV0bIXwVxsKoMcFufD0M5I0QdHqywAWihHmKwPwHobFLLjJfWKqgYIy2fzpz
G6RB28OC0NUCE3aCyPVwFDvZVSA9w6QB2bOeckIdR+3IUmUbaF0+HHxoLTnNozxksthCYilwczzM
LxIQCuGLvMie5aP/56qCEfUVz4/XkucbaN0pAeYeyZ8Lvk2ZY1YeyAzIuqLD4VG/8JpEdGzTnc45
1LrmKZrR59hfmmvR2bHPKauIdLrk5pRTt7v8lr1aQc0vYTxIai6MRq0q2wb/HUf7eJK90Wk3uf+y
5x0W/eBdtc5+l0MDUURv1R8waLJbHQKrDFI31SBEy1ChnG08vbEpGYWwimomJwuTgfb15+4FbhnE
UGs++DYZa1lLa85WPI4ltNXKveEEO2PVvDf2y8aUTqKUsXlI1kVYL85MZa98W9RMINptX555b+Fv
mogkLMwoUpSlmyUDyXtO7FLt/4Ju+176WIbtZJc24XWMJAihPq5eoXsEJ1WyUHsq/nLo3xogs/nK
HOqjt1NReSh4JNHmYTm4o4ufOqysjCJ/8lhKnN5iDRHXiNJ5zshrN69hKU9veH9XoO6NsxYs9GSH
yekyUGfYGWf8gCUENj5d9C2rCKuHUtMbq6K3Kd1TiBsiYkwYx+JX3HqU/T4VUl7MXDVBOhV4XVAO
39EOh5mXgj3v3gNFZPgLCH5k1h80O8FdpXgLbulj/9SMvt8VYvvZ6Bev+ILAcGIwWL2LL1cPhOit
JpEQKR+3lETCS8ZQqqgAZmFuyCSaycNb1Giuhzy2jwT1vJccdHuyRkp2azv/EGFK88gwYWZQVBGq
uKEx3+p1ccagLs/V5p5VI/vpPu+moQlhhYMoCZup+QoDWX6O35UxbmAbp8G1ACKThjOjrLjeM/4a
YAMRFMLZfx+v+VXAx0XFou/yXNtjZ/dotkaIZnNXc5OzGGPSp55NASzWa7NJhTWlF8JwVjqF1EbW
GLWAoYY2C14/xtO6s1ngKtzD6x4Fv5JIggOItoC+0ttpQEUK0ljVlkYjhbrPsirHL09e7gz4Hcqx
68hbkoKD5VRIJRkp29IpCTecAeqD68QW61UzigL5BOhHEtecgVYhX1BOG7C9O1jVWnh0oBzjTDml
oMHc/7XRhs32jG9KX4WR2qZGKzZM6wKjP6izhkBtb0Y/mmcS1xoxeA8w9Z4IyxYq/YQ+FMQAehPs
tPxBcAKPOOUGkXRy3HpBMFXIIh6sn3YZfVLEhKcf/BrKOb9UGwN3w35Y/YJmpQLxqlJUzCDlgseG
R3rp2pDH3U2I5Z8cwJltuti5AM/OlzFfIU8Qlih8CeIgm5zeLe6bwra9T1zF5093YdY0T4WxnzES
4pli7Ej2JFyS1B5HZ3HjvHuWeS14MezU3Zqo7T8c65qfKNOYsKPYtib/JLdl9psiPU40eB57wMqf
I5BzsBbuZv/lIV8SNG6nbUPzeSD+7Nz3sF1p9E3cKs21dIG9/09xNFuTB8CagJLk+6gqrwMqhRNv
6nbzbeOKv8ifAE5zotDlpMl8kE3Pd16+QB4lGYmEDAF8J+U+eG7YLONWnxFICFmQnrdIcmcldVEy
5raGHbfOm8whE67VZI/uXWbjYQyX3/OJBJ50ADqlBrQRwsAIVL7XWVIxY8ToH+jgCcSEkUcKDx6k
i0mL9G/WGZM1IxA+rhBFKqaCrCR13EebyAEMDBuZN/Hgj3aGo1zuJSVu/5/YTNqyiAeLrV9/zndG
rvqmFLhwoWUv0PjmqjrEehfgLa5X+oPWkGCHDmvlfrx7BW3DHHbxZLEwrFWhmekSna1A7VPVVMhC
liyAJvo8CIoxyGAVf/x9JIZvMSa5pbExWsF+dCpwvx0Hu+Ran4mOSwnf5mMrBwLmXaYapREMR1RA
MI5o2Ft75QYTloTAFRerdZDO+GYJTwf8220qBmMRzripgDFJ4j47dS6zaJfSh+gj7BmlHE5rcuuO
JohI60Nu79S/BZI7hixdxipLHVOMN1JoI1m9QHcFhExc0jmy2vqiQv8H516enXWb4ubnfW/TExop
BU/7Ar0FSfM9h4JAFlRUDwfc3hzDU08owGl6tQr8aRpS85KigqVDFbiuIqlMuIICBRzLNNFrxaqH
9YK02g+OSbmWT1ZnWsFLoltpYJrsX/Vn+W1ZpSrnOdrMDfx68xQczRfe9kkOprGWpJDZhx99R7mX
bqWTnqPWks/1fba/4rol6vN/ixuVZfiBXvJAnL5FZ+nLGhFWv+F0Ywvnwb54EQo72d9d69I9Qe82
OTVQYoezzifqKS3PIySu+g9ewMpK5FALuqOwR+TztZYbxVvIHvdnA1fI/RZRtkZ42GpmDkMMnXPJ
FF93L/G+Ca77zYn55z6AjIwwK20oxPGO2+cg5hua2fE6odeqahPwmVdMArua5p/jtFSgCpKQqkhe
C/2dg4aIZ00B8LtEWOBFH0L4UZmzx27vbWwLOsRv/ZlQMyJxGRAbu2RQjLUd8xfzWf1ccMEMp9dH
wIy92+VQOV70CmI07p4ZwGpt4sF+lFavK/YbhI2W2F6rUUyaov8Mcm4YVyI1jgJG0OIRByNpEJ1y
WzAXw++XH6lBjtzlmZAtsAgXWEDMKS4tTajCjnui0vJJFM1W5nU2g6VjmMUxJVFtDNL58rwEd8Dt
BlzGddxWkeVPG5nj4+QyDvt/C+4bESYb0O2GxJQxgv/upDYmPuvcgVC7taG1ip7YtLnDsxxAxOuu
gt5MxddaAeR6Pmh6lOt22mjYiblJVsPIr9Bs2lt8OUf0+Bj77JRGl94eSAxiRN+i+gqnpMZpy7dJ
i4/oSZndeiWgXxNMwRaDfmIy79VJLVqiOFeybnLSS278lhGZoR+Rl9Ifjgj4s0+U5txaSSzV7ZUM
ovIBKP9JkOhpI0t9IbEUcIFBhI3lP1quVhfVrXJ2Em4v3hV2pVS+1OyepUNv6HgmGn3h0ixcjfv2
QZzbulZ7ySKgwhk7oARNRxwnfSDAbgZJfva0rH/onAJMA0eYi9gsogOmIIfjRamew9m70ug6bqWN
+0aEvqYS+dXQYmuLnxWjvRCdUaMd3Qams0LsYG/2Dh/n8mMl1rhQf9ZKgZLPmW0bf2Nr6HWmjXCl
NRSQ5f71SBmf2f9YZin52o48pAwtmR7xZK4PzlK0hvYBNBIQQ/6Y8+uo4dqf7g+PiuqRc0I3XGHu
H2fMokj+C3o7bsXZZKZhDLl1qiPVrhji1imlyDbXwgWhWQ+6l08FUjtfFL/zmxc/7fh2M78sjx1r
VSR4VMh69U8zPfKs8yTtFcHd+d3YLgR3CyhQwShuqTjIiEOwIeYGCwzcrMWjXJrRzZaueCm7fA95
ejr2c8cjxSjP5Gb6rzFF3ttmss1GXnB+7miur/fDBuuxTb9uuqUGbq61g9R9NIRrVjzKoyi1yq2Z
mScPivbgSTtTnmiBWrgIfYFjg1PjcCGK8dOUxMXkXW/RMf+iwcNWq43KdIbSqepK1J8AznJciW/k
C0dlXslFL+cgqgSXoyVYEY2+bfk8A3rR0Vcm3+oOKvAI9S3rhsNYVM/Lp4R39x+HRTGvnfR/gksO
q6gkNegaM3SLlcE/rK9b4HpCsjCAQQ1rXMEb3bPZaTvja1943Mhbc0o6dqYSkYojBE0VI/TWm14E
40oh2QXlujz2/VM6hblEH06uh+ajm1sFTh87n5iUheKY81M/Adro7W47AzPDfUeG72ua7mFnzrTF
khfUVA+hVzgU11jMO3tms6lkjcYWy8zERlRjoC+SCLFpet/QmPvqewG/flfK8me+wVgMlxe2VSPO
KbvWyqXeSH1ax3rYF/ySJAvtyav2UMbKypzsj4KpOcNctKRZ1p2lX0BvZ3gSBEMGSeZ4R63rXQA8
mNDmUkoNssjZhqD91LbEHiKc2O7ISFURRW9/IdjSsPrWAYNOtRhvyaJltjI9j32PT7tubsuUIKmd
gbqiA+WKuPHD0DVSmhZ84roThK5bwSflVfgujAg4SKSwg2lJXxcbgenWIspURby8098SBY/Lf8d3
QQnUt8UnLLeeqL2/d8D1OM5BJTpj+HvTKlRcBhBc7nNyZPEl+NNWQKc9DCNcn9T9baUh/eSoceJX
ZeoMM3nbmd5lyBEwc1F4lp2MRwDJ1/WinP/XV1rxfwUQ/uOsAxWWhki+bBuEqFbgt5nLYpN1SBpU
fO/xS8IvLKZXjdd9Z98bz8NUINfXcy1vMCY7JoPNBJ7DEKRWTn8Fgt12AtGKJj+qAI/a4lECI4EZ
IpiJnhAEYQa/OUYVuItRXS3Q++fVg2b1sPFuATKZxdrZFm1OB9VXCttiN7oTrSfRbdGR3gF0x+kP
sYmH0lyJKsGRrlyRHppWHspQgHfu2ZEEg0pwydQLVbu9RS2tkXF8eRnrZkJFD96PA7EhvP46Maxt
5Yplakm8tljaQWq9aOn/VH5LPQWtgXwKRtGdxphFoEH84p27LV7H0Z9CNRh5qOhCuHf+n5qY04lv
hwrkGXtFHUuOsXc38fH/1T/4BjdLewYIkbRF4cFeyAzpO2mMijTiJbEjexYlxUWZ2QVvse1Ca10W
PnCD1jrtxLVzcsFvTGkJVr6Qly4KTOwwV+6PNCWv6tT5cVQst45GVjC5iOHy8vhWNXXMZ12LJF0c
wSSPbfd6UAvya0HAjlSQN/SRZ2AM5MVvJgQI7r0cS5MummyuNQpok87SRit/jDm1sFlnCiqP7tIR
7NFyVjgKMr2MYexJ/mJSbV8mKZOrau927ruPqp1CFjPD6O9jMz7FH7Y4Em+p/MUTGfuyT0e81rEX
SBDGziCmFyxSvy5vjkaqHSUzJX7ggn3rMhsv2V5eEhMUzC5mlM+ylJZSO7/FjPj7o9fS1HurYgOs
ZUgn2wqzZzGhUNgMlN8H/iKxRXynabO1vPka5xP57L4Indqr9NQL1j9VloI85NgppbJ2PktzID2d
wAlmOViIo0VAhG2oYmcx5w3Imuy9G79QsOjZD+NV4XPsswzjWQuTK+NJrL25tY76zDpYBeoq1gHH
LNAvqXrBUPEKkWlCQBXHB0z1IowEIeZxZGjlF4TWE24TgtrLyQdbfd/V3F012Fgq/lE3htvF1h8j
7ta5hPB3DptLoBkEDBKxHScQhUk+Zjt94kz6DBtp5actOKD1maVGUhM1pvQ7Lp5GLsd1Lrn3F7+Z
Us5nzdv7c5q0Gy+NAtvaxh+hsPhYqwxL5MaSeJeT5TFaZM11Q1BOx4JLSHpXK3zfMWln4S5PYqQh
pT+fYg37rJSkmM6zpTVMPt7FH5zBnavfYqoJsjkbzaWmlSi9O9OrNZ57AQ3aEDP91PMj2YW1GtTs
O2SzDjaCbL0IhRmfvFJ3iBGPLLweEkYv2lIk75sy7yc8ppGCLDbGK9t33gXc9CwKsuprnO98ekhb
/DLZmNIAmT5eCJjRggiPwSQNDvYRZfdZKXTRffxbShkEO5YX8CB5//fIU6WlFvitq/qh9THabcTh
J5b3r29zSZtJmEzxd2aUikviaVB6qG4G8B1Un8VqcMjH8hejZ5MPyW+aUFnFLb00ZVtkK3pTWtUd
U8pLGw7OK6wuKt0IlzzUoPXHrpI5NVkuj5cWomuRgVHn7El4NLKmusOtq3+Fq4//Yx3dmT7bk/HF
axbkFFHb4xdm65rvhro+JQOv1CBp7rpSVofAah3xLQebFHuRReox+b+J+1Hk27jvuV0m7/s4Jfd2
35Nbsc5JBxV6nEb+1kmVjmCbSxkOd39aUyZwECtLW7TepLKp4QRh6diVOUgj6N3QHbb439rPvzlH
cAsjfPu+QEEi991MTm6iOxeozUaFQFMKePzjQnVDyvyaLMR5kDuGH8nu6yObC47IDwiAxVD/Q/+N
TfJRmycxZsvQDHwMLN1fQ5KHt2qq19n8DWEzLU1ycXIkEMwEciGvlUuVemAXU07uGnK8W8flzXs9
z7sh8QFVpRext+L3wnllAkfAwZAevV3m6EYmFP1id5l3ppYMd24JFYOtjbnCg5CpIYVUeKH6FX8x
XgQrSz0ac300bdlYWpHyC1ao2pRo+xG6wGkk66Zrxjfo84OVS/8lMLUNexN+6N66vCjaal//lW/R
qY5GiaAR+krMOLCVzrxTEdG4Hxd/TApNuoJLAeS3jrn9YFw/C/w7BGXfqZ4OtVp4T+Th5TxBsx2U
SE3T+jbm3dmuP3HiRRsbKltP4//ElEyEylUIIsthMpng4PhWrT+rjIAfks2BB+cL+45u+lZsIRSa
J1crcdLvG9s0xEBsRB26ZW6t6jPkPmFBohVdw09dQfmpVC+ZCTG6Tx9nB1vo1dHoxrSMzQCw4fyA
orWQCeF099YzTLNbowvTyXPxUuFoUG455mG98bGpvqB0STEGQ1AUFGhMtkL3IcNUTADbP+4M3wCa
0Uq3YAzcEUIg/38shZRWSeXy/SvkvakjbvjZ5hIroIYt87UcFOZG48S1CTeHfugAevzE3KdShlhR
xzhBCLyXpMy0E31Sng6omFEtF6M/Uk2UOYrf9DlIduYpNrN8RveggaQ6T9pbF414E/1gDJn1BSbD
LN9fPeczKDP02KW9aRO+pXYrF78IU5AIzvp2eLAqul3G/6DMV3LsvvxfP7ephN4mLbNvyL3Qp4GC
NHMZUKR7JBCuFdz2q5PCXiDFnAaJjqHZHfPb/37I9IoHns8Y4s0ApwIxBTKWSOyzvK83WOaHR+rz
qHFSm3dU4FNNEUWvK8DsG7As9snODxSyn+QyAYdAF5/877mXnWnp5mZyK8cY4n7asjP6wHazU8NN
CKBNQYcZ2htOjjlzfKFXOoy6cfk3M14QZV6haNMDVc/mV3FlgBQlHFFLLRJizjIUZNdCUMYMp8S6
yMDWYI1fSYHST1wLbw9HwO3IW8gLx5jMdzXUaJLZO1acFlQED0B7G25LpytlzaeVU99CNTPtuv13
W2i1JefxBKkCgNQ7VG9L1lFdeunNdNb00WEZt6p0p6/CnIyXD2Qsp06XvhTk5hQmvOMdkAD2b5PI
idmEna+Wk9unuYgjmB8OnokG42fKHii52oEZ3jtjbA2v6MIEDOejiVY1EocCoKdfOEpielQb+LpX
U/Vr7/oZxAg5of5wOu0hfoEzXrRaTPEMUpa5YUSptO78MnPuT6H1rLepEqyKvgBd+qsX4HEQZ6I4
Ui6ZEYvaCzre8kjfWs5HzhZpETL93f0XdehNi7ep2FuGRNX2XWVt6bMMzV6nYHZLCQKUK6u7CL1e
7UpCXhXWtakVEQ58ETzl1Kba646DSvjm4hdNvgghse6CYSFxWb2O+2icx455DXXbrZQUOGcFaU0s
2gZUH+B80+iedKocbGFPzboV6gjtlXHY/CGIDxNC9PtT55UgYES3xktNvY0efh5mzE/MI+Akj6rS
PxUqzUXdC1HZRSXeDlfGZ4iFVrAxzHt8uRbWtIKTLlroYhNlMYfTId9yAn59aP1Ec830Agke/UNx
iLT2Rj6ebVWBI4qRQV4iiqoR9Kwy+iE0B/oBi8V7zKr7DQV7GMbKx9FT/ft1rMvTpIUtHeq6/lq1
0iLM4YQBTXwEOxpcOohSvi7n2DrwHzTy1axRpJeii4MtMF8cq56VYarhO185LiYfA3HbrSxtxYJk
TOU8LG6J3K4S+xAgiIsnzzDgmNOBmw38+KaIcG99p1/UdnCTSYhV0q/pzFRLkkBEiZ0//BonR0FW
oCvZ5RBFUsCkno3Vn34mExmLpwy0Umlkq3E1Q/hyjuoOLA8IibpM/aIK5TEHke+8Xcp6l82Pq6lG
FHnYTN3jxFBuns/QjFRFZFS07bLnsuceTiJiKogYLNoi6gfm+e2Lwpxh0IkekFehJnrpdEii8aB9
RKXqPRwTYnUDue2f3PHhS5qfrBVRhgFS6nt3qRO/rIM7/ZOCKBH494RW3PljZGZsdCdwVtZxANB8
/vZCQCCR/0G0bf/KrCd/aAUAXwsGia2wULLMeSDGqFfugYQtYMf5jPM9yZNhSJKa2LotHxVFWJNU
MDnNRqRBXH0NMr5prNzrLBsfhMyyYxw1Mq8DrSSYzUlWbU+9UkG4To8zqUjbRtyws7NhHl9KFwg1
/VOZnp446Yc9s5oCpp/Jg/VrVIUM8hq9gDjgNI8pZDfq/qhjpInYKJ+dNaQAHQYJ0vWQOnD+hZTr
YmUxCcqG2SwYacQvMPDJOq4NDnUNHfJqIGgz0qRUJul7SjLQP4b4CP0zprttRZo8JleTl80LhL+F
deDlsCdV0Coxcb7nh11p2oGC2RMV11+4KyaA/BlTVQymzUoBYhr64TBWSUOMEiBYcmMktLl1hPw8
Ll2oBAGeVr9GrZ3FHDlzgToEo3khuJohwWOsv171jL0QQvibwFH03ZTRdD+n+/dyvVUc7Iev8sJy
EnndLVv8sYH5wqepOscOLuaUJjAQGh96fstUYLnnA6vfG8yvJzHf0NhlIeggc5nDEGmvhipzt3oF
6L35t7ug6ZMaOkHNARSO58exOaeIAixBUll8Ji8ILe2e0RJ/2kt6JEvb97eICPcssf+Reo/WIXfz
muPuDmQd8oBQUPFckYix+OQ5irMe8HFuBO4U93PDsuhfJjgj/yoHtPiSJT1g3a806aViU1YmqfFV
15cnQV8xVDe9V/Jep3hO1yRjtf8BIa+/O5WwHRTwAAPckiS8yRejxual12xQgK+PjTJBCa7b7Ton
2oFiUB+ibZL1wvurZcc8b3wUvjKLrB31cWMx8X+TyyYn53zSUPsv3Y9yli67KeI1KkQivQk2IQhW
PpwTpphGXxEBSv5DI5eqddgC9PcirLaK3EQRe8r0RWxmtM/lMjEqxfVyX3A9F7D6MxtICS/uAPVt
x6uzypPG5n+Z0C+Uu0gBZOS1CyXTbF8rU0S/oCDJvp2lmG1F7FFqgHl/ZHjZSmSYfP+Rtqzq8L7z
lFMkKK6neP2VCL21rJeD4Tdjrm+PQAfjtI0LPxOlWnqTcRlFTuG93T+0BoYoWbTJmjlmh2PeCSyf
7oRPuojrYEcUbpAaLSHnAJ596Ys/Zt32F+j6CMGq8j/3MSgxD/5tMmwGwgld1qKQoLOmetqSuOUW
SeWhsJu6rMsyRnZCQV0lXa5g/+IFk97Wv+qPloS5SlLkTSYpMyw3Y1XmW7UtsFcdyWsGSzgCFY2z
TjZbv9Oaqe7/eHmlk+YAgcmkUTnF+AnbvWTHdeaVAQGqNWcaBti+DNrdwtnpyCwy5bGSzKwAxNJY
n3ffJWRabDVbpnvLvt1/v9lbP4hlltcXr/6vQCVGCd33it1JAPPdzAhSClrP+HK3vFMMYN2pwkCW
DMQPJh+TpIHnfty3NAea4j2cmgmZIhmWdGKGjNjL8y1H18TV2i732B5PVud6WPFiGZ+mlif9W+LR
p/2Ro31ytx0yGQRJgflALoEDqgYzhFFrxIvkzTfS2Lo5UTRWwzbc8KU+YoYwsdbBE+KDTUxYAT6c
kJKZ0Z7pz9o5ngjwX7l0e+2jcOa0ySTaWpMmDIJS/u+o5C+NMgdTF55WixD+qEijgR94zD55m/XA
rDasbL2C+dWfosX4FjxzvKSkQLjecyWRDFt8AGsUzyAU6rR/YYx5JtSBtR5Bn7mlhaIZjaSsar0D
QE5u3gz9O6wZkeBNpLEOC1JcPsFHsZBdAyqCF56Cm0ElMzMQBbB+zpX8ygTmcibWufFosX9DA+SB
ZeKSTiO7/tAqoww5oQZNYweUH3jyxHS3JS3egeeGr8xmgSNsfttFn9qS33MFaAJnN1bFMe0AzXu0
ZVFH5U0HOMMtuBFjLyhFj+QZSw0wzeSbT6+Ol1RSGWBZDObrPXgONc+yk2bc3iB7OZDM0ozidYgs
FhQRYLwnHkW1gfcZbnOu/w2CqBFcjf7FdlF+Ct7WKWxqWJL14irgn1kNFjPklfxuft7+w/R96i8P
stWmRSnQVQhRYnw5xcDAbpBMCS5GQcx+adN7uaFYRY2R/LEchxw5ZdelifA+EjPG8WDnHEAK1gkY
xc0stQJmgd1f1bq0E8YWCp02XvzmaxivsCoakOf4B2oE16NvvlHJTIABwYLWxW/eUV2ueTVzpsMe
SRYtKXyF+FVojGkkNWlaNtOTI8JC3HqYW+7ZchRia1K4EQBtpeN3FnVr01WiGEnfhQkUz2bVH7nu
iJzt1cUls8TQVDhogePn83S6qVeAMJ/A8ebXJdUU0jX+Qy7Bu4j3qVe45idmruIuLeJ3yklVfVnD
QdJ3tSQFO01rnO/Brz8LNw/+pdWlVwlQD5QQYNjx/Fszt2WCks0dvh9BTgJ9TMvqMR7T3v8t7ed8
MMo8jzMSchKvEkANoII2zi4PVhqLjoQ1JYg/ZwCq7RzNxY41M2g7uNqGo7b2L8/OJzKWlN3O/FKI
w5VRJfQycR500TcT4G6RgKmJHoNVjzvkkLhFB+VrNjPhgWz7iRzb/9ppiYMZRINt+dW+2FT+DgnK
W+8G0nYPfATkXLwTsR7bdqxPyV/PWB4Pe6nGsm+TSVI9BN/ouWfdCzfu/V8+5VAtdL36XU4ZHYtN
fNfWhRYQJdxVIeq6syj7cALcwvgWjEBxpBsjvV32o+eTkCirtpErdbuzBHWXRiyls5H8zmLvDHyx
PCd/DqTwgTRM5gtkmTajEQ9Zxl6S4mEekweN4gck31JZxpysBJxdWNry5TzF+5nzhR5JJ9XGmk0Y
OpShrNjmTh0BlN4h6HB9ra1AJBBJoxB2Io+u454Vz4oZlJDMQOgwIvgC7tcrHJhd+eXHEQ6W1pB5
7LlcmVCMsI7ALQ2KWMtK3v1cW9S3HqgatQkhRLV25mKSf4QWMtrNfQ7ZsDfEmuLDOyB0fVV35f2w
vzhbFACaLfQ0HZetPa8IFmBE4xTQLSSSVu6yKlg3UN/oQLVLxJlKnnzXmUa60VqANeFIdip9HLtw
3q+7bDWWZQiXwf9NIPrsMJJUmDwIE00BHNHH0Id2xwcaamEnyi2XBjg/CEo+HVlyjbjQVTJBE1Mz
A56K/LdIHLfXBuj/Zbg5NtsR/w6uLaDkk0zjo5cMVEN4sVAXfLFiKAziRMhNfcoKw97lg41i0lVl
kbX0GZ3iX9ntldpEO61KuN4yxlGI8vjgjWW2klFUaohyfohe6HgXdfy0KhW+UefFUPZJk0KXlgr1
/iMcsj1aLYN6746N/0EZbHCPyCuxvPQiq2Hwn8KiWQi2ZKldmYfxY7UiAnBqnIl+lUr2cbr+CUiR
isqIFwt7NgjtbZkgDomXa+JOgKQD6ss7L6neLXlEDvsTKsuuAmDIC2VIGlzPh6vo+SNjX2yGhmVc
WJeQfm6dq+NpgAB8Pgqs44OZlpm3JfQcf1JuHBeqnv0Ui52HSlmTijTJ3G4lT57lncG/912UoVAj
WDFmvrXwhJCcsa5z/9iljHAZD2k70limxxV/BQio7TKY8MioiP1tEDIi3KJgg9P3utzArG9oZrDy
rkY+/ov0E51mfLU9zbEyj5+ShhRRyBZRzZV8gyvhNqiskzfdbZNLuII4PtcJEMG0w32+iR87eIfc
69rBXF6l2pwHGW4w9Zo+01FLHaOtzVZ1BWCDTU+hVnhtRiIrtBDIj6kZ/Jmu5wRFeeP3iZ2Tak0b
O/zcLHAFDwsGR5C/WH7vCbWxZdkVYrNyLFh94fMQu1NYHL4H8OSi+o3qnOTsVZkANrfw5C3yMLC+
dFqO8wwj5xNsbBclOfdQN3JkF/9jZ2f1EMs9JR4nce4z4QE0Vk1IKItraO6hftAzZk4VN0qYAw2m
xx++Dh4mN11mMpiloXTpqhRSH44OQql7trdp5Jk3ZqgFIrZKZmeAuBsr6Ko0wZifFkB363wYgh8S
3Fvei0R8c6GaJQCENf1TP6xwpWpXwIA98gBbnXgmNmcex+6uU7HuKEsGI6ZZ7l2GyKgqmpsxKcJF
QlTrF2KxYMATwiBDBdIdLd+gBDKsAxeWpOAWB8jBvYUsHt4rRLi8nu2urHxpGasfLfsp8RLJqgX5
qJbyznJpl0gEBNt1Pe0oE3FFilQAh56UUuVrImLKcC7ranGz3d6gZRxWeideM6rn4uy86tKCiQAt
gFS1eNy5lopHO+8AlBWb/R2nif3wyqpFq6H9EwdjBQJmGg2AaGH+Pz0ICkmf+UQTNUTAyFclewPE
R6Smf5GkhYZ6yg9NLEPsj/hCaLom8O2kNB3CHlm7BuArXpBX3gny+YsmyJ0J9rUYBA0ov/KV5luU
fd8peKu4ODRgjcej8qyqIeGju3xgHjq5bgjFEhNaon9uyuwiVMCiMkE3GFFTArT78xT5CTFCRBSt
zl656C2EF/P8lX2T0BXO45s+1wbjLc4SrqVWW9VADyLcMpmT9AefkJHWC6LmnCxv95mA28eGjqLy
DmgzVNR3SaLE2y/UyURq9TsEsSmMKUWNbi9378gG6QsS8HNxWRwxlMDHNVKa0aIDZCvxDB8oPr+h
Fp++iHAMnZc6cCgtHfjJ07shbEDHxV1CcbzU/sjYyoyK5FK8FJ3GHuhi6MDXvMbrhKK44cf6HJrc
zH2i3pI48ucmsIMhp0cX8bRioWiZcyjOeNPe5VyYwMvD0ENhiZMMuls/b+XoCG0xXw3roJCkVfge
YZ+KiXDheI0hVsSjMoZ1ey/EmlwTZbB88CHC52oTSgGd3qO8CfYRbv+XynBnENhqxhPP5Olyxybt
04NfFdzuNerUseVRvDGorWuZcCLA/ObXFGALHuoCsbq6F9B/VYiw/8NchkqaAlsqnu90Q1dZ+ENN
RnyBW2Z6hbijQTVN0ngtTZACdJmLocsrvn6r+Q0jQJs3Rxo1GfpJF7bUNh81WeN370R2X3E1SSij
1131Cl+tjo5hxHivLC2CurdwmewcqBDDBW7SiL3zm/5wzwi0ug25oDxRkAW6RDCxDMNc0Fu1jqEz
J7Cb2yTrpJ1la004fQLMAL2m1pAvKtz6miCDDqA1cCdA5UmMcAQZzS0894c6J2kHwig12aiXB1uw
/bokvOdAGJqM4b6OLJ1jgAW3RGVKwl+H7XrtPhhiB6wWzKkBJfuFtw3pW6IbxIsBnJ0hQwnsuD3a
ew7sDu26cTI/6eRdwmLimSNNGAKR7xU8JNmK627rU4Z5mDhTMVHeN81daf4Cc6m5KsaIHQa85eSR
Dy92Z6+0Ouum22J6z86mc6S1I0ERvTgsRDQ0IIHgNBHNDXAVPI3YA8ZpzidWhYxyjMp9RlMUGcvC
o2tY53Imz20XFLNHXRU12mCN+BzG4NmiFdiJWCQqOoYChEJAUKIW/NBO97/GBWf/KX9B6n+YGqpD
DGZaqoFU6tnv1Cqn4axt4hiRZq94IKQOjmJSt89PNSzXlO70Bn83oILCr2jr2rhJUKyOsXz0yei5
rV6jyZ3LFhDMRn4CrfrNHY1IoxnFOqQChDA3k9Wi5FfvHYYXha3L5eIj3I2MDaFqtTDKjpeKT9wh
i+bsFbipW9TbabuYxlXA7yejqX9W9AuzIWVHrsH8EtHkYY+pPCl0rA7FzJ1xO++YmmFBfuqZXE3P
49Z6pcJyZO7f9Qevgzr6ite+MnTw8/7AJnC+jUO7Tg1HG/GUPFUTndVcbCGANoCh6ePmNaEIa9rZ
YDSyNpxJQXQzT5JxAX8+kVUEk4l88pft9L0PJkYPGQh+SwsouUhoj9Nzq1QV9V3CvRKVW8Gf5KeE
KoR0N85FeIiAyvtxDDWPu0br9jYUN8dqA+pPsRJS8ZlHH7jt13CdyMd9FQ/OKdvio+wa4lhVdXen
jcZ/W+0OBb2LJ7+ImDdox8oiMCXGst4WioN3wJ3FSEc3oBP9acj2ZLekXh1j8tnausGJ6ZXIYsnT
SvHDmvBEs/3nsNtbKB3PhOL+nQWGwIpBYKq8FD/2ygXH/gAXtdJD/57Sc6vEJlXdcs1yV6//YZmX
7ZA0BtWa1ROK141FGz61GQ/D6sgkLcBQFXVMki/TeMRbkHq78j6VGQhVGL/IRb28E6mSIVmPOACg
N7FgNQ7ujwaHzCiPHozt1c1kzn6qEn08QXeSxJtpwF35KUKs8mOAVkn5UxlStRrqT4+22uJHMlfk
s5rxZW1U1mSO05sVUxLGNPIRQQfxE1n8LXDW1QIQYeOvWmIYEXo0/Dn5NseycfDhAPajsfz777IB
myVmuBYf3++hhf2iVSybrDl/RCv2l6WUVs97sMihec1e2S7rpsu/SYbuXRNko+hGk10/SKyHXfMD
D7Z/GZxdhByRslErIWKKUc5kHR8QpJfMuwTTJjEgBceOuVW/edoYPZexfK9felmiopXrxWzusDbU
70viw82Gp7EpysWk1ROQlDz6kqI2mk+yTpNs1MoUHoh4x2llMfYR74upA+ECJcE0A85JH/rto4ja
z80sRYzkKEbSJIFygpXgbMVmEn+Bi0GFylxyCB9g3rDdZSRai0YtDzTc5o+XUOjU/M1gIMzylYPa
dYC3KS/2Xsvy6Na9hado8Uw+refXbGlyU5R5eZiwrBKHEPzHsFl+uROMkSqmhZ80QIqss3e0oLVA
DFMTuGQZYQtNshsRRIQi9jc0OG7rAAfzxE2495Ylk6Q1Dofvgvp3zbHAJTUMu34gndA7osa2bZPQ
l4Y/XBOeK5JGk5RH5xutn49xOupdkLp6FIBkM5DdjXh1enUxWekineHP0Qs0ax5hejkXZhWSWTRk
R0Fpc6uwS4xsndqaS6E6m9ngFWI2v8EsETTg6WKMT4tG8cc6H8x/KvOJB5R+8WgLjQQSObHI/fqH
XVjZxV9Ah+p153ahhQOrcn2F82OYH6ZYKksDkY+ApqGRklVjavqopuiBfJBTQ4F8uMtfjltBXt5Y
VTRBQ9VUNmP/iQqNfzRCY0jnvXBDBDhnQjXoT7/x6XWWvuX0xKHlT24PP7X5F+7foBKTdG27IMfh
/vSILv4vErgxVTEkPpWkMWSi9hKF8nbfe33DHfg6bDHQMKopn+RL3/iBU108lF2gd5HSq8E8ZLgp
Y0L9prjbjPhYHV2j48f0raJqUSll5AY6V4pmT7MiGBI2I9KB1eP0KfTrmaCIIzE7av1AOllqiFKF
8cVqNyoszVKS/8sRuhxW8ZkMpTUt2CEJZndFq3+j9LkHjX/TZm7NxzQyuIBdDONvtQXS5TqpS8iu
Cer3uivrafMmF/pHOI1oV2bEaGacUnvLf8Ia86F3uSGTzvQtYimZbwrAyoHFf473mlWJiFOIF7kN
xvzuDWcW5DnoUb5OZrrEA3pe85WPfZknaM3T9eRcLb/++C+Kr4VMXH4JuFRQlvaPCr0wva0pZ/f4
rKlWyxjlhm2tFYLhp9dcWwuXzYsO0GqlnuTItt7vwO/cJOWXzUqRM+ExhYKWAajLYAwrOtY8980Q
opg1fxEVunrPl9bRWttmHZFxxQLCM9z7MedACQlLrgNVekjRfv4nuMQ9WI72u+PPzlcmCzZhrBI/
TCgORlJ9PSn+wIAdocEwhtx8+wOjP/qatN8Ls7pZPH2XQWvfVT9YAxF60e6LG55xdVTiYSShmcIP
fqyPa7avUPIO82wPvZa3H4qqQctlQUr6FE1cOCCdVOX9mjmORJg1HFsLcp+cgUUaPPRoJY/fK2RR
4He8QuIMP0uAW3+FlhVXw/h9Mrt8HWwtJ0CNTtJWTurZk7frFnrgqGAXCD5h79SgM6Irb2P3iCB3
IH3Ja9+U7OGGHryYo40C6JJ2x6K07xRGyiRIMbEUbCkp+DZWDmN3qFIrP2iYXhnb8lGJA2wG5zYD
cHFcp8bhCuzi/bAYpb6KW9bVUfhGhw2Xm+VFvEaiM+PDukzW5MXXCspnoO3hKVpbeLUusb4NyuEd
Vs2Id/aDHqx/GiCVp6I8H8U8I4OeeGDi5XnuqcOarGASIJZIVdi5qb8F79QUqH53lmB4pgMOjN3T
nOo5+Ltnfa30TU9JuKnXY5paw7qMvJHcGzAxH+yRXRBl3QSTTTbhiX2SsYixq0nh01CLz3k1L1WG
uS6RYh4AeDwN3Im+KgBExoxCFkeaWcWR0nyBs7qz5/4MkwHw+Zy2gWh7gt7FStQDOZwJ9Pak4INA
IpBkl/WT7qIzsMFOvWLUyk/qve7TgXb4xbxowikw9j6noUaOl66+dVVf/oIfEVgz1sJnQFFzTEnV
voDrZTiPtE0R6s0ctP9C0hWWdZpOx7bkHfgA+vyvQfr+iLvx5NW4Zx1FpZ5nW85ubZhKW0BBTFQa
2+Q49ZHih09G2BqGAMxC0RZ6clkGcJbfvsSwg6WA92GiD3HsSr8IS508c1PPinOkKg73QQm07gX3
n4k/ySeciP2s/ySvHyxOKsx/WKg8YJLQQBa2OUqPtYwwixXSH5OLKoi9fKlvwtt26BLcE2ayTocF
3UwhzSA+Xsl+etxjCpwzPATi64tlGkjK386N+k0xWzcNcIH33tk/bMEPdp2BTBj8nihsBJODXbUI
aPI/H0k/JwVH+zY2U/661vXPF43IbBYku1hqG2BZ18gzfiFKouwpVHy5vGhqiRexo3f36jKq1eIc
mPD+/5Yl4sGhrU8TNk9PrrWlkecJk9UReiOdl8WX7X/LaitnRmrHjmhKa+NuzfhRG9KUW2ac12dQ
s61GQ9JRWM/Kudn3OZHaUTCvPcWruGda7KpKnkUTvQYgs0sNAbIYMoz0LQ/6RhysRAb2gOdEfEBr
g8MQZ/dtWvCuWdzj7phWPoTsYJT1Hv3m8zoi+uEuZsF2ZjAHTzLvGGdrAkgND30OGdHbVjso4qpd
XJ+TSN9s/9OTr0Tdp8ME4sa0JJh2HjDJ1O1iugd6xk3Y62ILFOoHFJFN74npYfSz/ygBL/dttK1D
3OgjEYwahuwH99H5zNt/zEgGnZtgdl91KeXaOyQwuh7IpS5W+wSw0+/SXjNZJKFVHPOhTD93OWO0
J7Zk1rKFm87W7yARZzG0S0Ss0aRNcsgClKOsrbwrOEz27Rgeqxz3+PlIhtxRwN4QeFKFgg2zEQj3
wuFsjKhv4c30dMqe1Rneo9DejRPQeFddeDfoYyYm6h+jBsXhfmS/oI5BzY9GZpQ7rsaO+2u10NGD
EOrbpWApc7LAvH6OiYMbTZ7/DsN9APa94jFFA2j1zhDe+qbPbmpT2I/ZxUeJYVl22Xk3HaTtAvOQ
jXK4zPcGoWKAci2Npck79RD9GB8qkRN2xdrK/mXrzvBxrRFgI16QYvs0aH8HRVT3AXK8SKsvsxaj
SiCVHP1L8CWX9W7UAcDWNhaehP2cMiEN3qIXqSHkRfGc3QIx1pwiOkEkb+CVP28y0ukJ/CWsMwe1
ReXKq1FEABBgF/VcRMrabbfgW693yCgAufJCdC1Dov0LT5tRrIQuax3Jg7TL9f7MNlNMfZhlNSh4
2FP/yrRIRCgL06JK7/VabzL1UNLO4Y8kNlbMkyeVhARA5iX7nubQhKFqP+VSPIIl1W3YdNNMXB5V
4kuig1GbzDfLrE3UrsUjLVLHxMpkMwU46qTjUarxsiqLUyEMSD3r3CASZP43zSnVVD/812otbqPi
laH+DhaRh7KGdTHlvy63Zb74H1sjnj53urS5nkGvRiqVnVKXOq4WG01FjZlDZjdFFkUcvhwwXqqQ
k24RmvHs8/xWh9XJtX2Ujz0CCdEPQitRfcZp0c8nZDQN705xPXmvcL27yOAPLv6Iihn3QPCaKnit
jKQm34FaDpBAbvfRHy9ZQfmEodl4QuT14hEfji/rbOwlrJEY3DJKVnhqnflBXLM7pHunmkPdKejJ
X/uHQ73cq2ujXAqHDYd/N1to0d6wm5oEzyXiOWK0CLYlemMJZRB11evDQ2NyFkYh/gn9ipE2d+TK
b9zl9JaTRQXWv85wv0HVulEtWWUr4wMioMpGKW/+dL3XXSlpvaTYXjFDvzkxDfqvx/Hemyu7KE5h
omBaKWANu0siTY0KkDtH3kobm9udLDP53oQuqoMODsqzEv4hm2LH8Z8DmQFU2L7J3V/kLjhabSW7
oXzwV0sRSISCmZeklxF2RWUCej5acoTzD5gjce6mIte1AQhko9TjsH8VG32cuCYWTTtoXBxRKKbH
8tkHb09HR5OWCS5+pz39FtY96hxcG13rtDvtRdH/xFUh6CjppN9GbfkZL9C1NcIEwJGZ3M4hfdy3
hCN3ahW3fJ4Z4V8w6WndzSkDr8ytUiXluL2D5M1YZwEL5rzQzJzs2LhDu2Yz++EN5GFJmLVjCn+T
Cm9N5fKEgmSJIRNREVea+ecsdhEgs1tNOsbTK7Tlu7N9UyAAdM+SwVaVhXLHRLSFq6x38oAJl+d/
pQnHAbKNMwQHIku2XSx7FPYlyqRdPYv4WMDnrBqo6daYn+1NMjN4c6nVnqLxSMIw0MOhLnCeJvdy
yAlLyTxkJsEWwxPAf0sg88HM6DU82ySIjzjGbSapwHfsue0xQ3fgkKJ8AtcDChYDEuDCW1cZSIQI
67fPeWop0DNrycmgJd+rVTNy3hbTchxS/6lNWgb96DPhIbESEgLXtXAyB1Lxuz7tBUpiP9XnScba
uA6EODm7A6u9K17jlCFeveagC7XJG49EIuNh6qcQGuXbLprPzpykFPzF00cfjKznfVwFhR/+nhFD
Y+FRYar2BtI4/lgZBJH8lGxYlloKer7tP+mAUYOLRTuCnZ5P/bC3CZBfs+5dX4qDQVM38E0bq84s
zubNFbitR9tcpnLL6oKDSS8cWPLm9bDpiRWjSZzAQtwSq/n0HVnNHG7bBISzvw31Ppr0alRto45c
NRIUTwqwd8cjjOm/V0yB5NXst6QM8s1A2CUPzW1AbykyN9xubzqT2WdmMwLAdt9+LcU7Z2Im6oVd
tzJLys9pNb2epFjVXT3qq/YG3rNK+K3SALJROWlJhJlgfXEJEeJL2iovPEr4QeuBOy/XrqN3hg4U
LTSTTw/CB+FPOGRP5gx8ohzJ1epDLf/Z7ag8ovy3PWV4j1qDd/F/PEDX43R0M6wzqhLFAortOpdK
NucUX0u/oXhfl1L4nWQ/2lUz6W084rEpukKhFWMWwF/+xqpXqweHZMJurwQ+pIW2x/zMMQfT3+76
gNv/WMzkVrnwtiLuIvaAuIt5NJyojdVLltwN7ZrxkzJ7nX15xkY1yA4y9LXPubVAIQmNptXRUPd+
tcXPfz5KtIwRV4Vh7DQlqGl315vWxjUwgvTYLbGZWXmCqQE9fzUiTtXps5Ps7BXqFKOjSumlMkzj
sKW6n4pzHNKtBIXN3BoeHlM6aPTsDafkVast1vNd5FbVhzquASKXd60EHj8nSeNnZ5W1LgY6swZi
N/2lbY5m0NzdDuYpVUkP2UGIJKQZhM4qSZa/MPamJg8zhHynb6LhfVerjDuJiFM5yvjAMzntUchW
1M0jysKbiftp/zPRxIwjkxj6yJQkDkEDNQayrogISfsC7T59QhD+vFNA8Ce80CxS07SDM9xz2eSK
hSjQ8+YLUa1KYfIJSaYQhXP+qD3IzxU0/ja/OQUW3gih6ZMIjcsNvjkMUN6gE+aZtvCTov3d+p2b
SwCKFs9lgp7aDFW3z/pRmSaJaEMBjFVF7PXuB4MRpr73rfE/022w91BwWLmyoLh/JsaOjuFQix6E
7roHuKI8JCwutEbdwINfhY3pkfBqhYHYg8xF52OVTP6bMcsZuFSoihbA911UEUn412RQhcdB1tZo
Qa2hDK6BnGDD2XwhdfyaoKe0lHXZRVFjca/FdwXwAYE1KI516ldoMfR9c7I8TA9/jYyAqxi+Thmu
Eyy4VD0LKDfBXXRZd+I/UTiSxUtwnHXiSQT9T9owDtnjXNGrIC2ZrFQFC+9e2iobRVHBo9lL1YoL
9ngrnlFkW8yzCVkB4jdeoqlj5aEn/Hjh6iMb8HbJb6m9UedR7maIAlOG7/rwiDQpLZ3cWB/GEcu4
eh2C4iTLrrfVY4+cRmrSoB881xeKTtDAw+jDlKEE7k5qxnARzqM1valpZfjF6Zv2lL3m0RCHfxO4
AmjoEe233YH7EUhFmOvdBZoK5wfe7gu5bIUngi6mUZrPZun2a6EfpBWjucxNCRJk2oI4tnvKGLjB
GoP/SUGUn9FjnhdHr0B6PwuYDaliVUTz/x7ITDDaYUzKTy3R4XqSdC6+d4oz2H3d8LZxp5byCwrT
ou8o/IhkeuGaRzd0MmjvVVS5ESrR8RkP9bcstxNd+bSwiNXVWRSHTuvnPr9Xb7tIqUcdIRT/u6Y5
QVHigbSLtELnP7DiGpVwHg1P7Xq0iV5qKhgwFkb5B+50wpi1z71Gj7uDnaYMAMhMuT4Wo75e13Y9
4eOsCA4a8ymV6KU0mLsQQnH2EP4mbK0qT+dNN0+1yYg4BDtl+2xoH2LpuSvaRoiejbgd0NAli84u
OIlSMCo4pBUKG4G1di1XnKuDJEogiMe0dzKuHvELQpqvrDpESFz2Bz/7IPzqsSL0O2lnk7bv2/Nj
sqA51A/NVZVRfQz5cSC7rwNSuaBq3+8co3QSyIsJWJX6gur4TJiaZonc8RorS5/wbC8sIq+70uDy
eZ3CBQAI4uUtXHQn5gdZWnjeOGwbU9R1rcQIKGS5jceEEn1NmkVzASwOT9fSjiiMjRx8LLAPv7Uu
lk9JMwVgnzEkDKUrourwYO1Nb8NplUy8ODOz/aTspLuoEs1dAp7URsE8qoUM9Bh+CvSYy7jnhQgI
z9nE5TJBrL3IK7CEuOWPLXQu4TNhrUiHTk6gEzWWNDej+bbHpuJik6aAdqQY/L9no9l6lzllH0pD
uccPlZPhLBEnw0msPULS+UPj8kgNToG0566sOM/PsrzafZ/IFp66uZzgNUXvqWGB255+6+sdDDv1
sV2QD9FKZB4J2ThbqgJopbTidKovLB9BSeQRpfp3M3ZwwFdsDK+Ra+1KT8INLVCCA59DrMAxLCFV
gQb0jOxj2E+rqkn74z57ijR1V6jENgJAXMOYcuSONg2GC+AEWgnrVObDgsefqmDC5urIaHy9zxje
GRGlidIJaJNv+cKIBMHEw9bRDVVokCkedEEbz2fvElboh7C38TkkazQ2g3KgXQrr/PztFAH9QVer
Pf3PQu+PFz+B977P9sRce+O0JLWLnbkJ3zSyzabobdsbXoMqxFqXT2RFna5aR0qrP8e0crZbFmbb
bWanbW5M5W0f5jZN42o0l+KCIrqBkFPgBod3z+OiWboPBbBIfB5BZbirqXLZyNPNte7a6UiwEsdN
KZ/SQw0exWj1XLCj+2LD7wBohMe9A2zng+aIWzaqbl+myRdgXMfMJRDFPsyH7EpMk7QW+zfOHIzJ
KAQ8PWPJke3FJfmlZqQo99drYamVbLFMuirs0ScXnAaAVEfQ7EvorMb6GeDq3HPQob4ZYkNa0Lvy
5NcYR7482zaCxYgGiBIPSXRaaItULhBjK7WLPN3mRFpg91fYKU5zN8Q+1CHWKnrCEbwKekq0hkXJ
SeVC/HdWpheRZtoIMSWRiOsb8zrH+PzziBZRzIF5SkipkKbF+uac2SzuOpn/TRgf3B9VBzJhcc8z
flPoemlrxHWFxTGHHZ9opgLjOQr85UqfSJHCsdcMFOJyW9X97edntKzjY8jGkffSYUyZnWFVMVj5
yYXyki/k+sMgCYPnxmoPdvthORQJgLUr+P1XJX7dxXXIrluAYUzSegZVOMXQdGIIyCjmXRDvKC9v
d4ok5tTWl7hKxJje6x6lgQHuQ68KjIumYVOUmDt0aoelXiSEK4scBRJaieYzYqjps+XvBKVFGuOw
5z5BW8H8QZLtqZ1EBMWr8nnsQoYloARWvWkO7ER8lWABwE0jurLIx3qp/g/0b5MYErZ85J5RtMRp
nO9ID/I9t9YqdPDgLC5xYFrGzZgQREpxcESC2TuHPhARrbeJQtkI8gtlo3kf7geJN8UoerJsvBSY
SFgkIHAb7/gGk5cXE+xT3U88VlTLOkF8v6Jt8tb/zTJdcunzhkPFxNikRPVDWn5IkA3xrZw5eEuL
RhKC+cbdkuaAE+Iqjyt/PPpNhyP7KdJsB/WohZkRwAsYX/xvgv85cVSo92q8uwKmRhMjaDnPXJLg
upxgcuf3Kv+bI9X2LEB31y3Zj2lAPIYXtlHflKTNXjFQ8UExDeVGq253epvwE0RpfnKcqreZojmV
JmZSbw4eT9uZpg/zXgubbJH4/hZZ631ypclyHanEgqbiHcugZ8jQKm4KlMrTFo98W18MkMJMFXNk
BceOFu6pYO0zjBualbPeWWIzM3H7bObyWbJI/anzGihkV2tR8T2pH9rVuphvoPcgVQs1ILeZUX9C
UCC2V0XznBUciYet3vzNBo2sY/Xeov9tmdTSarpBW109/Y71Hu6srXysqSfqUVbWaMcKuMCz2DF6
R78SKRRrmr06dRuLuPwwvnjcQyuB81LfjTpzWfi3CLWI7hPy/Bb8AMUZ+RmjKYzaCHp8i4V0kFWT
rnqFR1tPlXKmraCC5f34P0OaNcaRAoiF9AEUTyRe5eqCqXID7yZzOQgSnFfeWc4/nsQXQBXrq+oo
qTlq6dDV+/HtRe7xojXJ7cll/9COVXzbEw8d9hGt6iquLVF3L8V8fWVoK+uGo9ryqXAevWetMLFe
uxaNnhjlbN9X/5V/3kC+TEWvx4KXKM9gVPEEzds6kvnMnoPoA4mq64P1DNOcMwoSRH7mgBwkXJDD
SlFJRmHxGUiiQgXDVIM77D6W+qR2IYDA8xAbuNq0Abq8oKa5t3SCYf36iecNhPN4LoBgqbo67p/b
H5WthFKa0XceD41Y3Kq8+rizNdJNV4IJowg7FfubwWjYZIxL7mgdt17VgaNzPudA13PnqNCipBMP
s+bio1fkPkGDJsIKhYStbH40rBmMUMvhkLS1XfltsixTlrbiRJBSwPkIXP2u0Pw09P7l+DjylSF4
M/mP5UUMdCSYBpOi5fgRA7ojFEC8qkj3akYf+e8DSYUu/An/LVmxRLFSlWxBIhnWJuL8OszzKMJC
Ik/71hSObXhmKFHBCqmwjFA08FjEZufE4w5vuCjhQVUTv7eqDycUphO+BWgG75B2uNJ5WvYDBrBY
MbvtrG8hSHSveCqZvbakIcbYZSOBkJ0OCxcJyQpHpFYDP73l1+I7HWD2V5T+KaGx2eTuIabr1fFd
RJTFYhGp06jHG8FGmOyR97K4/vzRo4sSAgla9FfTSYlu2fm4CJiNOsObyWhQaTY8vv+FzXDihUvm
7JlTR7uTlLMeFFt5N6Ifa124XNge9kUPDKZ8NxDKB/hU8g1j9HjdwQqnKEY+TGxyjWXFwVKQne5l
lYnFXHmU4nsOSyHxDdFOz3Xt+7SxK2nZQy4pcRLLN0fAgHPJDv9XZw5wBhbmUUPoCo4sKb+41GLK
z5hPS4kmgmzsOOsGxEb4aqSt4fWNC7L2ztnMo5+D9kjCBwCpOgC6zY/ICSNi7O7arpfS5MRTUHvn
y4G9X1hLWgQ2gYzDycRY3339Z5MlWx1UMvpcoKJoCWa9LGwotzh/O5s437BB5qntlStLYYnyBnWD
/+IUpwurEqNRlSvKd5zSoCMFsmlXUpsfORzf2YLJ+6HzIU65g7MqJEmlLSMwOzePtgydYZ95l6Va
WsyYFZY4VPKyiaRoDoJfzQOTwlOp3T78hLclZwJczQkMu+Jg0hPq6ZtSdYm0TTdH9TJChcJ9gxz/
rKzUO9JVII2vfiUlfESav6AJpmioRullht0F8YVJWAh5buyQmrkMV1DUkI/Lyyui8s8SFleXa6l4
DyWZ82KTEbGX+Bc2GpOrg5ns5r8MOLyKhC4raUz1rC4qOrgqiHHiQAT9xDkF0PpEn3zcewBQjiHz
993irjQFTHYehKL0k05PzMm1lFY/RhYmdaz8Bl2pDOkCXPpfv5rQR4XfeU0vo4W09tLDcXJHwv9N
olgZ3X1we6sSyoinKprpHp2mDhDCwGH+e1ZVahFEcn+xEoA1zNC6AcXTp30f+mKAg20BCH4qmsDy
sT9nisTvLrEnEr3pfIYy5cD5W8Op0eSm/GWdKxcJo0tl+yu9UdHzFQP7yppYrQT0RYlA5L6+MeYK
brNT6MO/ajilWdV4RK/0uPCyB0DoQTZIgjdYX5fsuw8rCLcibd6KJt100u9auuVLUXqF9BHAsSGz
irHRXBMAFKlgsk+sg8Fs7PUzhVB0bPT2gptVfTR5dnKwwTjZPSuJjIea0ADD2NQTrzb1K8YiBVre
+2fesylPaUE7a1sdJ3ph8JgdaNr2UBc3bKzs+lNv9C5J1Jh6Cxy7ltpXIBOgQyEjJL6oHYcfH9PZ
lHQP/oX+Arilz9dhPRqe7xZ2f3NmM/PBqRLDpZXxsd0r1HHDSzGGTz5ChtPJufEeHrgVZj2+9Ji/
L7kRPridcjvd+N+nB3wpHIeuVX+kpRafNU2oupliq1lnIvgzMfUMQDs7BKBbWzzCIQx1vpcKLuqO
H5no0+OKMHd1Pl4jgel+qFwO1oQakB27gfHhjTD4RBXHa2tm1dT3ZgMNMOfQEziEqDCe1lWwJcK5
dTBZc8zK7XyjsilPl53wCYUQC4pubhYp2rrNRYWT7OqzAlxT3HvtPAgtkS/li6sHhL8a8LMrZALM
IemQCDL/NzvomPlsqixY+GOGXFio4eF+mSR3+HCNqSx7RRpsieT/FF+oVN7S1icDyzDhCq+8QdEJ
vDN16aL6TNh2efIGsmQt/y1Gf4kL0VLap5te74bs+u7HowQWlT3zWsQckX19giBa9veJhD/fapLB
upYtliK5bcpFVrlRJcaonoIdh2GLSMk/WYftxYtdkBI/Qip9FOpXRcVAxLdt8yJavgtK+nfiME/6
9A/cqgPEHMdvsuJgwu9RAU8lGU/HCymtzLl300O7sa72hffYx+KLQ+K+pMPif1NZoNbCujwzBN8o
acfjeUMuzA2qdeFLV+2Cr23ABghQdfdPFLct1qPQBMVWnjFybZ/pK/CZKnnBNIqssdnxnq1Q5Q5R
FwJPwWVYw+NSpZ5QjytvjaFC1RqpDE2hh6KvNPJjV53B9AMtieN5UlVYIUHb3h/ngjWFIP0ySnDY
37mFONeQndreqFQZLClnF/YjgBW36D3sg9Yhmg2gCTmT783b8Uke5Z2poM7XyqcnG8iF4y0we7Hn
WiJgCn+/JQEDxNQsGB06acRwQI/BqYtJlK20lMGaTCg0q1dhbolBKQJTK7Pk4ybNW8OHCv5Vs0Wj
5wY5rfkZzy7UA/Y0kkLhi1HYPHDafsCkGT0oBo6mxV4SaeeSPfpTLrzB9fnGza1uzXino1Ix+Idl
AcwHoZL5kvIap4Ue7N2yqQtHx4+b/o7fegt2RpvtHM375cb3OG2gcXX3XlBRakm4SY6H4F8RhLE5
ojyAtpDtuFka8IRZ35Q/n0dJMzPNxPAw0DeqiUdynLgndcXfSmiTu1JonlCc3IOD4hSWveZV/Izj
+07zlUTNnsewwUQXf0PuY6ZKlbZdiIp8gxl+/ybMcQC3AL6nFBeMnyVPG7rD7SHzJpFASCn0K/Z0
56ziKD0Az6+7OOBXfABUI2aHWps9NNiU3qmHflvJn656LmzipnZe2XPIeV8mrob+/VL9j5537H3P
b1snf0GFdHO88WP1EbHCUU5xB44VbKPt0WEHTCCMViqXMyXWtPhnSTy8y8KnpUGOYc15d/Rx80q6
KKdxJkfHnwLc6vUk0F7mDwxdKY5vLyRCtbue/pYU8767dgLw8dg1bGiaworZIHhUfRmZJnWaFPwB
kogugdYXsmdDN7xXQj80y3TcZ9YPZT5HV6mU23spkLHzRAKLA69h7JVwSmChTKU7UV33BnxUv5sc
O2rFbFhgmOnxGw6gJV1dSKWZLQLVX4ptzBhU1O6UiFEmZ3oJojagh80EybMe2IRznRJM8KJreLcb
N123X7FIlXsX7HE51p1D6X+EvcpOVumJwVfGLFIU8a9ugDfDDgitlU0FJHNw97jgRyUUCwSIb0hZ
oyzXaLV4LPg/ReLF+Z83diQTUG5kNF8IHIeT0Xq0TrdOru/WIVp6GKcuZkKBo/NVxF5QtrN/8pd3
eQzYLzKsALKY6V0hUJdLX7hJ/njaSSjk9GldESTZlLtY8jht8+yhQ84QOnGUzcukU2OUk8JVWCFh
v5ujOSbYcm3P/YLpU07F0g1f/OH6/6jGOwhJp8rsYvpq2K47+Ys+Qqi6MClke2X1wejg9vH0sMqo
CkElbPW46rFBVmnFGL4X0kPMmyrB1o4bROQei4t2vBezhjczui14IvKxU8GKuQ7rn+nM9uPYCpMi
hsbs7nU61MqD0n1ajisQ/TWZf4+BcSQMYnhvPIGh3AmzNtMpbe8rtbMm5zthQph9uF2FPczEnnVy
4FbcvwmzghSs79uHWSRvGOWmdfRoShQRxgiot6a6QLOpNqF/rrwJRzFvLkQhrnWL3yBXD2a6R3au
j/9CfDFnlVCpL/906IUobTyOcVeYrqy5QiYwtwMB17Y6ggZZYV/s4HAWHujNZ7lb3Ruy8bHOPrBF
Hn2Pi1qiCVlPZ28AyYKwfP360R4uxb1H2bRrX4y3C8ZHDFRYtVhmtGmnGgifKnt2np7BRWxwmPUQ
H1frpEm0rRG1pYO/9Cv3DSZXqT2SUrK0U6wSl5g6qKMjJ68bd56kIoDydqkVdTozuEz0qmsEhD/x
fABEzlSqAKeggFY2mJUxfNqikn/H1BzrR22y43z/dxlWkQTLYCPvXRGGEimly1uxzbwsZPg0/T9w
Ylhk6gvb7fCgL90a7ubOs2/NUehsvKzrd1PClyYihAMsr0hXbaWfMt7Jq4YQ+Ox7sqDfxBn3myT8
osJm5HIgfAuDPjjOEkYYM+myG6Dg8NF+OwHLz3WtLcE0tI9kPImvWznUbvixCTZFVLZ+/s5C4XA0
E6u7LZUuBSEm3Qt/E9GA9lPun0HqaprIauGs5BzhFIj0FgXTUdT7oqbi8ueeilBY5uobrGdahjPz
RepXDQ8HVy9Lz8me+kaGa6xGw+/KS6Ck5V97JN0xAs5bEqjJ15BmwnO4cFyEOi2w2OmQ/Oqp1lMZ
aKiz5pTYc2EvFI6uTaT8qD7PFSi0VvFWT7oLCE2tO1H9Pjg5K1OQuBWWk66Uj5WcyVMT0y69BR84
Nzn4ZZ+gGkYPblyBlm8HCnyK31QpwyAED3w5//EXs2EIapv7Y7qEpOc9KInizMdn66iVonRKDcOA
+m9mhA1FCU+IXGS6pk9sOfkqNheSMO5xhEVC2leHacww9LhIo1KnpGt+OnfRucAbn4PeZLI51PbY
y3nV0/ec2cgJXWb4Y/Y5VtHrpSddP1Jv6/FdwraoE8gKlu8RLhMYDvWy86+95UptE42T/Df93hro
48wK5kD/ti+vPZt5CdhsBA5Utv/vGcKYhkmmuOHLsmtvnPkViyCVel3YA+nqC+q2d7/6PZxmnzAN
BsmLp6PjNY0xN1MeqC8pjGITGh+lGW3YofEMEhwgJkhkNI3wJ6HUqPklzhzmEwyc+aMa6MzleMZ3
fXEnRyR87aGcsDUMZMJz8od1wvgqwiEIwtXYMVpYFhIsW+bF2ujkwU5uB9O0d9JEbFa0gRrQ0o/2
OMXnCp0Kke1eyDtVYLSI3R5ZtQDa+7Oe4GD89jP09jHtsXBRJBhOJICT9R2Z+/OiNpF9YmqsLsHi
XQLBVQcqUfko/3bX4lbszUdIn5ENZCOj4bWCKdRyKInrMw14q8iY8miNLnVW0cNs2d6L9O+vGn2+
xkJNFDstII8ZoJZT7i0fz/gZjuOM2XdsGA06rLJdK6qoOzf27oxprIfx1jp0iybnuf+n0vKxUwUq
4d61u8EY4YYBKNq+SldkEoDqtfq0+Jt/HpsG7zeTzIj+nEhkY0LIcUy4eSxL7kgH6H20upoanCbJ
4nOYSB7riQZNzUXlC1DR+hS3NSTW1ZjtDLuB1LF9pmzZjkZsRS6aRn8jqc/AbLhHBmKTQzN52ycD
8NxTm8TvX9NlT4hMP32nltQg6dHc6F1X17HTztCCPqjyBhLnJK7nLrl669bmrGG5oHAnsLFUcODI
XI/nyMa1fLmyG84uh52i7KeupbzUygMTmuKFUJblZI+cit3WC1mK2wqAprRzG+r52WSW2u4rc2BA
TZ4Rcc9TAb4vJizdF/+t9qYANnKW9sFa+awtsJh8Nyik4MAZXQZAuOozpObqcdGTh9K24tWJ09Yr
gQUK6fgTEfjkSamFMgIv/Dr0YT5hXN6EHwl7qOfLDnMAhTV2gxoI+SxnR/2meUnSapSE7ido5rL/
5EMSCyXcsXhnXxUMo5kECfoczl13ZY198AlEL7irkrVZ1VDFktMm0jsXxMr3TMEO+Vco3BBPoLCk
HmL4fcXpkOYplO9tg+AQOYRdjIGbPoBAUr4j2kcgcfGiI46UpSfOsjlKvKXCGIuCVRbGvTdbehN8
xnfzr8VNyhBjUrvi3X0JKp6GvG65VdzURmdnKC1G/bUtiDaPix/Pi9ZomzbyUj92Bj7nlkTja2uq
nIHT+f78tXLa5eWgtFir+mGn4qsCFmdHTQyCzlCJ3TR4r4BmcQWoNZH5mnERBgGUBEKPwhtubA6k
zbBWLxoZAwCPaNN1KPkBiXb3e7Jid8cO8B3OX3MKNPx3KK167pFhc+TFMCqMFlLLJtJ/ukvUojmu
X13OIram2FJ+3mW23kLNkT1AccNGe72jhsN1+1OpV8bcZhmMTITd1Whmn9Xa1hUWNgjLsYnX4DKs
ZM2qp7w/Mz6Pj4XcmSZ3/v2UG0kV3/JiN2Php9g3sTEkpy/QyonjlMfX+rB9U8ie+9DJCqmU30xI
HVtiBwqlO4umIjimFQBkl1lnZ9va7SwsRgLkyuUnsnjnukSxarA0jCQbL/0hhcDZbrX3n6Q3+Qws
ElyECg0dml2eBbKjODe7m1XZlcxG62sRU/QyrDEGWHtMdwjLfb+m761Si3NPm3WljALbXxKCTQnI
HT7gbJ4C8QKJqCtmtBSZ3u17RcI8PPlm9p1GKvAq2WLwdsCQ6st+s583k2q6oDt3MYtqL7Ra2UmM
UcpR4AujrpbWXOaOSw6vqVPgZHz4jA20GpY7fI7LjeGjdNyiXiu/blRzKGmlhPtsHm09z19FEkHW
FF6te7euY31zi/IIvzqy3KTPXwfRc1W5gimrAFVOvJxuRr92QFFSLSl2myb8DFlGUMK3UwgZcwSS
ghP3mX94GyFywiHqnuMctByHUtAyjVMXPAUhO71lDD9wy0vA5fEFqK6qq0V+xvnaeHF1qaJZihlb
l6uIZTY/N/N5My44u5/TsH4qd9CivHsDgSjurBDToJqaSfLw67BvToHj4Q8YCw+xJNND6IFKk5A8
WYFa+BMwGVdOV9NdVEj67zN0byDtSZcrM1+/y5T6bL0/K+MSo/+B9SF0UKpLVQBQksu/l8Z8DOVy
k6uRp2F/ZcD3paSf7NkR1VmL0D1Z3mE7pW858+jw/TYYAm55R1e3Ib5g93KDgjmryT0kCpJJBJaq
WAz/c2Rjw2RPW/NEDRc30S1XH1ap787q8cMyu8t6aBUS6QAsT+LCQnlrK25rJN80y0QvUCqziLIE
RRFkmHMgyqyeJprBvVSHEAPXwww0kcv+JqKGaNOLJD25B7kAeZ34zHqBp+nBAtV5pB2OeOb9HeL5
o7DgffekQHmwHDx5f4z9Oh8yHIODXUSYwPZzIk4kaC2xV6sSistx6V0U/KI76/R76qW1jnSjoYLD
oaT6QSeWEERAnorpjCyBPCJg20oxEjpf0pDrvFyehFvEf47unx7IO9rlyNRjoQgaBevrtmOw0ILj
7g/iVhuBQsPDFw1cbCekRmA94dlSbM+qYYPutf2rQU/RdUjCDKmPvlTE2R21GuZ7uZfw/jN+sNHT
jDA8ASL89DkWuSZgnUDDsTQ+c5XeMxbsw3gnjRd93/meEmSWBWsyfVlKFUXXTjUtpMAArDTntY5V
E21wOdRjfC9MOLGGnTTvupU1+dxeVabhYERGwevdeji7fPK9RLvDglJGBVPK37xW8KYLfMJG9twU
opt0wY0A5wkOG2yD0MZKrWhwOvy8hD20+9y7IrjgE6aYbaBTE5O6DwI2dDddWhGuIgoT6xuREycF
EdZECLDqkk7SgqI5lueQYL6VCKdFtmKuIy+H9S8+9NXdehM62QuPq8u4lb8w8dIMWVDcSy1B5Tvv
ntyOIoy08waDKvwHox4y7lNfIXqsNSnmSRPpHBRpiITFk//fR+juYSq88Icp9IrNeVkELY42c9Gl
ZlYVcCtyqlV76Z1XlFCz7TZqTB4pjY5PPz1Rbbtjg6TCh60c9Ne73QU776w0bf+9mN8/XMyC2Dks
ZSmfPfGT3c10OvzlAZ/T9Q10Fr487HuNm+cXQQZ0sGR0MaB3SMHv/IRHOwjbh04YOljU5p403jn0
9FPsrWDwgtwdh3+6PdrAJzxj46yshuJaFHjZ0jWN77Hr3pec3vjSsAzq/2Zqv0jLuHcPh+Qa3jwk
O1FnL5eq5WYYSYz9YwoM3kDREKsnNiF1WoQYQwDd4flX24SJYqKNQnsp1uk/mFWGKb3gtIaXb1R0
imoC33oFCBAHBJ4ttQlUlMnnuxGkptA7/0aQaEZILjqaxY1DYbkhIetD+Dd4GOuFhZCakFEjh2q2
hbPezgUqjIRSjSwMdh1H20wRKdAuItfEr1jwZdB+7UDQXsHpdM1PZbQuOU01apD/6kwCKB6UDSnS
a/GwKM8+w4BXT7EqU+5rd9o89BM/rlfKgri+ORz3aajnhSEw8py3R8bccTFz9mllJxoOEJAAaGgA
zfZIZzl6tzzrW/A257nPvLKohAZ/Cvy8TK0NtffeoKJjrk9tkW6r1C5BlKNlyYvcOtww2jqEG7d1
lbruqElDQx58hNfTztt8ZNCCBqn+kNXJJU+7QncaOrYqhgSxEKkwkSSbbyAb/zcPhbRcGjVxuEqa
RKGXgfYjVfYry6lXvelZ+r98k33rj/WkMCLjDFY4QSDfrwxlXjCSCiviPUkHuZK/lbeAYySE3VDm
qs7avhnWG4UgpSIIUJ9gbDWX3FOMbTTTYhWhwr9XEzU+Fs02qPRjkIER8CX0nv29ZgvTGqvyvLFW
HxnViWAnDC1We/OJRhw/hsCZFLuG2QbFHpbuKgreuPMz1FXumZF3A+uUno1Q7qWU6dD19Qtcfu8z
Bj9vSPwE2WqHCDhd9aCjf+L2zW//uB1OVkSfkSL6hQOsRLBdbCW8+MU+taIbEIEf/s5y9x3yAJkq
ym+rgCPuXzzmNUXg2qRhB1n67i7n4PjxoCaxvDFVtZG9UJfNam3OWzJJZVLCZPSvpXUDVNzXh12J
iyitZrdyP5QenPIcsMIoF43Q8BHnGoNGpGPQ8coNJmDwpRlUhfINW3bDS+jiho5kE3+3HavWJ15f
c7w4ndB+VWNAZv2D6PImuCDMiZpd1qQjkrqSGKoeiLeT1kbiB/aXe8tKP9FjblDVx3L6h16jEg/f
g1jXlHFPbsadJqjrqU1UhFscOq88LQSi9KRi+0I/b1/jpR3QWHaicXt5t5xb2r3fIwIkYT6rvZqw
IYIDWwo2d8Ef20liPzaa2wz1pLiVs+ckvdfYcdyruFuUeTrLcVBkAYIZzxtDJYniUkIQ6X7r95dJ
5MLWPxZIL7y6tfTMHdGeYYRxXIlGksMaGvxxEJh9/rqClrjz483O2OUzI8L3WtzesaLEhlQGBgKH
ZCYxu+0unfOKgxRRjwxTK0vGUQbhbPWrC41BU6e3B6LfNFrZAUvdi+0+vqagWkVOoh5sV1qwEQo/
FavCIQpGfLt70XjZOie9Bsvu0OGPNl9FeDkLjTcaWR8nsEvEvkf/vmIPoZ+FXqjbHYdzH7mysHDx
JNm88gE02eUlEPBBKxL4SHRUi8OdzdkdMrJ0haxg5rIwihtX1wsvDk30p03YI0ItFa4PqQcflYV0
T1QcHKp7B2KC61MuM9tyCUZt/fIZOuCUCQ5mk+4WOiKg4MM9SHDtEK2YBhnEu6dkLJpfwHgatwQC
T8Stus+ExZvQjWJhfiY3jlDnSRXxvJpuzBTT+q8Ed95fTTRYAXUl1M3ys3XEPGTkupcWCgRiQZZF
y9ldsNGqlN5MrqraUi37fcP0ozzmla09eL5ltHh9eMmusexYvDVSElrOdrSmFvkONi8ubeOHM9O0
Ac7ZWbdG4LJg8Pqz3oQTxnsPgY2w+9u8ofbBgTxjvmwVkrIQt2aJJletzsTlIBfDrBvreuqexoFJ
GIUyR7rMcvCaRYsx89l0Md58+W7+knxbWh1oh0a/SgZ9PGk74VAJL0phNF8OAAtbSc67yoplwLHH
Tm/Vv26HFtiiTcb4xoXjSbBm5IRH8rmjA1Gw0QhhDB3WZBCXF++N031kDlm+tzlNnyFLS6agBW0x
bpOoQnK/hF2vS6Uw2NkCSwozD1rBVoYLhr8+pb+7STRTB8Lf1K05ZDtJ7USNFOK9oeDhbpXC+Yba
B1hwjogG9wg2lojweJAbQqyJXHjTz5XGNLruRNMYR11t3fwkzULG/bU7tzf70Lt0CtYEBkh/SoVJ
10GHRv5xoIqNS6vwtAUpk5rgrwRPK4b8O1QiNrQaI1s/wwJL8Oum7mJa5RZaBoiXHVqgMslHasL8
DEFUpndEYfrhDh8ueMXXYYmx6hDJbeuu3Azqq2CQKNpR3qNwP9hmN7CoZNb0EalsV7k7957MgGYb
0qfKc5G0SaHsySXhVefdX8UZU0qi0UPv6igRx/tdVjfNl1xop1TbeubwE/GoSHSCaeZsSj7Vo/H+
MROtGzfP24u8s3wndeLwdih2cCIwkt0oNdfSki4RXN/oRgf8QN6FCC9NjqwPix1RABH/dIrnK4Sl
9DtR6ckkSxXWc73H0ohYY9Y3hsxvQbWerwaMvoQYO11Bnz2uUUnZQIuHwNaThZqpko4YNOOwfoiS
yhWBBkcVgk1YDs23LxPGyKppT50P97U9GpjOZS7ChUDLcbpXyb4es2jI3myxBO5lvMz5U4bdYzpo
JwIOP+ibwqg3+cOEd20xmM/WGam/DJi4zbfqxcHE5n6LMc3U7tXscNZHPG0SYhg3MSW1+SxQqT5S
LQtyIf7pGN5MJLkMRNgUG1VXuEh/6r3SSRqhMqWlc1ko279e94n1OqH8dmbM4Rijkdv+ejFWVKEw
5PhlXXZFTYDdzXXblBJ30IRAZBV3SMqiBgmmG24387UQezwi0M86mhvtLtG7KykLE3JHDakP6Vx3
FT4rVc63NvAmqCNcm3B4aIcavd7D32DdlpFiuDjBysqB3jUHqr63CaxaouRCMh5lSMoiZK9zu9iV
Pz0ED1a/wAAOW5fnOOWlZu0hjxFQIqfQtGsvlBxlYQbQH9FQZFMUE53emOwnHStt7XEk+bsMaLDl
0gPVFRka5SHCBB2IP+gPoYS7ZM/hUSU0zj2iI06nl1Bb/exam69CCczJH+zK3uy3Z/ISvLkbCdqs
MHZThiSFuJpMcFMptEmAoQw24R/xMKbXaAZP2Sm3bXf7jUXxmq3dBo9MP9XMvOdyio5HFPz82CpD
SJGMNjdmWGE+KdyEA3z54PCl9FrEDf38/rnxPjwcbkxjwc9l41gQsn9avXtSZMAJJejjoXDOAUti
zx645/JbOBt/hbzLKU4isocqCODrQcbsMTdaJhvFdILTWC78Pk0H+2jg2PxFoapwTa2rPYa0sqO6
8OXnTjCsp2aNa3w+8DQ0C7TcBs5E/+IgTR3HN1VzOleMZdU2Awz6CgiEzlN+Fssu1jJqPiWbfFCS
pcU6JXUNd4UveI9NLprc4csmHo7a//+TiAjzCGu66FL/4qheznwMbQ1KytjF2MJddVHnLf1vkmCO
st23P6Qxv9MZKuMwxBhc/ZBt0ZP5s3qgbNpdm8+03ZId/r428b1QKtL+7GWvMumVTi25l2LjhSG2
pYVKX4xlpOOhsD7ecGWEKP6yYqt2IjWQbPPCbxMKnjiEXpusiUdoCdpWgFMjWLReNeBZbbmLamPv
G8WzXtLmLvdc+CAozkyIvJKpe+9oaVoDYY9vjMBs40OyWKpD8LOdyuVNCUgT0bA6V9EadJHEcwp5
yssZzHqzE4jhIk9e8aa5txpd+E5PykOePC8WVY2ktNiVNBPxBDD+ykzi08Md3OAGWaPfu5Qs9Z0r
etDs0zwwERPSC8tARnxQ3Y4R5CI6C1NDFTZAKeLeA/44cNNdX86qISqNDuBtuP+WKDzl9gDRVdSV
oMBP7FghUrFXam0FaO8Wb/iGoaH2jDSc69S0qk0J339RcJwn6NqSfmxVAKNoLd+liszOe9IYIckT
ac7M/vLojyLAlVF6j73Za7NhlWJGH1xBIYeYp/8iPJu0+hdjjT6UOnp1r2PkvIoPC+RQE8vdEcVq
ovPLyu9MaGYtUWg1gHe9yxpY4oVNCSPAueKsaDVV61O48rZjPQAzUEAWO7QrkgRFItMdeydqEfXb
fHUGXhi0vqEpDrKi/07PURun6vIIFxQ92vLpfLJTDqCq0b0GOGfWJHGiR30HYzBpwMhgxMT6NNU7
T4O5TnsMxqu+OC0wjEj78uIvJYjUf11umwJdSVKEgoh4O1++GPnBeHDMwAg4aQqNyfH6ckS6MJpj
xFdYgWvVhmoNRrp+mAxJ2JnnOBubLsRh/uyouhsVgK+7zKUojLxjLl2Gj4pibUQHcf11JTktze5a
OgqJt8nFNIOQ/dIv7nIh9cihSohFwb8bBSLFv0r8Vz0pWe55qTRxJBYiYUWKzm6KL4KiMhvnpGsh
NlWDr0XErknBe64T0hFYRx5jtEMFoBE4vFzdIclUcNx8sh9KZnYJIfMMD46iQlJF3CbcUZ+nVPf6
UM0zUqjn8xkLxuoYZ7hKwPkDzBErujr7MkmxKEGNUcwUA+EyFmxrB6JjKDJn08pn1lfDxSpK4IFs
yNQytViXFvlXDDp0nTplkYuc8NeA6EsOBrcr0KSg07a2H/npIJuqHdG6g+buGg5NfNAh9kACp/cL
CyG9tl4CBtVt+fSbRyOlwL6wNIB22/oDgPTRcS9SaXYDbbvlAE+lMAC9ad1Vu0cfxz0M6gWAko20
3wUpBsM3nNRS2mNHMcQpHAa/OWSPEAh2uEiqRDlnKWhouvFK9J8jkhPjrNkmXmrh6rZYF0WuZSCn
R/yfuuEEvCN8Njz1BCpbweirjrwd0Zrjspr/3WAZ+JRNv8cnOUPrkcImeX0VkE5zk8Jnubt15pj2
sj3bjvtCS0gDb7b2fL2rBv/+MM24x+5t93lEaCOxBSJ5mQ5qKJJ3+l2Ez39NPd1/C0uEs3Vedsoi
5cl0FJCm17ibi64Ji+nXE1Wms4lQ89nDdOlGPmn823tdtEppK6ACLVz+wp/kJvx4v6UDsv66m8/y
xGj68S9wp+HGBVpwd20XeP95aA9MGxcQR3ApLFcbYxu+IPKsaVowPQIGDk3TTGQ0xbCCFHDXx8V7
5UxX1MlTB3Xp/tL5XIBXyPMGfTJkOKXSDUA+yvWbk7MxKuaOHXznaH4Ht+Q+eFBTFQls1bBH/pmR
pwUq9n7FMyQ04D0vxGutD+CclQynfXj9GeTw/R7hP/FvHa0vw1rnNdF5UK5Rvb11R93ppKi4NtIU
yZNHPMWHWiU7MkQfUdhKgHb0O8Ub0XOdcIlWxvuyEOOLOd9ojF/C24G9q329YLc1xlVh2x4y1LHH
ptx1GDXUivJmK7hnWF07UsenujK4gW4kJjV/rC7ibn+PH5ap8PKSOeyZzS6CExyBk7nb4OniQfq7
7xroxfhr0T0M7sFeWKQudCrkv1XcyQYL+Ex91POEURoZTl/IgOY45Fvdb98QAu/MGub3Qa0ELGza
NX7n9/hOV7PNLsWkTEnB2eyK/e5MOA0LI5MQZnrZEx0maZgxf3a9R0jjELw81yv/GxHb2Kil3/mu
dLkOCL4vwmCjpUMLYeGaXLgM5XP6LAWmZFlPo7y0M5BpxJJ15lIpgdUOocZb6M4ql25ndkSAkEaC
0sVv3p2UihkLbF059fLxju1l9lVixSApvMO9qBS0w0TaaQnWW7xac4SUwC/3duDn1B83mGmg5vSe
8JfK3y26m9lgO3NvDwzWFYVUcijjyqeJtKNOUnPlojHenyyxq+Qf1kyIfCZO4XPErHXw5vR7NLLJ
cMAbZHyOb8ta+wpCGa0BhBrAlVCY4atqkg2y75NtxTxVGFM5Q6XuVre4c8OOLYTWRpDMzHmEYPZo
GxN07g7sIIL06FyhMqZG/IFEFxRfukz07c2y5kPLSRnuEIVXBuyxh+W9cxTzav/THRz/3KeewcJt
9YtsAQLkTlwHWFQMZjWgu2I1fOUjZsEHGVxplS7Z4alJjrp5ExQJShzZ8UdDZGtclwCuU8A8Zogj
bzc1czOr2WOKW8L3AJ1Kc1OEf/fqjTuckKxNYVqN8/SwhbEG74KISIRfNDX83WSa1TmV3dJ56oBs
aSGGA4AjR3i0ew6aSeYuSBb6fco5JfWHNc27+M+lJqX8n0v7alIBYO4INkmykrQ/iuk+VWKqCbqm
0+DyyIncyyFJyNTalbU68MTvd3/h2vx5C22okaMXM/Ai6TTURd2rDBIpCRpo+LkfsGdPnMm+z8sZ
BnhXuxk6BeIyfhfaPfcVUTLy9xiLSud8TPMvTvUWzAyRqkuVnSGSCIbHVHNIZ1v/ydrY8FVsh9F3
Xw8kZWofC19rCRLw7NfMwLLITrK9NylW4w4Dh5lrt7a3e9q7jjzlE1cBeIrBZmP+Ib5MEutjow8n
v5pPZgghDWPSPV/JjQCjhjNElYf/Sa6+4XgfbqU6ICYpDs+6vWOQG1cwdz2FxXYb41cQxWYoSE/R
k9NloUhCwLUMP1wxaIfibv0JfBGQ5PSFCGNEcHQKy9r/UQqnGxItZ89drWUEnF2hREWcf+vF54UX
kIOnnCPvBHuZaqI3YDjrMpe26Bej4/sQYz+QUoZgRM8TVDDnzyRXZPFgvvVbo9p7TvRb3Rc3ZF+u
8j0f8bABlTNiR3v6HgGE3ewydh+OzpAsRyiAQ4e7XCd1DdieVO+ZGtcMgz14iH91lmBfdfxG+h1S
ukevRr8i7ASyD173Stjzak7QnwuFeb2BrTzPop8Q+gInD5wZaZOQMP3rNARN2xbSFZFU83bi5t2L
BLoBzbJZoviJc3WlMBp1b6K57eVCPft8c3uOTx11LiF4pwgFjGoKxLCDpB9ETFZ4zlCbkuunRIrY
zx7rd0sNQaiy5Qy/ZzMV5SxkctxWk8AYV9iNCc5qUiSZw8S56qe/7wbdFR1fZkfmV6ORsXJbbxSh
l3lE73khjS3wwL4tQLeuq9XtoXKRGOVsQK1M3sayJWUtwhcJHpdx9RpzZ5UPH/SvHpHXLffZe4Ah
/7A4RvdL1+WtRFH0NL2LWI0uN/gLcWEyp54ApR2W1mnHddPIAlrXuqFrCgQDOf5vINcGY7IAeSgE
J9UOtvb9U6OM/QgbSTXDhDersbCd1f+jTWhmlstmm7k90thZB1V2l/bzQmuQlkslKaeo8zAOOFLs
DGxQi+KHROEBoc6f3bIb5HSsWnc20CEHwxrikynV/xfzgbw9PiFTuMNMSBmuFKB3SsucduUKHM2A
GSGXQ9hH3cZggpqrSopaaF5jIDc1scFipINo1nVBb9i1GwI39vXk1zX+M2XKwppHvKJKiVvJ8FbP
jHDurARXmdEPlW5LibysgEwza3ICkQz7cTHj7Zrb9Gjnq7YaUM0qN9vXCfKsNayRC52exjF73REz
aBeyDT8bhG31i7HmzVgbc53o+IyHMFIkvdG4SXwWAZpWnHxMa90RHGhd6W+c9dBQUmlaAY1j4O9q
5MJZEr4e+cd5IdEvxN3BAtP9KQS2RHM7R2X7Z/4ovu8ZupvV3xykzz0wfxsaiS0vjh6O8iUtQpLk
Vqf3IT+PdBPBFDX7CwOipI222FW2TToJyFLcBKZgjI0SvxweWTgxYxT8Z9uJcF6T5iSTVgxuUnuL
xfOaAzyvjUv/YzXmVH56Mi9mUxgKpl8YlWZvdFTeOPhzj61zixxraTmcmytb21OocPoXCxMtqETm
fsRSvrc9pAIl3dlKJh1eQVi2c1YH9jyzVRTu3YxRP1GHgG8NoF18zNUJFvOVKisN7DbO0MFxBPwc
gdkfhmzjK/HaImeov7L3fGqH0PN9txVlFpdX4QurL1URrcbwBLNRolHFmiXDV18kEGGptB1lR19A
31NyX7vNmMvV/LS4+j2LM+RfkuespA5B+8Zk9/FbYJ3uOpqc8799VeKeADCXxvtBAOhqFM9i0mo8
dSWLgijmf1DdO2hnAQaLBOx8B+Gu69g5W5fJz61GjHLBJm+dpT9KTgnf7yn+TKijtN5mDMA0J/TM
Hg1MSwW5rSKFCGT+6riiDkm84DyY21/cUwOeCGQLbacTXq7fZdzCZVpFsJV287dPd2Po2H9qs4BP
W5crz/cxqydVVBKn68QoKZkI56HxHHXBpK4SEt80gVvAPtz2wKmNUQk4TDQO9+xiJmNxtQYe19Dg
usHKA6fiN8+U2yTBiHC+7d8ZrQOY4HD1KuXU9wp6gb1CEWkraFWEQuOCnOPVjoKVoz1cMbRbu2Ul
hlS4XdxPT0zS3sgT8w4F1lWIs/U32Nu8NsNuCGidnJ7EOsI/O0KX9gIqawZV5CysSBqUKLa32I1d
gC6PSuzOTKwLInpciPlC/ws05Fo/hNuSCCG4q4yaLBpL4PRiDqLNe0WGd2GyGr2fz+ne3QuRqrNZ
DgmcDr88DpsuObP5pEuDiCdD/WvYcwmBrooA7RC0q/wfOYWuAE7CC4bpukSfrBjYrCbu7oczMdPD
sOFoNg7NIBZKUXM/Eed9BrU+Yot8nUJzy1XYDrBXIKGruX0qFcNopB4bVn+/LCU6lvZWv0biLemo
R3Or6FfojLX74F3egeus8NrEx9tmO9Zap3B9jqkY7+RXR3HOhwEhY3+zFUSc9GV1oHxCgt6yUzPW
r0YRWOl9Hh3NPwocNejyqS08TaIBNfjcGSHokvEqKIDlN5tHRPpwvBOa6DIzC9LiRj3C1Y/Jam+H
jIBtuhx3BDo63GZQhW/Ud5CQXrAcWSb+tD64UVWA1Xkqp4y4YSghSQdQhvRLwrENJhQFx9Y3svnX
oXYHoD8t5oV8ZGUStCOq/BVAE64V24rLhZ7ivChnaso8Uga6XTlhH0cuclvdx3CcyaZTP1imsB50
uYTVwxwBnK+boHOas/oI6wYkaXybjIiFkMQ6359F1lM6ZzI0to04H7BLtxo+Y8hfp3/eMDEMLGNt
f8MLB5kPZGofj3u/P7PtSl+K6Qa4mTjzirxPq0aV550JN9kxySrbWdxqMZbsNggLlCCFGSOxzqkI
aunYgUvUlvHd6uf6qE6u5jZiUu0pDTttg6Itu0qqC2WrZpaNomZMAS87eZllAFz8IY+aJiZW63Bw
DI+iijyV1Yo5sxRQiQlWiGICQ5f8OFWRttiEcUTufrG+j3OvXjkI9MqfmQKTywamrspvD/uxnPe/
z2RsyTNcJsquM/dEswXBM/AJsHF9j4zywduWfgt5+dTK5hgDnWOvVAnLli0mkbnUvlOJJeCULiS6
UsTh+cMr9STxaWlQSxAgsbuM8qDVVPKuUE4B+ChBtdP0KOR0lzHfXzTAUqWAK8S5iKtPAHmmS9P1
QBk8T9WzJ7VFyxeb0JrBV9zaotnFH6uG0GkeWprQhT11Pyg42nFdNLGG+/E7Jvn4wcctvF79XsCk
PzMlhmeRW8qhjayZpG6Gxp6KtzPMIJ0KOIVD7LdGlk6Rj6Xe1Tf6/ounyToIBY6HQOfECytdfXjk
JX2revZOW2k3LP755gG1f82v8rwN8yd2b0zo+OM6BgDnH6c0YTCpY1yh5kXTFM8rK6iUVZ5OPqZI
Xs37S2NUx97n2Qv/VEN2/dz9ZejqXeJBlJIyNa8HIydfi47FiLRF06EDy1O/spEWTx9TRer6oOI4
XesFb1Z+pXmjFj4FGCVnie881dF1DVahPr1W2ZU3F/8QSRiIcqB3qDQiJxsAP4jq7gmdhbyo3TFk
KY7MKA+r1asv4p3QL4yQ+EqJZ/9iucQpt7femOk1oTOMjtfsNdMdxU7KVS+6RfntIcKFkQ1XRifl
M7cP7RiqwXk38TEpYKYlaTAqPDwo+UB0mfAaCjGdAGcY9XDWCIBxCpWElnPqljYgMkTlyPAsQ3jt
Rx3eNn8Kfq2KMAQMp+eNCrQg/SiRwdV9ZyJY2VUYqCZ3iCFiJF2+alVdbN0EF+Ve7Dq29H/LkVsI
XIvirmivfDNfXI2DN1QEJ+7Jlb48Lq4sH3Am76MHqQHlb/WVKBRoNtbBSmDXGHyF/jD9mGG6fJGU
n66/tR8xxjVyikPGq1rGfdOUheinnQ7DwntKUe4IKqvdkt+UH7fVqi1jt2zK5jCJS8g7l2hmHqdG
jmzPFsTHnPlpdT9hMxSCshFhNvNOAJCsMuTNj/FsK1MvihtRPdkSBXaU3Fbv8rooU7kQGsspObfL
U/SVwxJQl18nbwWqgyg4W/AVKindldlHUvLBjm9xkXIY/Xo5LW5dJyyV46JsaIHsI4eMENDW0Jxp
nx6uQOHRzt03GT04z3iRwBv0NL6RCiEVw0G5BeFr8Tspm0XsvV5NzQVboUXXC+1pT5KM7xciokkI
gbZahaDv1gsITOB6QKDgQKdh67UNsnuZC2kPf/rKhqBHPyIxL6rppN8onzkBV8qi994WDvFmWtTw
0DNKxiUXY1kJMnJvGzYEfWwELScAafXYnqHusIuFYv/gBvnYrS7YtjaTNDWY7by/3hUW22LfiN7+
jjLpMM6UtfWydRcuKalHReq0i7Joxv/7G3sxkH7AhbuTlqPFUUYGTOvckdru3sac7drS45Iuq1AG
G61/RFX57g1RfF/mAus6TtNSsEEKCo3xqezAPHQ1Y7S6/POQ9f8Ym8GrjOxMEUKI1CC3lyzKMRhP
DE7RIY9FlY6/GR4QWDfm4vFeCoBQd82791u3grJ6l1I+W7A9rMVUeDzhPZ//6HMPcJxJ9uOdeoyr
NTOEmMh0nCwXuTP+kXYE4HZ1g9DEnrA5u+oX2tFMIr8uiYSLH5tV9j75gEXOCZv0vZ2lgOjeV6PH
4AcIjxvyhufWrq1RGINRwXiV0tnjfJz/rTbW8ylj1E0BPelw7iK/WxbbqIIGhGWaRdwJQjpQ4xoo
4+IG1e+J6jYGujhhJReRQIuHtGO5AwGUV86/Cephosc7KVzqBfIzaHUK1/RkwDKsJbJhEB5po6w2
r7vuk5xjPyS5uAsPGZTsuDD9q8qHOoXSnUAN0NmVA955r3CqU/wr7RcF006CFMaIH0eZKMUnkfx5
8HmFAjdqf5xcf+NIIO9jznqhAce+YTIjlJzJmk1oveYkfi90bn4eZ6pWqonZ0zKKd/xFJ7Gm3/GF
3DguJ4Sg35/xUCXuPaceOu8wOLloXsbfJIJdKr8BLgRBRjf9vrY7D2nMayCV3tIJEmR4/sorgpxC
9rTZS2FG++Hmd6o3RGUvzT2SUj6LIPfPz8wQsi2Y5ZNXOmlYg2+y85ShyCBQDR4XYrGqPJ7AZWqY
sCqShhXh+5MQOZgeGsEWKn8IO6c6TV1M7I2cprtVtsznrLGit/2gkhYDIcepiTr7LrEhGZVNRupU
nHcN3BLHBJtRngsSc3AT6JvMyZqU/Cy+zaIHo8ms9c5Vc/4W7zjgQs6ZOm+ONZRNgZYfT+GiFE7x
xCRf+bF4tI5D8fCoHxwgaTFtWQAlhUeMJRrzL8n1Yx2x2Qgo50rdm5cVEzr15fc5sxI4c77rvKpq
t7eW++yOCNikj04UUEMrwBs5SyhYmTDVfnzqOjhugNEhC5SL3GnroW5Xzb3AsB6feBHvUjOzg8hm
5o7CO8a3nw+Kl3quhbDgvETlDdiFl5WU2LmV6ysSfMOAGBI250f4jo1zahvfPBxI1QHSuyxDLzDs
aLCTuHVkQkRWnzm/gqfujHc1nlv6gn5E6PcegMc0ncI/PRViUIFQuhBvmRek0jx3pOQT6RWWPBUT
rpH9I3z4G29AJFW36EEkdcqpd0ESmu+w9anEp2kMYWkblLQ85DlK+j6bUYpHUx/Uk9Z16v04NGd7
SqwVbIxcadA7KvP9Wxl6hbKsS+/cVasnhhuCK299RBqMtI9UYAA4fZOfCt4YbsLz0UqC4KB83Bu/
AFl4Ob6na2p9vVm0quA+aoRrdN3iZsb65Rni+xZuy133VucsR8Iyx5s5BdEv2CnLf8X/vxw9e+uP
2EHlPjV9Y/Vnpa/+vZLGWFpLoLFFRUHcZEJGB96B4j9ihVSqSRCKZcg2jiKGMlqFvqPPe2N7RBf6
6xw6Unsja1eIiedoBUo+9j7ihxvUTSiDJMJlEkJkSj59vnHOGJjkjlJlBNQc3Qxn4jH+RPLWaIPE
9CEwWW/jKHXCQX85p6Oc9xJlNh7iBzzEr/6P+wxZjF2Lvc3dp49LTi+cPzID0WIYKYEB3heY0oza
wBI0pIwXWAgsp63K9DRF5WCh7+Fy1EluQcOpV37Jqh1gi5vvfotadWU+ut86uReThw88fwHZEQvP
NdY+zd2wxyZsV6K02oeoAPoV36ZsXjGVElNPvRnD4OLxU2/XqoSrmEAtJxxBN4rdzsPh80JmuDhh
DqzHevrihWWkCbbiFQpavLFmTLoHKq8mjGzqzo9QFywx2WgQduQANqEygLZn2BNfjgAM0po+taMW
wX6WbOwi4HAduFQnOY7U4pSyRRzo0UgFtQTHQGvyHdxi1T2FZ8VglM386HkF4/ubfOqO5P+/Y6mY
5D4mfs0PjkbfiV8aOmTaRo5sR04Scd2xk+9deQzqrc78Lgis0w/ya2XrH9w5vwH9b9jVUPpeya9n
DJU5aa9gbuMNG6nFqn1jK4O9nJc99iiiHKsPAt/M/xnIdsC6PYzyRaWqtA6Gq6EJHZN8kFriYsbQ
HlxgxI5oAFnJr83SThXBlq3oqNVnVo6frw6ui9KzZC5Cx71rOpEq+LeQ/NkWJncZkfpXP4Y2Jgoh
TGb9hi/cUUXTYT+xHo2X2dccUE0lb2/ZtBgJW+nB+KeIcjeb4SNUbTWwbU/bS/Sn5+cvRmGYMT7f
w1sltSzTi6pHXyZnCoH5GrNjq8Bj2NA7NtIWB4fIaXZ5a2msORNp2dvVmR4AanxR+gr1/Mph70qS
llmwPuFvKmVbv7Q31uNy2qShdTiG1ULW3DDi1twlnFcL4j18HAFqd0rsf8SWX5eTFXx1WXd/k1n6
4CJBYd09KO49DJWItv7jHoMoo0Tdq5J6IU+Nxkawl0yrEVMSjjdtbYfN7hVAGjWeZFbAPzY6NRRa
D3FWPFT7Q0ivcKoebdGZ3P3py5BhvI5a5MOZ2GEDZcWwlsR/adqW699LitNsx6JzLfA5fPCzHanq
lAwFVAaC2unCntwy8HkDtkD2l+Zc5HHlixyUNgJkTEnuhK8rle/5jWXmKQRAahB6RizNnzlK+8gy
uNa8Cj/nykCg6rYy6RVLlOD+3vB3BaLCam63RM7Ea2aotVK4u4/9i52uQ+2cIDha1KuLX4W5EnDR
cek6wMHmxeZOOBcuwYs6SMD/0rwdivSDM5bgdAiJr+F0/eUy0Dv1DnoIohH3zzsZMKFrNR8ZJUC6
Hblk4hEGm6AHW5vkduZTLGo8NdObB687Ym4enJcrKm+DxJZTHGJV2sDfvwX9dnLB84u+00hj7FHr
t9BPyoeeRqNWI0MsUah0ND4qKTj2wIagRxS5wNqRKpJ8c1nTKatQhE+R3UMCvfyQ/9kTBtZrLB61
lNcEoMRcB55N5RfJW7V63xtDJ+96QeFqSDzR6dDKUhNIz261DtX7pcbeEn6bC4Uh4wiYs5b0I8O3
nRae+z6wIK8xcgKU4IwqtTg9pftJLtZOTjfV8px1l5eofbu8U5huI4ISxdtfS1rn8Z4R85wG1UwY
yDV0kaRFdfghXmZloqHoOq/y50y1HBiZz8EGNq+ODGJbTXl5ShfQF9vdr4ND7kElzucExE+mvDxh
jLE0cFOmBSe/0OR3qF4yaYxL1u4IQYABRdvsGbVlON0WthlNAsGvWlYTrHdoQx2TOmp/RDTgPBCO
MY1ioAYMbCqmB6BwdMhSfeIxiqTVb9jcUhoNX4/4CUlHsxKWd7uRgUoTUAg7l0zAPia7e6P1JWTG
Cu+M3h/VAHVjITSeOOsA/EZy+wvJbxE/+GDdYkVJ2f8Wj9n7vU/5C3mQ99ZjbzKSfqBYkcf69Fw0
5zei511T8GLQederFW+QgQE9MI2cbeHwcXwexAplMsYMdTiwafIe9CiA2pqRxdua88jwIwZk9FmC
6Eje714+gCD/yqBBhKUwx0v97aPhYvSt5rDTFNQtEvsHesUoVA1+qbQeghLpiXVJ5uiwVo1+pAM3
ouXVa8+FcK+Bd8OSl7hQF583eJkUx0EQONvL2MdOrXj5VOSytM889Vx3lDbIqai2RCzRn15eH0st
bE/gbSnpNnfavOnvSjQ2fmqTr1YdGsYe8YKBjPKW3YFxlHOZ6nKc3PH6ENVDBLoW4W8KZsThKm91
f5HYqjhtdBCijhdj1szzX3T33Ownx3io1O+kORjuZ1MKltpNGmgQwHDSFtZ6OyReMqW7+mHULIpp
i3LOZHtpx1Q2/oBUvT1iGr+AVI5O2FZyKSll9EJLzX1OI7t7f31tNrNr407M0ffN93bjP9rNse2q
xAz+lPHMmrASxt4Yav3T7KBy69o525h0D0d2wGytxxDU1KxZgEodqselLyqWhQTbBMFFjcK50uFK
wb1q6NXeNDtj5MSMyXelPeeQR9J053L6vRf7n6ME01AG8y9T2VhyTFxoGn1FwnwxAiKllzkogThH
v/V6yOQDg/gcGjfIkLol39J1pu7qL8CKMM//YJyIxeOF7dfVLat/eVnZV4yxN9zUbkIqa2HhY50R
OYJbYPcY9K319oKc6Dyrg6bgTi8AAnPJHAO0dJV4ruoSo3+8Q3thKu2PEA1WYrr8DirGn6ovvxPB
vrAdyVmvDK82UFRj9Yfxbmo13NN2FOsYE3ttN7jfNFtfQwnWnOrFLWILX5E4QbLALvrYl/yrJ0E7
6hvMx4jEYxDdztjCI+/kHKVpktaRGg/48nVyOKP5Fcaunt99IV2QmNXa0/Bg9kdIcLpe8YJ/cd3b
pw4e0KmyeHj9w8XzbAM8yK4uoMGISDRxgx1k6i5QvcSPuMQBkPD091f/R6ct9hQmuPynlph+jXax
735uMVnjzPTNmqLY/n+8N28fp+i+hYWw7w5tO0OBbDn4lp/9wtPCuWdPmRd4ErJCHqCYya8r+Huj
sIlyuvwT+HOoIJsx02faN5U4B0EKhaDY09RkPY5WCi4mGZTT+BFsmYRt+L+9JPcHWucRYhCkI3xV
C+YAseHEcsIyCNCuTqCZ0p2TpOOabCgJN3auteMbdB5rGQA6ppdLWxmZDF4pjFPNwJetkrl8AGKw
+JRUBHmFZncZuiFxJOWfzZJzvdWpMDxRdZu3N9y0T6uzdWHkT52SIsZDaHqf9FQ+f7yhYUVrGzs+
Xb+EvIZESoWFmc7whiPpRZUrttXb9NXfS2jm1WDishMlTiG8br7h6GbsRIBoiENgLgWFAMojd1/R
HBBK7Dc6C/Cu8bOZc5u5CyTN8cUKZzkqwKFXDDqWcG7gDxn3jB5vgLCdRe+A74RY4EYw4EyHK01l
0sRFdY/6QmVO6G0pqBE9srwgBmp4Y+64my3KWdua6PuQ27/IyrCP80mMsTR05QRrNCPhZdvOE2Lx
VV+Mp0Cu6Rml/fd8ISCkQk4yRJwKQ3jOPOvd279w0zwdTkTPXPq4kWgsgp4SnB2zO3vcvDR1pj1U
hh7+JGP9PWcRpwGJjq4fadiA4zLzIOWUBx6A1jL03lrRmRCvettaq2ouhxzljZUZIhHGo30FpkxQ
k0ss1ljRLeOElBDb2VHDnIwyLiCYtKfV1rx02afwQk+87ZSSBlLJirg8FaYMLIks3w4iMr/cE0HY
2REjlh3NcS2UIxXixQQNZpbH+92+in8ny8Iot9JL9q3U2EclN0MyBWMqiAQltjDt4ohuEVjrlmpk
fY1MPg7jB/QzeuGKcwXskcyInk5hhQWtBrefLNY/elrFTSaaIccTyNiQmOBJ7WiYVqvCl3uJ2lJY
AiuQ9zce20WTVqQDmozlVRcmT9N/FEa5jJPOlh7pzRmReAZ4ox1FeU5q5NIEhT7E5WZeEWjJRYIM
g2duohD951lZyXjN7TN0WqUGao+LDKIIPKJMsoKz9Lf0dBFK1ilQyG8wd/gDwpvdwBXT5Ez5KVnR
/hWbiddX1y2QJ5XUwefzHx0OGrm/WuRBaxEwBQY23xtMkaw5Swa8WIAneBCzsQkcOZCQa/IcljHf
/nUfooumefmo0OxK7hFRKO4z2GfdcF7I1mdqkIpR629l59IBc1RESAGRwH69iN4uLZX0cviu91B1
LE6YLTEBIMiJmr6GI+5HVPip2W5yf6ulY8VUhXIwcCHNsg5cCLrLRYrykxwWuU9FDWZBNLXvPilM
WAqfrtWFw89r9pVyQvk05248uC3Ws5FgjvgWNyFA0C8vkfPLRux0EFKuVj3423rKD5VytkMCCkmo
s3IJ4OzGV98HogEohVQtV/lnzYRwxp9eioTuMirWqieoqJLNXnp7nUynVB7px8MXe1rP/0JT89ob
3KGIbAZtqZb0d9jXLX6Gv8v32gazNF3l7jGQX98WwWhqt8TOZ1GoTCU5GYZmOETq5uuVGaK3KRnw
K+lOhKbYm28i2Tl0or9RbQPkmX4I7dwZhJ3SpQ3KdgaCCIBnWXtHUvkdGlhS/d0IcRKao4XLO5sj
al9Bjhgis477yrSdi5GU1w0GTzqNxSoW74HXEDt1hB1B2ZERLbF5Eu5jL/fQ0jPIsFiSRrFtb9Gi
x6yG1O1roTsPkyF5GVPADnXdA6v1vwH0MChrpNZ7nDTaaVxYpkMVWtUxdGZjI4KUlCys0pJD2Xfc
Ow1gxvEuAoWMnynBT5aoT95T4BbtYh2mZ51nyEc9BepXzCAvprzNGf22XJM+fnl2u7V6xvjSi2hJ
Ubg050po/C7akvVWc8Bu0Ipj9VDw4xNQQgE3HI1Fd4AuE2/qM6BUIs8cJbhzkjxyhK64kkpOYmFh
FmjXH1ypzkOeCldwFc8e7w4QRmMHPfy+zdwmJXNkAZbm3pbO03h6cOGORowvAydmTB200cbTINEe
3Ud7m03KfW+HGQzkmIfxFa3YZCunVSj0KJDNYhlr48+nbBz0yWLGIU4R+y/NQFe8uwaYKBlaZak3
wkBJZMjqT35SOS3VY1GsecJtHOETrkvlMXq/WmLu0iolcWJiNHyI3tUZeYBqdVGTY/tAK0i5iWaA
+HN6qtawSKbZPxTCXooHtpbeLMTvLMvwTVEoCqZans0Sizns68mFzwD5zgyI0riwfHVzi4gco+cl
oixPtMjxOnzMVxMWsq+idLO1jAfRw+sdqQ+bfJLXTOo6r90ZIQdmb5me/j9HKw3zqMLrVmyZF7vB
+leXe0UCrgjriFEmSN5WkYIYw28qP/VmLiUFBr9oC0R/ACeXxmMBtXJMjfMuy5CjFwUPiuaDzCdY
KBYU2xGDtjPMxoSZDwC04wPkgzQAGFSQ0RYZEmjrDLIFht6Z207hpIxYGLEGHJpTLO7oSdQGFQEc
lyKt3YbPiqQVhX7zpPJldw52vtX12yarjM3vCZZrKDzhAas3EN1RD4SDrzqoqrVmX0RWnTZDSBSe
do2WTCGbMMmHM8aY1/L9eOgcy99/bZbHFeJVe4FTGjVNJ2tSku5s3voI8JapI0nBVqHxvOpuenJe
+3O1ylkEUnWn1G5K8CgFuuMX4Td75UyyWcSM6s3TSwKKTWKtLh+m9nITsYV16v260PQcxibwOisv
uGbKqHCp51zi5YZQchWGzosqObCW+ZzyUXMSDKZkzTP7viq5XD8f7SzDQ5FnFSnedZyfhI/xRN4C
KuwN0XhACRCfGevlneXYlK2Xp2TkvdGZy5q0RZODidfTAKEOReJ6jg1CRT7BJXrTJQBq/e3RFBJH
d5Ut3xmnHcJ3vOoQZmfwB61LVH9ziPTDzIxrPCUdAL5mwWzH/udtzRvT2oU+pZ8l0bSQJE+THUpQ
ls6zSfdoO5UlSdSuGAhndESwwgOT52MsQ1kMXzggRr4c30o+aRtvRHxCvBFXpLXTFo5ZW+O55Vwd
KWWRQUyCMggGgb6eNMY4W9E9c28+LH/Qq8r6M+SKtR57NY5/ijB3NEsUh7Y5je3P83kfaSGKqg1D
tO5eSZtGAROy0JQklqRfY+G8BbcQZwZsfrsiNZdAizBYfN7UZl+H40jc9/+FnIWqG9Yoa+KiH6hg
ee4W6Xcxl9YKeG3FxX8on3UX5JvTBk2BwgcYX/hBxUpXkQjDyporNx+c0EuTXTO+8xcqTWGLmKxs
nCPxiMBUj6tHuyplEyZ2q7FEEdmPNs0nR78y/l8/wIdoWPpPUPL/XxS/NrE/HcNQImj79RMSOTDq
31QPEgbO3tAIwErNTuwJQJ/PwtSg9dSYPZb0vtGx9b3I3Agvfp/Ujr9O2uHMqNevXzaIaIHVf7Li
002DfyByY9XYCotDR9qv9+gKc4pD/BDBvhhsvMiCcUhCvQoJlV11Y0Q+timMQz2FAz9coCivJKaZ
vLaSPS6RyaB0ktAeBAy7QTJvP1xxY7K9thq5hPSvMMQ/tZXGVjj7lnH/N9cbUzJWFAnAssUILbPy
f+N6aKhS1Z4iZ70YrypG25QuSQr0vSEW7Xx17L+TC2zxrtkJUbDL0HTLXlvkc9Oj4Xgt8MDD552V
L9H7OyFj/NsbjddqtfcvLkSnotnSxWjpqxtIUau96d/6MSzzs1h0LoWca+1y0wl/urM+zv/7+fM5
RI3quBTT3LMgYJ74nOkGdXDan4mU0LqnFhTO8x2xz5fpNf/p7k3LWr0ZFLgZhiZ/55Q+7KGa+kgJ
NeSl/ZYoQQRN7t3KDXV7+ZujWmTl9aOUn66+WBcrzLV+f22iCifzkzpJZqG/FKBLNOiYPk7AiwtU
vmqYrg2r4r0YJh4llyElo2G1RxuW1HKzLzpVEszuHBEmgfXR3KyIs1YdsvwlE1akw4jTjNGXYsWO
MBJgsG+3pboMb1Lqlv8a65Okj6oiIKrpAuf1y4yBw5PxnJ++zFjWgwIG69wdTe2pmPOnttiO5NHT
eFV2NzDa3uspJOZdhsRMGJMgsUtdtsJScBUkawA8OdenkqpU6pAWff86H805bJ87SN7Mcs+rdbsP
HKV133k+BjINh4nbjwT3AP/QAV4RMAT9zs3EkE2ptoDvx2TYG4S6rsesoKvjCbkxV290H5Pjil0M
ka1TgxLwLqa0aX7VJiC5RadYNivyHvHEqKXM396PSnKByil4IjbqiOVGMqah9vgpr+5h4Qc3Vlcj
nnah9EF3/KOOfEVs2BrbcjzoK6TBUYNUT93741kWB5o5XpJpUhTadbLVOMh1Bgqwg1sbO1qMzDcb
1fW5HeJ6w7nybxz+JEtKsa0jZU2AVVvh+eBt8Xq80+JD0dvK4vrG9xEK0sMAKsTM0wMkPCSztFtx
uclI4HcXtaMltmA//UU+b6uSAsuReIfsCQxYCcOwbzWL0UfW8mUyyXg7G/3h8/JM371jNJ4yhGro
+rSlPj+XJrLXA6uZ4+CddWiVWGcuXHc7uTDo1b0sAi0oJnjDzKNZIZtflCB/O3y3h0/VDIrzsK5z
QCwPdrTLp6OMpnjujpAwnlHbQ1rKvSGPyYw0cm78xFIFhEZL4IOrDE9zbMXoGQ5+4q0DgdLFpRYs
+qLm3Ul808c35s5G9y4GCO7DpxFuTxUKdsn+fYtL8aWJbnW9q/r1U/v5ESJ9P1fVOvdMGmzG624x
YMSJ20ICziQsmRNaMs6z2YlD32S2kwoyyGwnW70+Ed3mFh6QKsMceaDjhXyue0PeqeausVANCIIx
VMoRqV9cjTBynRj4xAd3Ti/KE0VFbjfth2DxNMs9MJh8FmglKMNTyojRDTro1GUf4Nvt8ZZ+YzIN
Lpe2lCX1XGmUTPo1qke2DWVCIUCeKNa5nvWDl/0YONPmy87RFnvX2OYWLFXIAviMBspkcQzpPMoi
Zg7oOmyI6o0g/iAJ3SMpf3k0YODY9kWGvXVbPc0y3TRCJNiRgdj9jKgjkRV8zLuIsfwFSLWyHw9I
jxSlQTR7RPlolSrHKmZ1U58gIM0ZxXqn9vCWUYyh3pR0Wvz2R8TMU7rHxttJRuStp2O2sGzCNUqp
vueOANytPkp4N6rNb8taH61PLXdUGACoioqci8i8DeKVmwdaS770WCYUbmf2ynPs2I8wrvQeBWbo
iWIZ+I/d6joMF5Qbfa3HmPsO9+q7rBrZwuuLR9x0tGdOU+QTykejkJIEyI4SpMjxgb7A0WXpdOjy
e7Dtw7aYSqsL3DSRk0wuQwb7NUZwe8AzQ5U2E0Tq0TxmJILivOZ9W8TpXb0XQK0BSK25/8wM805G
PBrFtpunHTrFjV8hEPVdZPfRRg7YTuSTd6YVh2VvjJknyJPHyNcja6/CZfj82Sb70LmdMYL5/gl4
yiGPF70PwSpi12ZffAZmIhQSsVU3sDQNTdKz0vl4damlcsppJbyNfoA7exMTBWXKjIc/O8MmVHAg
jKe0TRHDIPu7icJfnYfGMt7wVJ/k7wzpVOd1pz/LW8laTtQq2RS9ry3t65mnsjDLdDLXzKEGWDiE
fkJuTnPLDOO81RZikh28nx2pUgild3R71vEgI2SxtGlNRSLlD1iXOQbNXWE2FaOqlm8b377cTtyH
jfDh2msOqNOdRzs3V7FcvBUf5F+6qW1aN6WwFqWAbPSXsj8LghvJze70NYPXXZ0kd00MF0TeO0pv
2FqPn1Dmp4zMjwV9p81djzkxZS+6riY3JonJ4s1hEVsT5WXnZDV5XqNV1fOX4lmevN1RH2pHNo9D
BYLEox2EXNEIPKhQE456UVytHc28IgsGAB0gHY93u3cjIz5Zg57zEsunigRHBojarNW9qaNtV1lv
KQG0lSj5ZXcq+nIHf988xOcb87W1/GfsBesQgst0aVKapV96+nRyNqAauRTKUYL3coimEuP68kkk
+jnHY2i6RdG2BOA0/IkvjqzSs9Hl9H3OjgZ2X3eqC4hQ+/REOslpitQu26sUh0qNxmO/X6T6PBQk
ZqqGaV6L4x16RG58H3VFKEcUaTJ3Do+1J2PYd8/LMBHEAE+5C2YKwXA6MPgmqNfmF1OvRf1XB8BT
qCkwn9ErjX4Ckr6CzAZK3IZINB5qR0SyR+THtJGsBtnyQ2YjzrzlutBYfjMHEsaOYr/oHN4LHxFg
A3zEITL8XGi7Rm8nWR+myegGuwHPvkmfneibihVRgpUvWmH1zyDlk8fk0sZ9VapQuBtfhAUG4YzO
G2gdOzuF/dTlj3t2PrltTecMkpTGuLKmDWq3GuHIiQWNIWmVuQIWfNv7Rjw9Zg9+LbXP2u7eX2yZ
yFlaNWwUAuwzim331hFVfrTd00MXFYh6yCfJHWeJ4YNLRQeBLjL7LC64rw5QNr86FxPuNNd55WJJ
95zcltB5aIlwCBTrDr2T3yUYTXELD8qE2SbvyqGXthXySLMjy3CdMbM0w/okMwQPCQ2eIYohKP8w
GfiM186qyWOaLUlDSA5aUc6mhLemtwKZUXvZcNKRVOLJWvygNd0g1BxslwH37e1NAJcSwBwooCEu
17RndMLw0xKU2fZp+ToVtKwmiWZ8nyVjaJrOyqkBR7sB9T7CwzDNjVRdWUOxjTa8cEjK0p/xQUQc
vP5pcBnMg7jWyr2EWJ02InlFRedEmeOrCgIPAfkxHIGiAn2eQI4LHpxik6cpW5PwDUlO2psGIo0r
SNTmYMxy3erhIJsAAubvnwplhaNpKv7zLItxhrXoyaEi1Z0EABFScq6SLtnP3aEY3I9G+iXdIp/f
p5fgtPPnU6Ifn05Ob5nCWliqN+fQVuA4vKcC8LPnFf9zum31pCkPdn58J1TibrH+Sp1ERZxcq57I
oliLgCyDlJ0QfOvo8x4qYTNCG9Gxv7IfVv/oHL0VNJtZ1xF5vB7rVeIyoOYx9NGMU2y2ux5vhPec
QfOTIaGQbnpyBwWBg04rvnEPMXL3k0kERYwmQtV/bnGh1UPxdt2gPBOGSBHsCvy6BjQwjCBdvt4K
eiabrwKN27mSI9sHQarWXJpwO/Fxrs2/iDaW+Mox7dELFvNK06ghd3rg7tgtBoWrMGYjXz/uiKCr
IWtYu1OJ3BAoLfICyFmiMLVJ6p/DTtnMSFVTrnL6ktvHb5vc0Sjt/0lxMkOdKpHScePRMUo/+vIC
j3HcPe/+/ux1Rx/DRWInZ3TL/fXK4Ca2rlm/iKAKeB0VpFp8KEHVL+K3KiN5jpYRemFKPSX8f/H6
YOcrluYu5kOU9TzvCIYg03eQAA8MXe9/V16vDPwOnNfcz0SZiTA9LyEF1dlnvCdkJrBqe+3orw+p
a0E7eTt8vbjuEUaNGtCLeOQQ9xfDqphWFUa74kFq5oA46tTsj/89kiITsCjlkBWaPOTxHAHDVXQZ
dZenhslv8u1kOc8fT2cztUuH2m7SZzXA2P3/01FqR+n801cwr2p11aDRGa9Ys5BDm6LtgaWxBQT3
One9QS1QaAuzFOs7qChK4V+PtGSmzJVTITOTrvw9duqGPMERFn/ks14pWtmB+TGCgvYwTt9URYrT
hUaZmPLyasiIrXdqLkDkdTaSWldCYu6yl0fEFujGiwdHxP9l89/dyLZxnTLeCyX2/UIEBufsy0dR
VZD4BLEMvtOkA2hnshhJCUoGXUqFnfqv27aPEJvJH/A17yUShhAx5z1QP05GC2S/brpdq3H/0yjb
qDGgWOqQd5sTta+X9P0+auaSPXD8LfjmI9pGHF9jGnpqcrzc4eFrf3Vlidv0xXHnxreAIHT628TH
O3APaBSbU6oIStJ+SnCT5TZDjhxp/6J1oKLYC9M5001/qfEL0nInQs71RBKkFiWV1P5RbqfG1foZ
i/HOyImsa3nTZHAJI5iyXBWzLAHbzs4kRvMJZZPo+T62TA16P0jV21C69MEw7rQTL+NrT+1T/+dH
p9hReqfGf6edLN7d7mDzJo+kn8FlZeZVhEZtLtsDxv/FVmkJIkWYHzw7xgmaoQvTP+fRRqurUTtQ
oQ3vLKFiabusYafeR5MqqnjW8ImROZ9W1HVL0rBzqux3IK5RtVD2LDdrPQpBXonLXuumzJ7t+gOO
DgL9FI8WwZQwAlNnDCZ7gljzrDJYa+GSIaWLu60Y+7MJ+HMVcVyNTfBvGI+eBjcLhlpqjg+IWAQa
A5WBoGwk1bqQNKfU+zcW4vrRc1FGyf9XnylObNCyZ5ZpLNFzHq8K9cKYtClqSchObjfb4gw6v0p8
YqIuqHcHheD897lgNQdvXcVSOr+5ZEvpg/bkpk+qkWDzCzcOmWxpl60E4RJxCmgSAf6O0vvBvzVY
Tk+fCkNZBjc7nRyP5jV5V7D4P1IsWq2Vs5ucWrwVjUUcemX7DY0EEdM4yPziy1BgTZ3kpAxeii2e
wntcpak3+BZTJPzk1QSJTEpGQPX+rm1skqqC0d4/285327q6kg+DoCJAVDLarOPnWgSbB3Wa8/Wk
nZBRGZAHL3KYQ58kGtvX/FJ3I/UQyJYxvtbqCMOGQT4wz54BcHK81q1t8s3B+gWdRjrRZ0jLQlXa
Nrfn9MM9IlVmrlOQKn2JdsVJMQIZIXG5k4zJJ4zdOrirEtL0h6vXPJlywMG8FuZ6xIYhp5a0W02z
q/aLHcAF44TAW9JV8p0T5K3+9rqu/ZJmw5klNAtK0gNAJ4l0uBsuQya/21p6k8qN3Iv7am69G1/P
+3xSu2ly92j+7eEHIVp2zuuSipNEIQXNhZ2Pl+H7TxydAq+lVTSqRbxb1gujbWpDVN6UjcuFr3WD
5g9QY5eVzeX2sIBG7CMM9Fw0QggKrqKRxIKayBnxyhZeHVUUZQJQOHdKQbLJVJUYrkX0ukwN3VYd
Pc1xKlr8mZn7nyjX6uJaOpzMm/lhQtabEsS8zayvTOWPUtX6YZnLKSnarlcg2ti20lWC7pLa1fFv
hFtMZ6w0UvlFjRgH5yZRaS9wiImMGKoiUnIT3wUz5YOAHVi3KkfRAoGXFNJhGgDLoWqNTSgrkFEG
IYc50H+MidwP/PYP7TJCIxMLSNFlyyFUCX3rzxLqgImHX8CfnegmnPSqiRmYgMu71SII3Om6U+cK
tOZHXN1LRt3SMX1TLXxuByYLQhb5Cm5gFHU53068r5CAxP6mxPuYBp5GmWyRYiqGW69+9CjBhqbc
+L+LvkFydXgYYR6woLIUpURNo8e3aTQa3CUvnuuVx+34wXtDtdk+AeKm4foVE7NDdeSuiOtsTcv0
vh5I9m6nh95tf5OPGV1DBIkv+qfL82fRtULaPSvZ4lBMEmr4HHLT/iRc5h3n4oLnJv6u3M6Jk/qr
13AB3OguLdpBhveS13SF9xFNRorXMduBCvY3Rfnwk5YILxxLcU7q6oen3paMjLCyWAdSVaLxRjnF
x7FGcwKyuxvWX5WOEXnC1Hg5y7BRP8mm1n1nPia2cY+iOJPQu1vpMEcuI9aTYIsSrJUi6Db+48cJ
/ctvytPKuaSsO5IqyR7H6JprMU91DXkfok4A6x81yK1/cmf45NaBry6FWwXb2Z+KiLK6hsRPOnFJ
IqGhCvv8cy1ltBOEbu4trV1j0pN/ES8lNaNDJxxjpHeQM5FWWCVNQyUQT7+j7goBZcR9B+SQw8J7
tcUHXSEsWZMUKZj5BEoOXLlmgXK0OMPLN/RpvCRDbUkPXSfwrfzxhVvQXOmXs3qmebJEScPD0Fvv
+VJLla0Fid64qjILYJ2G5ExYJP9MBZTjQWzHzai+7i/+f4zRhcQbxJ3yDYaQnwLRgy8Crv38OkA8
tBriktjfQGmKXEjxVC9vg9r7mty7l0PUt/usGN1l5Rlexx1Yhlj/4c4E+WhFXVuUa/OCQscNAWBy
LjEgTNOAJOeCUdzkygTQVpqO0qt18y8OY+OFgkELRpZwZdAvQ/Ojy3WZsLcTFn5u0mT9kRtbMgzS
WpLy1C9mtt6oNr9rgzuEbuaQpBmb7KnKsLkN7pvyOxqbqWUUqaC/5ooHi+s7RcptiN3ZSTWs4vsG
LW/WXTLMFSxzbTvB+GkWG81WczLc0tHh+0Oefu34FcHFwvrXbfmpR+mAjl5quqkSEVXqa8hXI/TF
gFyhQ73Mrk/5ockHQFiYFopypoJg1B828/daqFvu87BbrxLL2DvHsbLad5sPrtXO8PvtzNbsgMXT
kqFHGIM4T8AzDfSNNXG9vK1wjrVwFlx43Ob3gKI+8H60jpsUtcyZUujXxuC4fPukcCRmHRNZO2wD
VK6uvLXEE/HHEf2mTBWhOgXh7MJItfshJc8pLKFU8d1WRZ0IJc/ywyD0QnmOmY5p/w2CwOiWmQ3Z
5XPbSP7XgGnMiLWY4+Ibvwz5DxlIXPQXu+zCMHvf0b2gdECtfyvisi+7QKDiQAzxHEmLA1byds87
t9A/Tsjz9WIs2dagYKF89xRvBHu1DxgaQg6pmW0IhyMa/wrZtZfNxaVeyZSvevY7/ssAEvH/oi+Z
Y3sKFqagS9WjeGtLhwTEYEXDlAKgBp7e8Qr92YZMqeLpd81mRy9BrkALnUAfXH0G1KgY/pn2jUp1
EIcprjV+Q4cidZVfd9Uu1CsGTlKXHatMn4SKnv5SPyP1Hbm7g73wIyfJXRw3aJj+atRu3yIGB268
zfz6hcGgo43PzJaG1H1LpmHlydxdDnS7bzy+kkTW37XXA+ive96+qEy9vTP+nzet0Hk71cNsWyt4
gcl5CTtNQ5f8E2PTTazQWPbpuhFwZhCzV3zcvImHLog7KqZolijKxacAe/9UwrUQ9Zdv1FBc8jj5
3qBUvqkcimzYWydVDztjZMJfRK8Yk3jMM3am8QDxLu4Vn5+ymPPpXvGZya5+XO8eIMX7DkDGO2KS
vweKlvaLsse2wyewwW/9GrQsYYMVF81/iK7KmQIOa4SdPKC9+ub9mQxSa3SJyDc7FKWyLENTgj9o
gfs8FLX1u1J+AmURAEuAAkZ0Ffx/Isw2+JIA5dl0q6vlunDYgZwRDxIFyw+z3qTYFeg0Dam5h4vW
0AXbbenoVLIcsqJxDn6bcaShWwj/0yzhd12LiFvvcJZdZ0wL1HRfvau+YhB/VEsQS8v07irjhRRE
hYMUk4EFzclmquPe2hTTC2uJ3QOa2X1Dx9G+hoH2iJT0xN7F8RByjxbRWQdfgWYJZJ/6kun83JCz
67rNd+bMyub5u/AbOToUPe2x0OsU1HuEF3RweUCucnxStbfxg0vfViBXPq73AtqgK4BcostMswBS
YGMzvmiHzdn0ezi85It2mAQnGXL7b29twI8v1is/mwGrZ+kY4fA3dJiD8tZvyzChJoM9kclIMYDF
EMvvVFKjApl7sjdtOMzA3fyyW8tsF9erGPErgHkKSk7GZi7/dwaMyWAkYLcKY8Nzy8r2QvKsWGAe
rkKZPPsYM1sz1T6DrkSHbeS7e9I9xshjihgTNEZKxPdPJwVzCeMo8L7U+A14BYAMfljVmt1GYJJQ
3CfZxx13s4Yl3V5/Ut52PDpIKE9KQuUriIK6Uftwr+tMK9mYzAyyim+78OiuMCxYKneEaZXqBTT1
5x/emfSChvFvCrXQDZsxwjmdrCnbsL5F704bwYLnmx1wN0wfX0he7KKR4aD/C8rUUumcgbo6rhrD
cEewxebaOfsdZHUmzNeuruivmW+wpFRIy+c4DhJskEH6QeOtz6I7Pgm/KudB725NWtOaP35B22fo
a6BMEp9WUk7U4cKH3RFU/tpNhYCsGVYsSu8kX6JFVwtgxqsvJ85x7PUMIVVt+7lIPxrLAyRr6Hzf
i4CiDBes+Zznvp1Rn+ntiWRPaYT19zyFdDHKXs70CusFoLUyWVZJOJ4sIwQ/9mA/jNYK+Wka1f5q
Q9h7qUUj3FpAbuKJ9nK8+kdMGkwl4NG6H5teihFgHzU7/SIqvpPyRHV8XO9Bbt95Ti0oI39pZTXZ
AEsFE5HPDQ3QjWuhKGdvUA+i1T7Hm9FB3vJ6ov8WCI6d1GVsAgCTYzReQFOpwGw+ZamfmEDaKDfe
NbBuYQEqYB9Cdu6jE61qGJeAb2tUuIQ8JxZ0ET9814W5PAfjqgB+hDXaOVVJ7Q70jMzkHLi+aVQX
J9z4UIUeyMxNqUGqOq5BHQj+6xr4R0rHbUqZ9FH/yk38GfTSvREQLkoKyRKt7iDimh/d/o5O8Er0
+Hu2LEK/iQMBo8eVr9htGyFM8ysNQQtWLKMHY9kvA4lL554IXXUD6ukeH5tUk2UQ73toFDjVl7rz
KpGedPhHCwY+Fd03mC7JAlDVjVpXj/94vvRGkOj/mc2y10yi51Y1lifluymPZfIyTI7FpEjFcgxx
fI/lMGXD7TM17+KfbabFpLWlkkB8aIPdpOKdCQDGwS+VeVYyf26IY7gLnx9UIX0Y8xgmsSXx13Zz
imrt10Llv/7Fcot3w1Tr68sFtpiXMDBJ6dDQkrEEdkr4PnJv7fZgjCkALJi1gEO1JpeJNtei9KBu
rfN6KozsiRugOfsEK3j2HJOc8s02IEnRPi7o/9kngVZ59H65GyZjZQJ6RFRwvxAAoj3KE/p+2Eqh
TS25kyYDy2L+vLaRa90F2fSYtOiSxUDGeG9ltWGUzGF51RfX9lR8CSRTkPLmbm9BM0dBTihMZj9h
uzCId9UR3LgohfFWnLvHrf2ao3VXkxCf3hXg7C74FhnzhAVWNPXbArwucBFNkOretVJKzmune/bE
XbNA6UC7nB5RzGDA+plJoajLcpR9M/bExtWPAZjMgRpkgyihLdSz5pzMZTvw6IULkygZ/HGd6Raw
EJ9zEd9/uRPjPnxCiYHNxGUcARRph6ppD/sc/I1XiyEIZaMw5VyPJ0Rs3bP6/a9dJlLJPaFRNj85
Bsd7pYAVZnrNAoIxxhaeiMwL8wbn8Ee48eU4yg/JpQb8e87tNwXEzwUOXaskRrsxnoTGhwRSRkQV
j+IcnWlfQ3MgW13q63KfTnofoZbgTDwNbJGPboGzLJnZP3ATsxrXehG7e3tULbR9XcunX1uA4pa5
XkFAPG0X1AvxnA3gt3PEYs/YBM0tJQG9KNAuORlSJPNVksLLSevsK45SuE0V/q10hDTTxZGCki7F
0Iav0FBvLU/Rlt4uYgviXVP7OeaaWWPwGWLXHO0xVwFE3x8ki71AuS63+KO6k5fWRjI7KgcHosRN
xrjEvFLxIehsogzAEdesliIlzDMwxr8/z+CnmN1im9c55t1MJUtgwhn7ioAGmD3/wxwoAolxqV/u
Jx08tLIA3j51nhpWEQb5q/N0DJu7zZfi7xvUpG7N7+ZpIsWV07MPYF5q446tOHYGXtH+fRr8Wxb2
5joJKHdysr39Uio9xhlBQe1YKZ7gpF+fgho4GNe45rPxOsUTppzWxVAtz/Qos9UZd61j6cek2x1E
QnQkmlwSKWPrOpcOzCRShTcZeuGquq+KsamLi+iyU2+ZOtOQM4P3Azbl/CrMuyXo8pqYTeAWESfe
Tm7IP8z6WB11dQmup8EsdYUDTQLxVtQqZ5j2NiXrlTyxy2Evj6s0X1ky6MF695w4k+SLA0knsRIz
G6L+vKxvcOsNfNqpG2ZizzWHA3OvuZ2/TUHAElOYF09Vut92gXhj1JJczkXTHMISA78IUozyEOOT
zIoryVFs5LIOsalkGNDzk92Ok1v105odFWEUWMIDxfwaoJuPfurSworF+R6axhBeuJ7UoPuACfff
9xrMnc3msWzPT9+Sy3MBZhhpFa+pA33TlVyuN4xUw2JN/px/6q9CMkV0twZduD3SNwjOYZLGN6dn
DyfjwTkq3JsNgAMbn7SIe5iG5Xode9328P/lgxtddEtk6068BsoZ/Uf6Bi0AMLM84lC4vocojYVW
tZxxVSNq173kqicjUTZ8n/SHySSrEAeZQ/hzzSJ4qXHBuH2Hb7/3L7PLAh0LFNQDuTq9F4snOepu
lwT5Yc1PImZgGBVIp1ua7MALbDEORYXPpq83JMoKtDrL+MOQnD6K76a8pRIiChSnMo0G0eXWgvSi
FYFYD4e506vnQE0CzvNVGmOv4hx66NttROL2/PHQ8ERvHzPjmgPsn+GYicS1DnsbElipMJTLw6vR
KLtXdC4vAqkjofnGqW+Pz4kzZO7QncoXHvM4ztzN9KV5f+RDGJHP3qfUmzsMVDNIAM/bhKfs9NQh
6zt+BTvfYZyBAwLrO7t2VtwXObkWy0nOkDAhHIbEF7jKXw1C0uylqj43uats2TaXUP3gPuD2/pyo
qxLWX5fqlhqiZTjWr0lIqhrGxqCBVwKwlyBNHwDpWF0nPGIsbjZA20lgDIp63nsOmivx5VvDsz+U
AOAXkEqweVIVOVxBan2GhwA+EKDRmnmSushaVXeqNLkhpXCi9+72t6ugMgYj+1dtreifdoyN984i
waAQ+/EXvVv0ym58E8CwOcYuB6R+NvR0bzBF2btifAaA8l6mXxM2BbkN5rinRZUrtcotlXSvcecy
XYsdZjdJhjeItZs1UwAiClCx4iWy8r+z/oOT1Hjk+jiV4/Rpgd0ObRF8w4FUE2xVJA12neuNmUI5
l7+QwUaU3k5sqdH1/dw9m1A4ZCvAT8ZS8Bk4OMx4huKJSdX28813zAUzgSmqYGIylqOPGrxydcAV
TDI0p93LLsyzmIdyhmlcwkKBqEDs+tJ+nWpQYxBc0DfKBF/m1VNiDssyy6LB+4sI3lVm8lqtGs/x
JDmHl1nMSSVAEVFCqF5MlMK7XONyelisEVdoEkcC/WJdhlUieVAXowVwz1xxSC3wJMwakDVKPZeP
5oz2H/hdtLfhan3zY0N2dV462BlUjHbZqmjOJIMM/QaXqGBTAIzqAkcaWJqSQaIEaTLai/v0qSJi
IYShUehf7Kk/R2DsFG59ZJAjrxE9ufejRDHKgsLizCOzB6vVJCdutjRx+nkUN1ZYz3psDmo2iW4X
KBkYnJkgBelyPDsTkfqzf4vGYFSOxl9NUo/9ESn8Cx1EmYb67VGXY6rfL8teILP1JiI9y/fvRf7h
0DjjXM3ajFED729YtsM+nGcPXoAQ4075Gtcb8k72ucoLx2z4knrLxgG9pZ0EmeN1P76YWYmHGDkP
SYU86kTAtPXohPkempzhXmqL5h2IXAntDaSudGkT4uCuUB8DjgnfEqmCq34iQhLrihb5xQ2nrmT4
NVPOMSLZ5Ohz7HoO+13jNQ45bhKf/50o58X0NtgAmxDT4SVyalcvp/BBoRL/qtFDY0XerG/ak1MK
UFjWsvgwWK9iRuxfyx3Z85VN5vrOrkXhtmv0O6djjgDknAbouBlfpBbFj7IjwXLOWWZU8b3T8ddk
oJCG7eceApAs8bL23ZnOO2uZMz7q0x2epTrGhWsr3B7OSTA+zva/nO82gSIrpUQ6HeAZCWkK7tkK
6n3ZfVd6NwAQyrwcZoREK1lvXFyNAxfB7De1kVJg9UNn7HozEXiv8pQtXMvBZ79MoIUqSSjL1m+f
kDYubWrZjEgZGv0tJW3pzM3zOnr7XQJNjqmUF3+OnPOQUQ4mjWmldN1CTbgSU1xRaRTdEPD8tHfs
0ty5cBc9eYRB4ebWcOFlNhmh2b49GPrMUYPtfC5KnhHiV5lqlLJEYcIjurOOJWIdtbhOdPbp4jYE
5GnygKlDWFSfd9xYNwJQze1v5vG995E/EoF8aWN44ig6PmaKoU/qmt2xx5+0MVBw2VXZv42/kYdF
KAgQ6nmHK2Gc8arxC4xtBPctTkYemS5ERY31203efbGRI+p6N1UTEbSP+6IPkL31upRJ3D98aU/6
RshTf1P6vUv4roOtOcCBQeEsk+Sy/2VkMxYMQ0tVk/rvDyN84NuczNyGGYL1hNxh/2UviMMYdOvc
9mXNuholDnxVS9ituwI2oOkGXZCR2EbPGrvWrq36HSKIfOqZ4ttafon8SXea2WCKEcieSUJUEHhQ
zkrsZW4ZmH8uyvinihA/8Grv5YWcQxvI6bMBGjsFUrbHv6TS3W/X+ypvmzAS9USUMGelGSWI13r7
TjFNlLA5t5oDBsv3kjw1Kn9qnIU/grAKQyCiu++MZGwX1L5aLJmTyUS2ASf27qqe+u0rEn/LODUQ
FTlfwQFUuVtuQkY37NxatNKoWx49suy8OEwhwH0FQnYB1mBy2l+fr1sAQtdK3GKXNF50vCmVAWVv
+LYrgS5qHejFRnixqN6E5vl+8N75dpdr3NsjyBuEyi/PDUqmR9BsssZaCZnxm43P/RhEnoq3mExL
VkGWO/VJzrsz+d6AapF0EqMSiH6s5zeKbsaTjMX/u+bcMch8GVX/q98uhmHWOyazSv/kyu+lzzD1
SoabaAyaZ+qZEJTDt1orhrH2SEUDN1JA+TWohcuQWi1y2yBqTAXvVBIVogDu4geCK6faoRqCFqHg
9HD5pJcxoQGKsJQSG/eIOFPekFpZBv6fAGn9urCblDlAbHGbqMsCzhzC6L0rSULRBOHsvyOJx2HW
cmGwEw9aN0uCrOPZS4sAjaN2y3SwwjtAUnrKknhD1baV4uTeiFVcHnOK7I55L/18BJb33qFtvOyk
ME4PLROUiqhRud3ATJR17wDUFU6bbv8Zw/WjAzwd/4I7VKIBjZCVvkvlNB3QbuQCBUd1j5BubwBR
UMkn4W6qlk7KrLR2+T6UA0ztrXr+tctzHWEhg1elEcQpVvegiMSQc+WH2TQ7CzCLx8CKIUdaGVhl
gFYf8VJMqZkBvj6c8Y7XD3zWN/IBJHJ2mN20E/lZzx+22N3Lv/oZF0BH0lZuKXSkW/TBnUFNlHk/
Wgb/AzLegW0nIW7CD9sIyma+FHXMR0t5rT/dip4lAoTEGxH2Wxvwqw4J5p4b+km1xS0iWiKW5Lcv
SBQ14U/xk4zldyDde+VngbcIfda9dLcCaua8eWMqcPaDv3n/yzC61w/gfd+Q9dIVl3ljcFK9FSV5
j20twxWI+zouFVJ0QDu75sq3Qb9JY/YwUSKV6qwofffZgdc4BM9kU33WxoMbQeKYOZdOQa2siiZr
AWPm3KtzNAX0VvxYM1fWHR6fqj2g3fIdV/96J9Pa283Tp6rKSLlMOad+LgdeDEXeBPT63PqKVCuu
oF4ecjuHDhRtHcu2HUMlErx5f8UKcAgTjSUjOJsmcQSBbE/PEj0ahN4K+mq+8BoeTvZFMoHHWVoc
fRBa8hPyMLFo+xlon6Jt6xS9FiSF12KR+QAu9u75oMTJeWkPdPGuDXEFm1c48C7z4nQebRuQ2ETV
EBOzItkDJt6AEQfzQ1Obv8TW4rwQS+8ZXS+M+9eNPvp0t+FlqAjku3IMGgMXVsIh5SR0J36MlbIi
H4OJ4hSlK+JNELeZNv8KRM6dI1qtT2e18ojWI90ZhQw76cdTHFrGV1SlvjAsYxtnwo3b1MpQ5Z9z
Be+GE/2j/Zkwuvay6RscXqkaHJlX+2ZvoprQ0rF+CVJWp5nfM/lRKLJ3GIevh/8Z5UYqK6Ik68nz
WgjST6oCNgvpICFSDn0HXCalNY2DlOhoXnPxi33pg0E5IoTHJk4SARXJCV3C4J3PPiKjzPeqdcXk
k1Sxe5apeC1SRy4QRSMBRUzal9SSPtbNx3Vf9yyd0ceuV8AgrtGsxVmKoWW5jo94hjgFSfkEf52j
4j2h3PAgN9B9rVxHl8ADjrEawexd2TQYLu05jnvQI2E9rbeA6Ihoe1oC6WKLM7/XRRcAwIy3r3My
AO9Obi6ePYHRTxL0P9Z9CZpXJ+WAiLDGy2E6HH0N8+oc6yeXu1+m7Z6wi0m9K8jgGDekBuki/o5x
i+IBOlKVirDS6htEeBYBnOUiyj+aaj8VoCwX3rRMVWaL+p0NZOQBoDFzgH++ADE4mEqBz6nzpYIS
uOcFYrhFh12p2SMD8wyfd/MUdK6+PZx1VYqCHZoUC4vXqO0Qu4cUoVX5h6/EketxX1XVfADbZM/t
Va4RG/oNsInmKDh/C48vq91nldULdhJ6TjijpZEuOYCo8BkSbTGyVgemJsHsoYvyw5tYF+HSjBbO
3s+L2/IWTgWbxdQ3tu8wbejoCmsm+vgN2/MGz2E34bdYXkagua4s7vNRxA9guBj6rX2kw5nX9mJS
rMgELvS/zRWamo4nindVvQZXb0k2DcDHfvkOI8dD8nHNnqQ0ptGNIGNwjNgOf5Pmi3mAx4pWP0JU
d1DZijBSYf+X3JSqFmykgyV+KKva6rP/u7hw+22ADphvAUMxKXNXeNgp3rGoW+q8gyRFjTc70Bod
oLtF1smwGvKyQsByA3NpJOcl8Btrd+YJB9r/YfSFzUaldRME8MTFX6b7+HhywewceJPSBb6bqBvH
LZ73eXmpxH05x0C2BSpLHLrzDQq1sWe7piwtH8y6xFmkCIrorYyZwlhBM3cfHiFRD9cQ8c6S1jqS
fzZazSIkF590EG9aUOJmYdfLn5Gue+GS5MP1fJOYxvHzetU/DU3t2cFFL4e/MsYkJg/dEn0LpmuO
HdliHW4IdagXloFMZfKifOsBEg51nl96bV41mYWz1C2JosdcmAB8+j2pknQVLiW7CTyS4yXTBMQp
yQN+BD33dusN705uc81hpSnqZh7R6JZI6vwpDwkfBnEn6r1RLDPjO8uKnM8MtHSJmq14IhCaKddI
hSa3S02SrJXw5EpnftWOki9ENu7A/hKri3dfyS8m1/rEfdMQ51sAF7yq1fJknE5eYKUaJB1ICaW4
WEyGwJkqbYag5dQcfjuHx1OyXU2/XEP/InsGUTzpPcMxx9ERu3ILH9NSiwici7vq52I9APjb8LHy
jJ5n5fd2QXKae0mwR5Pu4J2OmjV2F7AtDxYdfpb/DEkjfMmojwpGr6xWa0sQX0bGmYkih0JFjwqn
6F9C928lm/YZiwTPk89wAClb7K1n4iBmIYCqcdFXdY1OUrfef4vOMD91RSjwcDAAOgYwkoQf3arb
3D3qXnKt3Z2QwjvX9lI/TLrk4H2OsDfAc9UCjKfxWIUTGMnOu7+cMVei1RF8zX3gPMLBQi7zFgGz
jR4j8y7E7Y0xf26D7xwQLjQ/oC/rDswqDBwc7/ikkQmW3TCSq0n4BcTdT+GooVeekQeYoXeOV2VJ
9q4VhIAfpopNL2IAeqJ8l+O014U3ZrfLI01aN6S2ZT7DkTIIZZuB7GYs7gJ2y/HoEveSmZeNIW70
tDD65945DxvhrFKxr5zB0l3R1Thx7G35NV26H8ScR1VPeQtWl17kWN5IEt+po/e/lW4Ofk+1kWci
6xCxpIQ0efTT46AAwuQ46XhNYC8cYMxhnZbT2yLVCWydhCHPtV9mCiF5jJgPuC6wYRy65blip4Wf
7L8mcg7dBRclvK53/p1mtSD2I69422PhkG2qtzTuh7oTkLTK4mOKniZWHduW5aG1JY2AReQeQPR0
hHRQQDcddIPwBDgRz6tX0kFQEZsHYa45X8Dt4khDm4t6KLumt2TKeybExT3G5i+CFR1V/5MgOElJ
CNEAVkS1Hxyw/AM27hBWNXDyCtX1VjC1h4Mub7eYUwjHY+lUtdz+t29ehZ44RVZ/lh+OPXShmNIO
9J07hPIbe45bO40wPHdbL6Ij42nC7MDUq+5gF/UgTaVWQ6+jYPaTT4N7pLIfn2HrtI+Ortt2Iupe
QKc579ZtScEdIp8/RvjUHD5YwIdR882nf54DnqoPprmvLYRI1ioO+2+pYPrDVKz1t8WifLRuiE9O
B4zUxn+ihn6fEOuf75gLG66P8bIkOhIhxixjPh7VMD4tgLmgaz+DMdutrl6pnemWdzhMcJLC/cc2
Vf7RvuTzmZrlZR76fJLbNajt2WDuOcQnhsNhagJEov8U6djJqiixhgC/7Vuot8hdqUUKBwhlk9c8
El+ipQmkAK9Fj/0MGQb7j7+ZHvwz882amPvCTyG++bkpRH/gUogC/X91lmQ3SA8rbjvYLvyKStFB
48GBcmPM39DALj4/nv73+6RdPqC5reklxzgjXBm8j45yIgi/vTHE+gJPx/623UliDov95Xas7Kcv
HGLR3KOYkGSCqFgj0Ig7tSJL8xnbOS49+9tUxdMYrh3d/u2NnNtxtbAZEdTeesaggmHMQalBQ0uB
B3zclA+qHPw2lj5w/BjphFQ1LbGCqn20yv52pzLylAxkb/5pEFkvcuxqKYm+RrzzDyMJuP7bfkJc
xz+ORYSYwdZSdaS0UFuai8GSSIKCo80UTZl6KOjwrvgsRib7sQYi5Bo2Mk5qu7Nto0RrLNPYF85Z
8cfsWV18KFYTwW7NJ//Ssr5S6K6/FsD3THIs/A9xR9DhQ25S2O60iE7BGkfAnVoWP7yZ1aDnebkD
VNv7NgFOcM+O+Tz8pYhi6DgC8RSpEew6B0Ib22IKa/opQcm/a6YVbUh7Ryfp4LrTFyBlfTM+HUny
Ir4SiButLcnbEdVZza+3DNZmdyz8J5lfXDQHeFvTm0//1sZf+vYxu1vKdgKbh22AtNLLtgF+MQiM
dggf1L4dE4gEXB6pD5FSuEBWxLenTlT22bfQu/N86fIfB33f/I5YROzundAtlhxfEjC9LwShWWWA
Zng4kYemnZyQsrZvzQ9Nugz+auJUo8GJRKhIkvFH9GjhVViHU4fuhxWptLVDkxXyYSqPbdAfpRsl
VYuSFi1aJtIR3n9yL4LJ4lh+EF/3cgCrNDcEWGCvQ4bD47ghIG/ry89n4ufgmIyCLKrkNh/2/9lf
Es6nFIX7igw2zUpnLQ3I+w6D+hwOAyIY+U2V3qMxciWCMHoSS8KsDBaExoqnva1uuIAx+2leQe42
G2kDPtnvC/ksNd+/II6MyzIumX5eUfX2PD7eoRMFDqrivWVrZDhCMu7Z9lccClcB2DYxpKd4pXHQ
jTy+JAzliW03SoyzSBsidJG+YDwOsw+3Vq5eeoNcIHYl+rCgcNspKDsyN5SjMhLnoxXY6g3IdOIy
YpwinvYJrWp1eCs1hj/6jSVjQ8piTqd5FjTjoThVvMvUmvEx1N+Ss2d4QApoLJn1V/DjF1+4pxDO
cBYF+7UxmroTJJk0NvAP5pBMbwfl7V8awbI6Oca4AN+RPthQFieh3i8VKq8q7UwOHGq+V5FfULLl
llvwlKM/gZmVPuKbPckUpX86RwAVond8c/4lBIfwwmy2r980XbP487ua8XnOova5efKimZtCRMis
c1VEF691fJaZQZPHavI6VstF1bbULrrTZfFqw7iLMwtqxc1+g4+60YjDlTkvvGpajFm3Wyk83vvU
8aVKUJLTqVNPJJgGL0lSuNe+9Cjia7MCBVP0NJpb7vbglpb44+tfgPwNymx8C0YhS/9RTsBawlCm
4l2sKW0Lq7kjFs9YpBqR2tvbBX2lLYyAT9H3teE8HhVd6FzaJi1a0h55VbyQvgbk+agGlVaPj71d
Y16pASzHOf266WIdQKYhP1G39SKgeM00BGkbu6MlFZDaMovXli84n4sOuvpL2iCheesVYP5YRoeH
3qlS+WnGYupV4MPB1nsHO5CFaC3si/YoUC6AlCCyH5nkbO7t9A+ldpF+/7tz+XAWeLZcRgChZuJ5
GoTbzo6AbYJoKVtK0qgUat0ekx/S1Yloj4FTzaDHlERxQKCBEHKJ4iOOxaK5oRnORz68j9RWshih
9RtkWDipt0OPQ2ueoB8d6y1AcPh74eKRJKVINU6R7YwJ7ekwJXIqMOwd6WUfQDQivQYWps3f90aA
zRPhUuRkFNdQ7ScMyiA8pQfpaF3qsXw35FVYkANgZH4iEkKs79JK4vwst8hcfJCm5mou0uSQJNn+
WgKAtjzjodn2TieiZ77Uf8ALYoi6pKvfUTMHYGgAZEFxRTk1z43zJR6Pe7hCiAjNUUvEIfDk7PyR
wrPN+bHkd6L12ga8S/24iWzbEwmnSqWND0sCNsYPNjp1dpcf8XIvtNS30nfJYCvoY/7Hs7MJalN+
T9AHNdJkZs25QpFIVJ3a3DhIe5lPosR2Bp/giuNmqSn3flK3VFjF2o3MVrHXGSPraN9aUdtCCpDL
ymBEwqSjNxW1WALmlbvfwn6OH1QWtNLoYvbSW4MA0xhVTvF1ir39HG/ES+2HwA+fM6wYMxRm1IK7
ITkdri7f0SurSwlcMsLMhEa+81GLiYYMOfE1RCWunxAkgXdMxrzj26zO98ZaVjbHWkUbWMNGGcBV
5KpV6vlrkPYsbxPcONkfXkgMnejzYly2SdLm7wQANmEa/xOvH+AeImc7x8Lx+u+siG17shkVmY+2
CW8NS+UwfMkBoJBCe/LgvCpIHu9OoUvaChEO9C6UMnkOPqfz2YYgD7Fjz6s5HGjs1XY2HGwep3/k
Z7ECx5WyzHv15J9Xsw86atUqZUBGGgVGBmIJ9sPJ0TJ6NsllI7Cz/RHRjRD3jl2nBeBl5JNdsYQv
VTy/pBndscyqx9eiWECt52OmomN3BLZlude1s43B65NtKgmVcs6hh3LLLZj2aSC4/XbBc+u3/ReW
bY5NN1fiuTopkqGC73lBX6pCg3YA1PtJXj5CUjDXcDzzzcDAtXwIIAOHxDN3HS5+ASXeDBuTMgdM
XtrXvu3n3GpfN0B3EKXniVm7fvdqHl5nS3EnbBBR5/MM/5cQCdB4sqAUYAWeui/syvR0+0a0f8Ww
NBRaqxY7ajgM64Ueyie2hnzAq8DNibyQngjEy//RUXnci8XDAbtMaVdZl4JvQBaqDNZZei2w+LtI
vbYm94nZuwJboOSOZBw1v5gNzIi0GgfW902Y+E/7+L3kLUnItyv1tK067SsJKNfEC/nV0jqj8Y/R
mwZ+SYY4aVNLUwae8/D4sOANnSM8ngamLFRPNl/iCyZZeYFkRek1gB7OsKjCiRl2cLz8dyXR+JKW
LLZsI97FUP/Oyd4Ya2hWHP4SYZwOwaGCvJk/F/S8wMp790Pt0pS0ydABr2/2nZyWiJ89ZHFF7qN0
IDXYlC4dbte3HuISb+t7Fc9evDOiSaZkEzmSaDr3/i4UZlhRSDx7ZgKE8y+gT/r6ot4i/q8EV3xl
4mkEbORtfd2wBBD5OR8vs9YTTFB4UpDkd95oXmI2ArhqoWZ6glmxn+pDfISJr0IwpqtfoqfjI/ZD
wXiemizH2484KrVRu5dmrV6Xa/XsY8KYeFiYeeW8EGesooKeOSu8jr2VB9eLT/bhzmk9RDvhs1Ri
UtDKCS8L9smThck9mvcrZ458uLfE6ed4CVpZNqZWtgprTfM9OVg2uLCIL2Dl4rhF5udVmSSb3bXM
YMV92Il3x832gT8pTIrxaiyil+SoKrauS7RDRMfE0GkfpW59cNxmiAVkVXu2LsZyoolgmFOQh0ze
sSSyPpmOYNS9UuML1TDsH66lif0mUvBGU9954HxIi5imtYAxGeHq45F6wEXaksUiF/QtiiVmF0kS
ECzDPi4ZFmHZiws4B/iasM5M86Fz0T5AkXBt+jt4fRMjEue33lUaI5q9dEriIJ0xpsY1MeYXN0W2
HGeRynb5MLZCTpTlf8L2+sGGyHwtwXFEnuX1bFq6dpeWS2F6rpGdwuKTCz10JcuLvGCTNgLbTW9p
HdwBFkGbMgmVRL//T2AE8CPDXsBrni0rbB17bd/mNRgeUhzN4owNo5vF7ptSBxHvmVcd2Vj42EqV
sj22FF6Tp4tzRwkK+gx+EkS/3jQ5rlWstsKVZnLpr/jQ/n0XfgS+3N8K7EdqYkWurv4SH7UhdbZg
OxbEAf0oFKq10vdh/B6AD8t9RFBprch0wSvKA2y6HwQOFvbHUeLqV36dwJWwd+72OYCmqAy082LX
H1KVZiYjcz7Lg88lHwJZ9g40C4yvg6n0pUnFKWmWq/8qJO8fiu6FZsig4KGQHjuP9JF9JmHNRpL/
i5oOo/MEtERlzlV/6A9PJN0q41sdtmeh5g7EiN7P7+PN438RhKHSTf6eKCi2C8lFoT7rqTaI22OF
ddMkZbTrI+r1PoPOTJy+AKunrUvWH13F0nW5vuMoZHl3JV9KF16yU3bmnZi6Pqto5Br3SkMksAAh
rlIlzIJ3BdR/1roB64b0OTl1TE+N2AXSCb1oqQmkk8GXrWRL0qqTExwOJ0OYC3Hxkc1z2CjcDfIJ
2Bad9k5wiyPl4pJVNkN6dHVGVFyNeu6AA8jLZUhvBtzA2DRYcWuiWtu0Y4t6bsUIZ/8zKKFDFMjF
f/5YNX4i7ErF/R0TSxW7bShMZow+7YV7DXo+RdAg/rASzJwllwAJunJ9fUmj9BEc6h0C5ulvWY5v
fCsvf8aGGd4AOkRc+VRk2q2EHm9ttTTSwFP+N5biU1sJ56+lLzHmcrZnmAGLZrkQCeropdMa2KuW
AvT+ntiqjRDtP+zlP+lblBQRQFXtV9h2yxhWcz5/ofT67E/ZwwBewr1Z0IxQDiSzlbu+YUdrYDcJ
cryZV8Ozzv/ldWKVXdDrm5S+cytuqWVBBZTdbJ34per9T/wkwCljYAQBJzv0HK5hkyWqmQlttTSa
FOcnOnq/J1o0qQXn3V5+ABiePue3xHmaHjWhgTXeZ+oDiu7b8T3M6CJ/H01w9gvTKmkyE0c0u+GS
aXe+/MKK9WFpcw9VgEmsXr9OLVW0OLwMEPItWELCPny5uiUzJQvBvDm1Sh0aqwm71syrMxDesfPR
BDdZv5Q9Q9kt/erfeXboWdtb1BGFYF/Kb3QLpwS4TrI9p3KqAL5rEcq7o8rtPLy3eH3Ktv4mwgUY
sYIzUXkMZBhSz6tdJ3BQdUO0wonceAWK0JHLH75oSn6AEuSR/b+dmiXNiDLcIJQe5+icZblPdBET
IJ0LMot+SLOSB1gt4CFAYZwHs2Y1kOC43Sx6dazdtvB+UK+NnV7nxhiSUpXPR37fP/KjP95+5JlY
QKeomZiy+kTaiAr16BUHrJ+mb9hJqBdFe1hMcksGbDFJzQGyulX/vE7cYLuh0Q31w04WspoNZCFq
L+0CiZdfIWfb3AAOwaeuk3uaHpHT/bSoIeGn7gA48EKFWj9r3V6Cm4L4gJ/xzAFAJOkzQvVlL81O
xyZTyOm39vhQApw37A7bPAtBYjY7gKLVs+cKUK/AjhVF3y2Ci0PDP2mJrf+6OsosLJsX5Ax1qhb3
0yOmZIq3OCgfOnZ1Gm+aWM1SVVcEdcfBlPOS8U8kSvl9e5KgAxfDYZwkzxXHOGgfU7HJQylin19V
ZVUWirrm64dHCj9Oh/C4BLNxKeJBx9BzMdn1he6/cktkB5c3ugbumTicZ7FNdmSnFRDhqhIbWSw8
cokGlLAozLXDTEdmSHm3K/dkNs8eSyZMna8WC1x+YaTrbNjlQCE8+gPcr+yvtTn3iI4RZcwmrXP3
pIV2+PLHBJOMaO5eEEE1Tb/fPeHC6pQxJVi+O7ROf7yL5WMcmeqoMbF6CXFKEpqk9AxZOtJ4iaSj
pipjGWJuZDUnVzi4SYidHqtrEWekI8qBWKoxq+RO2ATw9hLECfFUA7a22yGtZj8XukCoSFk5SE4F
cu6fiacZ2wrS6E8MVJjkM4iCHPF8nwZHQvk2+av2QTUEUyr7TFuDS79pu9NqIktufs46TET6yAAg
rw10LC0XfOQ3AZPP/x5IlU3Sh1ao1chgs34n3pcUNvsRPfEA/gCYylN6KuyZsi7u1IFpNYXlHv74
n245fNa3/iZJM9xqxQbWYAd9FgeSdWMa9zSJOws43AESMgMjyhW9A73EZTw8Bv/pg9HTT7KrWvpS
WhbTpE9SGqoGIvBeJ/ZFCWuwom1pwfAy6hXQN3TFeKVmMtRVgdYfIgB4oiaROUPLusCmo3TxO3Sf
nVohyOVCtijjYsH22Q3/d7MdWGA+1ZHmGQlm2Pae1xrDRDULJvrf1xqgEo19Zfyqx0h5XwxBPiYp
f1P9RzoLu7BnY68W/aAajVyUNmBOe+8xzDEKDaUjWJg2UCTRcZPSNKk2rdH29hsPmP2IJWOKlKAN
hJ2S5XcnBUg19Hn6ujOxJvfSVQbCUZwIE/9qJPIyD4ccaTKViSHzrU1qWE+LWAquzhgcujzaY+FH
SZrk9r9KGPz/j6KpCd3NquhshiOZFmjnNgVnfvD/93cB1ARNmF7574v6G3ExdE+Pya1cHNnE86v4
Uqh+lN9k6oylJfWQHy/UhpxUob4bHKoGvZtbcU2NrZTFEyPQTBnZSj8Iy9qKQYfqm7O6cdUZ1SLU
xLuHQ26/il5dwLG1O75VmLU3qRu6W7lF8e/5WN2VCif6aOv3+7cWudcubR9dv/p4MOYSOzGUPcIU
1VPm/wZJjFZn7h0zbGjLCy8ma7Pk9/4iCgsVhZcqTKUW8Tf7E2NULIU1pcOl/7QGBLpp2/kV0rca
2YmsgPeh7MPVa54goe4aZpnw5HijKhHy9d555pdhU8i3YGQn1wycV6NoqrAXVvEJcBMGLdIbA05L
llpeV43WNvnY13jSXUGpnapVl+7dmBBhHsSLbI7vkSdnzfguFZEsQ7PH9q2/CmEj5Y+GFwAhOHgy
dhR6B5DZd1Ym1zq5/p7ShDDJy7f3FPXpp6GX/Jm+XTMgEmhaj+ABO/CpuCZGoDFHp6J+M5cJLN8+
L8KPb59eznRWNV0VPRu/rNuWwC6+kP0oIcWFrF10RyOLkkNMsoFpLlbU50iRYYpLwLJUyCIYXqui
nC/sKUQhZEE7C89dBAZo8Ygw0HP9n0B/BPhJeVV+NBnu+cElMjf18OVkGuE7AoQErRq/gzYvCHd+
CX+b0KSy+O4Inaox5R4kMGyDFLny2OPtaYRDG8oIUDl19LR5/sHhBLH6jO2mUluG0YMYfomKgacn
3/lD8r087tb+au+5THNY46OfQTfAFGfeN0T1dPKC1xrmSAvsLhRY3o8GTE+e3Rm3HMF4W5lUD4g8
YuKzb+VObck+Sv9TZ9om9Cw4rB7Wraor1I6wI5lyf/8nMJyd7GSog7mTO2Ay7HqBCbo66fN+jb5C
ItjOqy9EbCjB8gviJ5Rnd4yYy4eTTgOZ2nskPb0SzPoBbNnnUgG8FC40BAFlt60hgo4MPQzl60ln
dLC+X+TIBpK1L3T4MIgCAfSIyQte9T6PAE6x/2TJJB9R0kCllaz8QOiSfzBMAZNjmYpHqFfDI5cn
MNjsjTXPuqd+ZTcgvyd3EE2YUy+c5eEhY6EsdKEJvoy4rmyZQTmvD8B4O3OyUdFJuhKro25g3Udq
dpVbKQMWVW3xIyQbmvwNvSxVofPCTqW+Vxmh6/fD5TKdTZd9wTsoLme63JC1vT4uJgWf9UJY1u8X
2GslMRVLah42rNGbcYTCDYEXqbabAwAnwW2z5REUmvnPll75kTInIoAF6MbKZJUggJo2dwoCzS+3
QqkLpN2oocBFhyymOoGRgXJvPZ2BRm+LHTwQNvfL3/l2hQMeW1GYRJsYUb72UB0l6B/Vyne5Fq5q
Kn+Mb1hCFgqAc9xY9LsPRxwxikSH0ch+Vb3aVl2YwM5Tbwcm9aJVDHcQMDEaez8ukCWZODF7ERlr
IrqFfZTaGC+kFVLAksURSAIM/UnuNnZ7FHRvW2iBHWq1dLDE+4FwLkYp45KvuEbj82vgNEy52mmj
pODZBMYFTyxi5pHbnyd2jvuXhmQj/jhHd1LJ0nHJvg0H0OX4ukMF9YFNOuHXu5QrUOISpetK63UM
M/8Lu4dKsCswUkIBn5Xh6lbQYZXRBVPW/BXtUMvnVLaOtuw1cnLwWpMsCPYkzeWV1SKSAn7lDAUP
VIIrJV+xhiuxzysQ8XeOkzYCE5EOW8tcZJP/thg5JxXXeVKDGaNYospFuh3MHuL/yB6dHizFypb3
XYbAPq49C3wisAY2vSsTZgnp35vaAoBzLijwTQAqiPvGOZ/Y36ayotjvko2OoBuoUTkIslzGuFCr
s71SYhfShsQlxyS3laoEevHEpL9c4bvGSERfHkiuOQ7hd25uO5gDvKV1lMHYl3w7psRoaCqTKTWe
PVkQJIy5M9MPeJkyRLeCAGoLbT2YOAjfWvb9FYWjSXIG/hqYYUJpOlheBmDPSX4vbB1rqYCiN6DI
yHgbK89fl+Xi/gbvs3u1GB/0+OaiqA60FC7mg6CwKPEYNUSpsFKB/6uzZKDOGKbOb70uARzBbFkE
YOTLaG4JT1MCYenFvAom6+hC9Sei6LcSZNwkKpsYMfzOF08Jzph1uMzpi+xUn7RkZh9lhAWKp05o
wuD9nZ1L5nLj2cICAh00aKXmP3CZcNLld8wrS9KJUCc1g9qg3GP+KvL741inNz0Rj9XALbYw/8AK
0bDqHS8Xo3dXGatYsXw2etpPBDm6hP0zBz82yPONuhFVbmSfy4NG8Rd9Tz7nA2zQ6kO8oXuIBYCz
Ufv87HIWzgCEZ9AWFs7W9u+tpZ2TauClXznWLE6tfH+pLILqJdCuA2HV53mJmwXWVAI6W/mfU5zY
Y3HOmPcLBEDFQt85RKL8ySWycQ3BTHf2JSdsngXrEi5uhhU4FUq7Ir9inUJFErsaYtVIr4J1nrXX
x9yslgyEQLs+K7p55C+iU2D0ya3rtFpPtnf9VegvaAixiOEbAvv+S9iXUsuLWt4ySrp/tLDg0Xwc
Zo99Xa3XKsP3SOekwoxL9O+Fv1z/5D35EwRyt7F98LGsPfCQfeIc5A5gNnVH0A3vZXkwvKogE5vx
FESLdi1t0hMsec5+liNyCeKfVPIAf7tFlDz9LvLCBX5p46d+CQi/r4GbEOtO+16nJc+9tVztL9Fx
w22a6InlTTCabZAHtYHGy3V9aow3wCNsQk/WZRJy15Spgj5ryPjA9Rhhwj5r59J5zaKNt3t+TwuU
2y+zhLgM1oLcT0O4vATKnJg4X6/7epfXaGk17fpGj2E+pr3zoF1FUgN83ceEC5y8Mn+yC7mCvAbv
JxLewqoXfMWKmZzTYUABaku3+Z2Ms+lW5VlWpDnLL8DGYACWankFNRL1MQlmmbGE6+NkUcFWS8Kg
/8rCgc606Yl0H1SOK18tglgEOqHao8v83P+QmkAPMWPvfCuDv76lnvcRxcAvbySXbGNVgi8cQr7t
1azQdRHf66ORM02bJqmzkVjWqp66mTn6zrUJGKIQLoBMAolKUL2q+c8rH4UCXX2cv7NBnvZjv1fE
AKpWCTaFFpI4nHiHpmXz9E/kLlqmSvyYluJhcltKuvF/rHes+EyPwbFnOX7X7QfrYusMuHZr/TQG
rg4SjQcv9WzuGHBFZ+KJzhRVP0SGnfLw1wPRFoBLXrZVDmITXAVePCRh8rJa8t5VbzA12K4GIE1I
A/dMbkXjNXFp2+qsaEckQqzjrbPJ/t2vjZ8lSAkr6QaWuA6iFdMyT+mSk6EqHEYbjy5cs5f2ZYCw
8dfqpOvNaPbzugBhz2uGttq0VvRxMLyEf3gv5UOsCxxDCJtsvuGWNtHUmu9MOUu1QzJQalReBAVR
K3x1MRoYXlwiuWVk5ec5dtP97TcC9LAKTBMQdCnofEvpFuT8BPF8kCO7QcjxHEuTLM3dBepkf9uK
GlMbE0s0md4XY657SpXt61RGSXedSPU/1aQ+wjKc6ar8e+bbIDG/cpcuY9dK6tqYhELwI4RlTjRH
7a++XIHZcmPOFB6k9QEUT9270V42Zp5EUpftF1g0kai6NkIv/WkwgysaWgfKxcDqs3zzJBeHs8/T
IGnQoC5WHqfEMwD+U03P8Gav40qrsbt4i5KWwOKsh5qx6H3aZjT8kk0JHaY+ueMLBZuyP6xdoSRM
nuFPazuR+cjqVaGYDTB7ZhwXD0EqzrwsJy1ZgAT/p7nW+/XYl+os1ivwjyY5rWJnjbTL7+SBfLqM
FR2iE9kPhnarh3WBOH79EMwjW/YY+EfvYHo145PTXPTJS9cSuGpc70OP+a1lugL8MDKrejFPPk81
f9k3PecvLb7wSiEfOc9Y7/9U+uEvNfonkNZbuMxRgre9wfLim1zGE+muir66oQg1eg/K2exs2+s0
146xMaeKNsGQzJXu1Zr/uDTBDpT3MqOFWXy0BZtzLddwyGCUMSujhDlMm2g57iC+2PjdPqglprJH
skZl80K8qD9T+UHzOKN6gPibBnItTlPEs+VUUlRBO1PW2/Eq3Ls1WXxjI6JWskNxE9FA6aiq7YE9
6eNEAa54EHGUrUQjeFyCnJlQGIhSg9WYA26qCcx6Y3Dv5vOgZxAfXlChJSNSaFg11A4NE+cHjtcO
OkFQ/bOgC7ypJhIbdi4RXBFXZ409/CA1fa9m3o63jLoXhnC9sTmwnKbmMkEce9O7n4ZVceVbJNHs
I35lK1TQADwQAeltc2WoqoJkn/FKQ2wNhL7971CoQhYg6xI9UZOeuwMnKOGoZRnTrjQMCgIvQncK
JyFgqbo1YJ6jVaOtmgiYfuTZKa2tc5ZDmh9cNfWREKtjwJDPrlEHyW6jFpN4wi8dwRzKG6hgLsfx
SRPMuEF2DzReK/hiiD4P04KJpO8Rit1BkqBuS9NRXkanpQy5wFsvc1Zh0Zhpv4fwERF2za+H5I4p
tFeAAC7aQVl7aNOV5YoNg6vba6ISg9pDd6Qjfh5xLQd6iyTcwUzPzzjLLGExRGMRCsr4qdjEdizF
IaAi3Nq+L8NypEkq+6USKoDrj0LYdrsJMdWNvsNl2H+hQ2sbIPZH2M8nMOBGr18m5JciGLIw/AuD
QATGGrtsx1xEQUYX3X6HzCVPBpeR35QJ7Nv5QGnkPCrOdgWL4QanIoYdBbllVP8bb7caE6pPsErm
zVzflAJGnDOGyuifPpIoJI8GCny4otWFP+ZsyL3GOTp9T6rGmBl7wfSCbpDqzJPbV79DVW8JPSG1
gRcd+cMnImMi4we6r7T9jSnIPZYE+UMCC00KoVWKOKY2ThD1lsCVIhr9NgcldzRVK0k2uhv4+R9c
kwrgxNCTVrEtVxWkZNjBITSLCjEgruYRZ7PkdCsCQXedmjoovZ037BhnTl2eQ3eYkJ51BT6fVQpP
vtFm0XQqYFbIsfKq/NQZOaKJSK3/Y7WL+tlsCmOChJGKhFH+tFL0CwNWpZoHol5ZUDLdrmA3GI9G
ZpoKTppHON3s0/iIL+FGuhm4wyDw6KWYqQ0sYSO08PF7hcxpXIMWYM3CRqLkdx4SXQtLzq9xUOXI
NQXIPmA9UkzX879fTMe3MQmUrC4TK9bmzQtRnj86waIrtyh6uzkO8KsVJOpWcrQ+PDIa2TFGjWlj
y01Sd7f+GE0WoCB2jeOX0U365VElyyCKj80LsecOhNKdEySAHThLXXdMp/2IYg0KxTkXT6XtyFr5
FF9mcjmS9aT8mdEeBV+dkAuHXRa3VYNoIgM58vW04pgrnR5KopwepdFLYTESvxUkqAvzVWnIeEcv
yh7pUFIVwMXnoMm7vo/GWi1H0Pwx3vx7oK+DTr7kvjf6hHVKcQnMPGIahmFSZ5gwz8hofEzlCBU/
sI9y0pGZkl2npLZ61NIGpq9IhTJGEeb5fgZmgJRwW/erlSWgBxfNgNXl5Dm8MtwVmCTbgNW4CIJ+
EfUgAtuvVu46yQtg3XVSb9C4Nxaz1o6bAg3/0zyLywpJH4kgQWbrMtW/3shsvB3yN7wbUlAm/PMK
+zHEGFbgDcdaO/kKdt05FdEca4i1sM2Z7uvQ8gh7rC5XhbmiWLfaaE7+jmWI4Ao8+QcZShETJr+c
5vARjPYwzp2fTxLaubSlI8ZhrT+3/vUn3VqAG9T2h/Woh8+NFLWzyqt+GtLlRpSd7MvoQvDMQicT
BObRgzxC9ewuNxubtrMmZsh/sXeHROX0ebK8+Ikim8txzEY5SwPQiHeBSwZvsgC/UsdYXCGdd0Qk
GbPDvy3FHcVfSOI+Vq0N4t2w2G5dxelF2RMY9BfFslt9PSsNneirhfgDPLG0Y/fe5LT32onl1dYM
5+79h6Z3qsc33tIqNkw9lQeAP/iDtVU4SrCkVLRf5ynjEDu+1KY9ukepuCQ0XvKWisUhxCOQbenG
F1uiSLXXclaQVwgcRPFmG/K1rmkOsEa7EFF9RdW3njIj3+sGsAeBkOCxXsR3XfwweoCEIv6xePab
UYQyoyl9iJjzofYsxHRscP02jk3Esky5lDv0mONMbsaSJ7uE+bhYmL3+qWDpvE02fNNhVfFGN5w4
lO0oC31Zb/RAkW23Z/eXvFXBVwV+q95bfvrk5GH1WX3XzHuHvavcZwsEWLJvRXa0mSQfGixPzfDv
LQ1sTQiPl4WOPaQZO2pSFMtFF+nGGIqsL8gFDO05my8RWalwIhAMi9iNoIdHyPUqMQ3L2XtV16aY
obmNMiedfqp8CTSqAwpsRtfHS+cNr0iXsMzmMllD/sq3toVmEhDNaT/WhcuPHNuyn85mAuTkRl75
qteNjYFPvViv2p9+tvgYmbBhMhJxAgYyohnL6nqngdwWQZsMyPSk1PFSiFttOafXYNt/FPw0u34F
2kyYAlQa/H7cKI5v6YP78Wq0QMSbIsSiXGjMYaMgR6kxAPYaUm2WuAVjETVdK6fnA9aNZDmWfKEP
waPDFFrsLiLlpqcaSkm2ESZsG+DftfAidzJBRGRny55H92XFdHT4fLf9biJ5l2RzzwRoxhd997wS
BRmqSqh3/o2CxPffP6oz9hUtyk1tOBOc5SB+fp7DG7ZFq45FUSAhW1W/C5rd4PRVAT1x72b5arbq
vWb1vUD20VImPgplPaW9gvXsxWDIf51SwO2U88JKsCrIlAddcpS+Q2Jk4JhcjcEeAEMPDLdcoLsz
6KnoDd6ijGXfnmUgIlqZU2W4k2d8A2+rIkIUkYGdDrhCm+eWmRJRpyxD04yRX2wVNCnCQE320Nio
1JQdRBZbbKbq9ib5U2TzCmzoyGS7wYgGCMMdfa8BiaP1osgEGujeg7L2N4vel8fI/dzHSEnr8QjA
N1YjOK+oYk/Cxmw9LLqciDQyDqljqGKG/rQJpS/DMex0ofvC6Q7NBixbPEjeW5KXFRYaeDxBJgev
qvBTaf14aozZM/i0FXAXVcmTKgsoHQFaXXDKusKn1PQY+DI51s4TtB7Rjo3gZjExMIzh1V21LMoM
rZpFFr4vEMOCyBg/+irC/k446ZdNT3mub89CvXpVHhBwpmAQIYVuJMbX9B/fJ28agBFApDiYcOSQ
JUwoCt5Xfvmc3/AgStKI4+OJ/nuwsXP3romlKKBhL3n0QH/Iu5wK9vLOdKF9j3KXxYIW2lwBtOR1
jl6xFPMbZkbs4rJ05ujxvLvCwYkMrWGjHS3Mat+64S3qTuh6bJZIKHYNObHQ8NOFP8kQv1dwvGaH
tgC5WxY1qjJoVaHMIpv5IcXVrMyDzP751542FilIdnuhTSWm0W2Wohn/DtlCyR9CsjBD4yPpXJRo
ncop6qzPFVJ5JsqbLS48v64K6wwvKKcqY9FFsrI41afcFcq+ikil/b4PP/yzRKj5w/Hyo4Gpq+Tv
n5+qFjdNREJ8UDylcAXVBnffLkIP6r0RhHGlyKmDF0FRG15CZVixEpUIRfuesTVRbPpycqQE5pKG
xDx8LMrC8Y5BLtG/3yPydxuvg7CGcEaC3/fttrqqjVAXBKoMPAnR7ZQs4XMEHnUSR9kg/lkCCUVe
hC9zSBmL1RykKPuP3lRqRz9LTOhmmlJ7DuPWnFBx3LeIQkIyYQIvStTWbfxkfUEfLwPekf2ZnL0E
tqtL/pdoqmUS4sCY0oYvFtkd5ScOu9Szwp6ZBLERR3ovFK/62S3tVRKbbptTYYWLhRgFt9u5MBsz
3fG333lCTC0U+JKnZWZVe/dqfrhFe51kWLPbpivGri6VmvD8ZB5ufrLY0NjpobAZ3+S8yJ8A8UjL
1pawZxEtG7kqrBTvgqQVXicNmKH9rB/yXrqh+mIiHu5+AY+83ejAzVop8fPLkjirqqr0YLRWBRZM
zwR3d8oWm/CHdEZkGx1Umi36FQgQ7Xw89yzx2fxlmHUYpeX7T1O8kSO4ia3z0OGfh7S+jQRWuklu
m0ULee5IAlyvyFAKTcJxfezIIYJpBFxd1KPU1Ji4BbGf8mj361d7t0/UKl6Cp/RAs3ukeu8NzSyc
I8hu0oxT6rrZmEbsXfPOhzAcIAjdlcPTFbgNyn0sgnonfCnY0d0E0soUeOmz4MC3Y6OKsWOWozh6
4Ry1uCft8RqH7fz0KO5idwueYOg3a1UxU8TbHaFehO7LKVWxGWcmEVnv+zZzrN/msBuGMqO4Jt8k
INea80HYqu+N8Jx/oLQqbCDYbhcmp5Pd6FSLK8P43LHlFSai42NUtMnwTRsh9r75I3NXIsSpDz7Y
ee5stYIjzQuB06eAiR1Z329cvDIVAh+TW4smk9vtACKqAjIeMDQOMFSkiUQ2c9HZ8A3VaAQaTA+U
LIeyH3yfzrDFbdoR5MI8xl6uAY1zPt8RE6YBrnc1smYWhVWxI7E2H9jX2xBIiTyXb2ZrSNR2t+Gm
3wIgomc3/wqDytfYlLVmS61CEPwwCKpt41WdBuIsmMb/R8wlxzvo2/k1+rIusOemmaNAMD2S/CK3
2MZuWqx9osKAZzk1ZWK0o0sXxj68s+1LGZ7ViFd9FeuN7qDgnFnPU1qhH5vqQCRaAsUn2HKKhnid
qIgEIhy+fHBrsMoxIKL1WbFCAgXgCNvYvRAWwTIEAdwf3uyEuNoi2KqzDAcaDqKKmZ+76PeNDuXs
JayEcVx67hmSf3K2Hc/gohLrZtmwJ9fEXojP7eHT/MUAdm7zRJrhqQzyM6g5kISm9WqG46LKCISs
Xtv+k7Othp+DmpN6I0YX6UahgkGp23AwcbDx34O8THjPMALlyB6duK8WY96gAbPKk6V5Z3zv4Ohm
CgcIdkrXFjT88i6t2uOdnNSUDs31VUcYbzdyJjN+l+gnYxJLfPBw67mTdtpIbpz5KENL/fqQeiK2
+1f/45pFdJBNj93w+h0SGF27P+ZEEZi/yVyfq3/zDOzTgIQO6n5JV1hyDTUwIUYYrZWB5ube/o8u
SUy0dpYeGmpPz8CdG69wF0VE/0yQZGbhp4Z11e9GkzcA9FP8TFlYRmz5lRmWBeQ1e+TCDbX/7USw
iO41HNT4a62ePpw0yUCRv/B4wXYRa0X+d0WfdUybFEDmYmYMtuPz5vVnMYcdQEXRxh/pOEM52Zsd
/53mFgvvyH9h5noUHFRDWuLT83wIwqwOlOzTi4gTayIv0tU4JT/7uCS6TWkmuwAxGYdO2CPmoiNC
cUbt3NcFxwc0TvSyRYoonrQ0jWL9k4YWPOi2s3TAogHXQLQAVCY/XKsdxbbynR1J+EPbjV3qFMRq
xQNsfUVXWn2LsmvNVuSlGf4RPu10p4/gitcdfsrWZDSzeDtFI/HtJnW7JCzf1nUX1/aUnn2eWe1d
FfLD5dPHv11t+e5tsiQA5NxSsbmztJNwnWq+YrLf5iulznWKW/ouRFgLRANTzvljbEq34sYpeXM5
8W5LUpxRbQIYhbalkIjp/v6BOOIYiunvLaaCJ7jCSfyF7qMvNDl1wsjZ530MD3P/kY9X6oAl0DOD
43nYO7/Ad89/xpOiAwkA6xHMvJzResEnPVDcQ5oj0f7BtT6zZrrNuhYjYrTO0DPA47Xa5++Uc1Sk
TEesi41xyXvHOgTmf+iexviJr6cQR5xyEMKIH7h5SogAxPk5X0GbbS36TF8i46v8r7RXGvPTICZq
uUU33z/q7O0rWoJqimJPTDBCkGB0n80mf8siRsDg7tx0MuVc0nV+Vu/XiQNcSj6UZ2QY8lixKDtO
tvIacRE5vAbbQBofsAT3iE+bwp3ulvTqPU309ivln/nBr6fioEP2I9tQ15KSlI0u/+LrlV5eXnhy
LZpSDXfDGEtnoPBbu9YKi0dzpMmE7+2971QOodZjsulErPu3LHa0AGDdVnXzwDZhAjm/bSqTRI9B
Pc6UTe++3imKSRw5Ej+liHNdr/4vFF62JVI7zWIioOrP4VhD+Udr4dZMFcA7E3/JUo9y3wR981eh
vjye/AnD6ZDLQ4phK4ZVYIUSAh3HpVqM/eGUegQhQ/Yq2Qb6KsNTaoqrfN2sVRNweV9i8z1CiYRc
ejFbeXxtEITkan3m1uiYRNXksxqpiJrLvEt4J7QWj+XNHIJ7UZdqPqqAGnJiRNMn5p5bilx2JGgE
VNAyLSdrPJS3OyGwJFu8czg6AP5AV27BSHUvQ451zU4MzWvLQPdzbOMakqg2yiMks5eScUZnpWok
9r1M069z7Qke31ZQ8cpunTs+TR7oWPap655rn23QLhv4OcsGDdoO+k+eaSAC5io4CChNUHxNlIk8
WqQ28NL44+bx+SiH6CFECw4KoT4fciPT2qHMMzgnT/0MqSfnLw+xhU1P2k8L50k6rEjcNeOMwwu+
QVStDruSBj0KD1YtzOvNCgq1YvjaQkIj5I+FCVv5q3bi/a3ppmC0NKIDg4H5wE8952WlCJkxGluD
hI08yQVMlTO/LFVXmcKZPzxBgt1KXpF2WrlZISQ/TP+7OXf7o/4IMDaoo+JroefHNdX4m6RI8BNZ
2Qfz2vx2lpzdoIJpOWROMCrOtIM8fENR3xVvttaJ/Se7QD096yHU3JUez8DpNSi+16Zth27W5t1I
hlNCfhPbQFBWh2pqZfMOZRfqBi4ppWrcuCYy+eCYXTdchPheVA1hPo/oyWmDXLhm0Ul2GVScyfQI
Zy77k0Dg5DAjh5htYcUGNft8ZFcTPsGS7S7/jCkD5mDypsPIVROYOIr93ml/yz02CdvSiP/bgjN3
Vo3VoUJ1JTiG8B7wK8c8b1P+QXYmpf6BUvwDnJI5Wt4UCC14V4QxN6vqyXDlG0mN8pu4Mn6VIHnT
/Jx0H9dOvtFtYrNcQxLw3xEZ/yFspGjIBv+SILj9ZiJ/90+V8tsupb4cAnWb0gdZqMF02YojXyL3
ZJh5I7paxYX+hez8Po7itNz0pWX8OiOC4OI3euZfrY7bryXImatN2+bp8urvzE0e/oovr1wLmtjv
UW9L7rYS5st1Up+vN03eS15PcXrX8ibemQutY8T5HBzixNQX2peWglobrgD6UGYHGQr7SmTz1nH7
JWizvvBjq20vr7AtngJrzFG2nz8kbWAMvABbCxm0AxBHdqiqsBuOJ9aC2bwKwtb1XrTTrisS7qS5
HXMBWPxE5shCHtFulpCmKr2PC4ovx783KhGK8IV/ViBilA1QacH1qyiugYPRmsNuFapVcYU9dVsx
+3mGzv1/sjsTjKQ5gR7G9j1kV3H4K5ML7BwjnL4WpobrTO+SiEMpqINfQMGm8/JL4N7y0+LQHNr0
N2TxCuYkfakAuCAwDpE6O0XJHnubo8YQa3e6UcK+6cVEKBXj6R0N+nOdACXDTlTxgkCORGQp/Aa5
kGAe54elhM0msd0KRkPKrB513r7C9i9kTkY2bG8Tf7zc3L3KFdCMPShRmSEB1UefjolJEnrvGx18
84ZctHHxtST+OsmwBrXgx0UXN+qTiJ9byxTnETNn0mOSPpl19StUmLwRLR3IIqlzKGoizaXqHYgJ
2Ow0Fnhc2mON3o1eGU8LdW3FTI0V341Aq58YC+mbAwofaWfmjOw1vFEhpcAlGisjM/QvApiZCsRr
otQCRIOdwRmcGqE9c4hmAR0mU3Ck1ei3eoWC+eUCFSOLpmSdep3VlqqCNdW/oe5Y01785MUW5AXR
bbIxdhiqzrNnXPbXvfburGFuDT8/PNb7solUBsLdRGI+uOTrWG15kt7leBowTexPTunZyXdF4sBp
H/HYnqh8zRnLf/97lDO/XwQxPhpYO8/0cICwXx+Lev0DD1lx/yCLE8o/GlDsMqssEP4gc+62tTHY
46Pl7R5d+wMctSn6l3lNhgeKRki1bRERSdWu77/0yC/vsc1fvH2iBN31o4ZfUGUKiR8UWkIhb+xX
zy+4JcS70+M5KVBC03YwCsYXAAtebwdmSrye59Ifu193Rx8Rw8KYsxTxODiFOB+WDB30IZlZs7Cs
JjrS2zYA1z8Kau8NqzEmpRTFbedUps+3nx7lr3VRzkdFfVmAWb89xAc27XehbZWpXKET/rrdBDXl
OR+Tspn+m/pwgPqHvXKiThMV0zVYkEg4UK1mDVhcv0cGFvkLlKAgkO41rFT+DZwL/XPU1DfjWYDB
X02fSTPVMz0hdnN7mXVowY6mkGe6tccp/AmN0XznQEbsP2Yzll5kyWao+nzZB6jvYLK2lTOqCFgd
A0avCI8VGPSyQO6p9661HlcECvs2YmA0dyC7jSFDsKXLcN/ZyjvTH9DqWCc1Z56a7TP5ZN5ebEp5
iIa3oxOnIhZZsFaTFp7GaXta6hjeG/XqI6VYsKTgtqd0yO/mNIKMzYcD9HT9eu3YuldD5cS9o7Rq
K63Y2JJ8dKfBL/w8CacnrvtJBtMbW0Z4No3YbYUCfMoVXWcNtdszKUKu3U/uU9AP/bFuW53PBhM7
eUSuPESZCGLXh+Ecirn0eMUfKZpmkM4hRCP4NpClJeNo44NXLrfNYEqumAhTBjgyN6EvtbtZJSId
WQBLUpThjIoRTUg5DNIfbszp/BKBfIPLvKJRku7OuBs5/dZ54NuQjXTfI8SXu7fAQgZVgTxLwNRX
b9IhslVzT4sSYpF2ZAjrIw+FYavjmSJGXMwQdmjIhe7LHPX4P9ob7e3TzuTH3/+P1t3Kjq0HlaLk
84WHeKxeK+ViEMZ2CreQBhCVocHirVoO7cChgtPlp6u3FMieS7dvQyk4Udm/htNMoLuDip+dv38L
2H66KXMY6lqHPFabPml4TrwKsXzsFb1vailAdElfk9rI83CrY5ir0ZADc01qaOTGC30X7PWk+DYO
oObRyuiIzHwOffbAX+7R0NZnDB9OFgqNb5YofTPX8I2bIl/tpIRQ2ZoKChBTUHZAry3cNKfsLoII
tq7+soP0IEap1aULfymgRr5jmizRs8buWOJl/5zZRzjM089za91IxrFTrYiYuWRLDNMAJ/G3EH/E
gz6ZKdcdw1ELFdYfPq6Xeu3iiRIjSH/JLbpyiGGhbFsocamzk8QnHS9LDvZe0bHukasvI4rqzgjq
gbDMaTll9/wYU8++wYnl3kXcT2kzMOGZ7oViCrxIJASWkVrKo0Iwzb8Dy/IIvPpe/GQrf5V6FAIJ
MLbYQnvfeEY5QksW7/AQVgNTWwa4R89fUovdJIAMudI+xl/sVC5Ivs5TeSYkrbCMeAMXOuXic79n
AfyJTNIO3GAwnwANx/AKOH5GUGGvbbMfbmzgFlIqKiom00dIzehCrEB2bOrxc9d9ZUenSDb8QNOr
DqJTUCVQ6Wfyee7QBtd6EtFaV8BBSx0QzdVStnpsWRIRTznKLVZmJmu5sF/cS2NcJEE7TfEr7DjE
g+7FYR5bm7keVaERr7m5F+wP4hOXEwGStliK8XCL7mPeZZe+hf/LaxqXHOjobHfGBmN5JuwmRPHT
GA2pecXyoF8sW5nRCRK6E8cmNXYd3sZqy4o4gXwEsYsepMWcdVuoPieL4/HqW0QR8+MerwzafcrX
J5HsAjGfX783nfAr5bxsf1+D2OM30ziaWX+m0vvc31V+bzp5nS9vvK3MmGby2nrj4fLrtkA/LtzE
BZ7JxpFRfOQauGWqiYxgo6yMAS0eVB3VeMgnaUkJKrGwnUb9CgmatS3wdUR979jUlWfX8X2lxYxC
AOpoZ1k+0GUiIlpo8yuIHqhtww0JAQ8Pu+40t89xZtBaeaWLz2YBaX9b8IP23teOuxyakh0t5Sr+
wk9vntJEHYBfKyRVGUjRPMUyJnsq+J3MhwwHuMRUsQ5YpoQ8dHxtp/S2HOphsjaFDAGDwg4vFVCM
+L5P0Xs3TFNRJ6wkr7jiO0Tg3FAbXAJFu+1fdHo1d4EPofbLxsYhUbUNcktgVoNVlH0Qvwd/SDow
IKpD3tYmyerKwIECAVoXX7pXp2EQzooQ8EZmvD02XxvK/D6q8AZqW61cB9qBES+WDWylIQOd8hJ5
YBmFw0QeH7xfWGlJaRcC4zzKkuwyRqK6i2BZRUinUcHVVVHQNgMrt1MmzdIXm5v1kroi6lRhZcl2
t5llMu0ullzLmTiYARMYYXe2fGXahtT0ud7ZAURm9IPNuM1VMhRGTVM1sTEGLrKy9qZdBGaV9eF3
4bBGeWjx6cR0uuc8iK4z/A299kGZWn2Oixk5bGSpF38aoqc0Z5NVqVmLvOmItxxxtTO6tPeh6VXm
9v1Nk9zrMwoYlgZs979eTdAKFEGoQjFRbCprESWjBofse05quR8veIVvS3/rkw4JhfFNUIfnX35D
RiHVYxd3Undurpql3mOMYOFvghEDTEawW5lgMJf5Myj748yy1hgMQ50Uq+DilmE1+Y1oWHpQTBHa
v84Ck7l1R5FuMZd3WnqQGgc8T5ee/ncj5wJwK6sS5GXVQ4FqyOzkSHbif9Zy29Qvy/W7htnFnXOi
S/+whgOZ0XnzYB9Xo3OAk7HtuQwtJxo4ZemuZLm7/o1yG/QrhS/PxQbThyvECYgS6fXoAzLBfBGF
v/KkCx+lOv2UE59fgK+nqxyAFQn+uglchD6rUDxyB1nUHQA/RtnGD6Ag3V/PETueGyh2XH9lsjgy
qIKCk6s+Ko03LWYyRwG8cJrPvQknmz2zjV0zowA6kk2FOSC8oItBKHvCX/oyt/jLC5te1zJnOu8k
DB6C4/wnOQEQeTBfp4tTfNzvGc7KIq/M6qb2+hMfVAJlwGU5BKx6x270wiAL+yulxfyLf/oALotE
4XLABlqm5uf51Taamys638psPI42EhDDyFfoZ0o4LnPqUQET9gxQ2pu96mjdYI3uIGJyd+y9zvbE
4m5yMhESewA/Y9KSq8LmtdtD25j58F/pYheEAh3FS7sbVZQakgQfA2A/XBVu/nRsezfkqkrpSdGN
1jQia8kh3MpxfrkHrcMmRlBcoN7MrYPvXcPco7Qum0i6zKjeaWhSsbSrFE/OZjicPD148MgYXkK1
tNBloODErlJ6VdySW5hR+R+Vt17446qm4Qu31XlL+vKR66wvxxVX38Ys8WXqxkJKKerrTxOEY6Tj
DHI61C896xQxaeoibJSlI/SulcSHY1CmmefyVhgltkPa7sLaaKPQDjFDF8tAw998T1aeTQWrh01/
pu+gC+/zPA/M607AOzJD4ZFY/cHml5cb4JkJ+F3/MGGEUOGmFrRJdSVPvxrcEvh+J0KzDEJrtx1W
8XfRs4pN7SNS1HwunbqHEq1355VfDtdP8V8fqs5G1RktE0NlQoPfIoFlpXuHXlE2hPNXKK3Kfkxa
ElIOH9SlWO7dhEqXi5j5SmD56pbzBRsTIlcfC//hE8vynrjGPx3jTkqtgGxffhf+mdPI+iL3IZiP
wAap66xFysCvfnaoMnch0kG8yhXOoSGxmzWywYJjMNqmLnRBWlj5+xmhLd7r1eOnbN84hDUTDdEC
WSPIRdI+Q6erbDHk5LzyL5fihFhaJml4rZm3lfMKOemPMcJPavOd/hPT5zD7S4QSzZT/mAx7HD2y
/touPLH7WykUQ+UcphnXgugBEv/hQLVYWuVgQ0FOk0TjcqIuWhgb0bfHMIPnlyAtZyYTY9qxoCTM
+vaUAqUcb5Kxs9suRivBYNOWAfdgrgaKiAKk2Rwf7z8MdWtA6+sMcFxmzmZ3Gau8eCrNK9rBdzYV
thmrafmUcR1yAPs+bIa7cHDGEm9070KTai9a0YEYBqIs4uzvrpn4pIoTvQH5HKYE+22fgg6dv7A9
eCZNjKUgbWAG4MqG5zUhUnGl442dI8qn73+DJ3IdMw5MXGxlHzP4JX85nL7pdvr09Zvbq/3XAk5/
7WunVo5VgW0BQ545CLQc1QaswyW7Zmf5flFk4HFhjcvWctMBczaYNakJX6KABGRp8F6HbcYN1FsY
VTw4R4EzVRaWZD358dwSCk/Rrk/Z1vQHBmjioQF1d6Ee29kiIU2JMEDS51C6kWE64ScDORHHb8u2
pyEtWkvcJmfrW1KoDQ4v6qkcIoz7X8cFg5gAgGrtXVVHrT96tEJGjUIz2Hhcg6uDH6UqINbYvtyg
17KyD/QCrcHWjjrdn4ZKZj7cSIW3r0YhEaQFnO9kt8vsLJ0fcQtwBbzQ6AE1bDphni/zM9/wRJV7
MZS5jUxg+XJfrf/1F14Xq+nqxxSY41ICi57YTwkFNPaqpUKmOy8RzBOxX67g22s4MWTpZRbcw0M1
BtqE6nnBjsRmd1JR0fiwShbQNByqFqgWwmqnmlu7q9gMFvhSX2XNTt+JlR2HZbHA+7Iw+xsstFiB
hgE7i8ghwWu7GWq+ZxTxsXrOrO/C56alxKuXhZQm8f3ovMUkZv6DK4aTrIA6Y2IHqM+ygmZXg2p+
95IePzEzSSKGtjO2vol6nSh2pqQt25h2Bga0BKtDSeqDpdvwiqzqAi9yRvZ33qIyCUuZaSPaZcm2
Ap61wKLdO7ikeEszH8WHJaTns5JdTY7HvZlwR/nBAX/UkVnl5hnA9VnyPsmyEKSvgACVC4a6uBdH
M98o2AsyyzpRoLXzLjjR4EqZdZ3eGXsMXtdG39h8FQHLjT9F/rjom0kxZ+gf66hlrtP+OLiALQhc
AqMaHI7ftHqOnTegwDbhj+EPmIfGwBdPuuxfBSQ6+NddB2/PsGVQgq04uTLPlHOAsyFdvAUUGd7t
jVyu9M3Fp1+ucOEweQ27bOmHyfNnD9AOiIHYFglTU1qSeeg70HqpCIjsJsFk3ep+3b8hx4blobLj
Cje8TYXfAXnw5O8zJeUJvvF0SoYXFRjiDjK/gzjUgkRT4xNTns/dfN04LKLL833rD6DWtiins19I
lBRk4ckjnkwG//lbuEFdNYJsAwKFBomuPOYxQrsRHd7NfGkboQoDrkYRfjhYCQeLXkdOE3bICMsX
2vmoerlJq2jv5MRb05pK2Efi8r8CzBtj9DRfyDzh1eo5OvEu+C2OyNLYO13u6jSIlawKy1tbeuuG
KzyD25IIMNiBiwQIh/6Ri2gfsA9uL5+VNrphIHrGaUKUPmMizeMXy3NdQlMi2qmzYDpTxLIWQ2Wn
E/LRguNcBG4LG+S+T02n3b49c2LEY8N/pafunzVwMZj5m0i783KbzrrkMfkRkfQWvc6vjdMb1CwT
b1fdW+v+S3Nw6IPYxQbop0KVg0eu+8EVaSZ1jzFMshn5w0Ui6j0PT3D09hqScsJ980JbYgY/WH8p
5/ut0fxv5NGs8i9CiUX9k/QdjbBbp6UsqtXdaja75f7F2g7g65BZZeWWiymlAIAgTC/WpsbjkskX
+JRFBKyQsZIUOoL6qlSKJkG6D+o4WnDlcl1+8g+80q43K/j8JruIuSmPJCTzSh+ZO+TS5xhLMJJP
qaaG6XQpBZmH5QwpJTtEAC+N/2+rSN3lVG86X83UaG2V2XrqoncxBiWxBNlsx+a7nrq0tTvfbK05
2Axl0J1GtPvD/61VpphsCZPq/8MIykWkHo2Y+QqqfxMDO+QPGR8q2xcxCnZSCDKNuAQNMEmjXgKx
m/c7bMIKm66mXq7t0aWanpr4qCQjXXQeLZ7gZKHLkL/Db5xrhYQurnMkq+vvWNb20BuwfnLaDfw8
lU7pzWOfBUOufDACxot/wNpJLjZ9AyuA6YES1Sjp5DPG36xfWWGCpbkTSTd2KFkbNd9tR+NNW5oz
KU8Iac1gUSjQhW6nNe7MUbzbFTFUjL9jIiCdO+eCRuDwlB+ndV7RMc+kQ5u+Nw1TL0q9JT1AaBeR
eaEskXtWrp1oFqnYsYv0oVrPg2VtgoKMoxkQXxyKH9F5YipjLRY/8y/2lmT56KtQlgmNu2CTg5+8
j1+YD7QIe/FBF96tYp8SD+GmQcNufDbO++TUIQuOSc/dE9+2TAPCy0DlecM5u9kvP7bMMk3cVbXm
ikoDdESiWU1aTQX6NHeMtnLtmIjLqVswqc/Xy2T/Q6vmqXqMGaFeHCPsI1nML7PmGqoey1DhI1gb
uXJ1BHY0k3bLTEGiKflZoG0ba+ks3C8CSNbzWs5arVSDasmTsjz277KCl1of6CW8U7rC8Xnu9Z/d
5Ui2YC+BjW5wpe8Sqlk3vI6x3z5cE46nx9MMMgP0zEJbD9FcEBeNyC9OEjD2GDFQPKASC4m/DROO
+9twz3fta7JhI1YZRmj555H0IdwizId/O/NAUWZEJRh/RQWosmqdXDEyRMS5oAHcNPv0laEoYAXF
syPUf9BDbCIg9T7t7jHU4AK7idfZ2O0gKsIOrH4ii9pmBnO8cnPlV1RlPSzC0zEuAy3t+8r6vp84
o6IIFqjvpLGX65Xrv2AbUROxjl0lKVIWFdwrNTM9O8h6tvgD3htL4521p1q51tFlHXBfSLeQGOpC
ZVg42EdWHyzreCDw85EQgQjMslLBx+WuVkfXUZNg/yA20FbLQK8HBGeztc6E9PFuXpxZbiT6oaVg
/mF9A8qItNT23z/WIoTpsF8XbDiDqeFHCRzkCr3LXcsBI/Dgzhu3H+g6Jz5HPPsvRZaXwWIZ2KoO
/yjsNQFuxe5N+nxXSp/15lBWQWYKnbUNTJbg+PMYwQlIVxiDPXKqavwvn+L9PkwnU2tPLN0dqZLb
FYYH3VEqegU3oTIWqpGD1WS7wQutyb/n6RmFwfpEi0T5WXrO5uzxiTpw+7IeM9aLH4OOhJncj6Yk
FPTh9BqbufIVpAcibYRLq7cqdTXq04jPMAgAyd4h9JGmQsXLMYSBQXKqNL97ZWHpJNnvgAEejlmu
3M/SuZZblZ9yifQxb3qCmgS06ZNW5onoUOVIcDwqhGRGttVZDgOyHnifZ9K4/KQuE5QFqq70x2U0
jHiLfu9n9o2ACguJuPxIBQMf/Rqi6Qs15yY+KoCgYHkQ0k8FcTGk2I9b9fM6hfQuZs/bl9xTxNfI
2Ep9Zi9KxObzQjcqCpQ/VQ929ivfTj7dcav406ieCvpzNrGuY04FrMLZ5Gdb8GrveNnsuOxEPYuS
9Yng1L3gZwTJGog78UuFBUAcxCdPp5rBQOaytEtnBr3NhKFq1JXM6NuF5qygYxB21bWu6hKGinkW
QdrwF9yeg6eNEIiNdnJWgGv3OwA5NRnep9o4Ezq1DxyVF63TvqBJ6l7qUx6nwdXQ00DknmOZApWe
kLXgPsjrSbkDxdbA4ksPk8CnRhQFssvOHXf0xeEpz9Kx4AWSP5/T6UA/LkxwcxJUgR/LqSxK/iDt
Wb5tIO3ECSwN+oZl4tzxStyfiv/nAEgAMpSDnDDEsLVlanFZq02ehJbFaik67hViv/EYzHreScEE
t9Cx2wS3hvyXEMV4DgLPXP01Jbu2m4WcJGq/0wjvwxWBLsR+xtpVmAm3n6rurxA51qu2D/WXgQap
yBL4V4Y7F6Q7EhL/cVs5kFxkZOz+91y7MlKWXxtVicIVyGy/PrKXGU5gopxjJsXZB4MM4CYkKLSJ
pxAFmYT8Ouxx296Z0kt/5xMSFj7CUWwNz0pkSvIu7AuoECJiZ5pWElntD4YSy4uwnQzQu8e+fQnj
S9VcmbvTqsCCCJWJpNKPRVUHvBmwaNOiVEfq2NC4LdVzrd0iyMN8r1CINb9Qv2vfzzaWSICcn9AQ
41edf7VsCLW0UfiPASOzELsxBB6mCa62SWYbhp+g74zVQ9SkFe1EABtgXbemrxYaaxC17LFQBmUu
FXo6E+GwwwE3FVHQBmF1GLSpwRvwzAk0nnhgfNEvd5scvBWMHOWyfseICQ5bZQFz1YRTGWOIaX6m
1ZYRqBZ5KxcmrLt9mTAv3zby6him84H277zMjfOjm99gjK9dJEm04vu+U2RGyqkTkuEmwLkWsaXk
PujA2n06p9xINtJ5Eho9z5+Ewy5/R8NGmdoRuHU9s38YQ7bTWY835pjymbPrn/a6+7pv54ZdRolY
enhL/AHHK/Pr/Wnsro9BTUD9IV/YiFeu0ojnJF63hnJMSrk+OgIFBXJoU2/8LPNvHyp6vs+sQni4
lGuiTe4/t0zbvpKF2CIX9siAyqlKOBAoXz2eHy5TteRyeTd/0jGxxtTdIOx14PHZ9SLTMF0Y/saN
7hTA32KFZiPKRkCLPEIZTsXeorZ8dJ8O3g4oSvZbpJCYsFc6Ia+rQGE+X0Iq+6TWrIODqim3o8vS
nBkI+RE0G6BSUVzUYnynBq4NHF29WZ3h0LEDJ8oly9FtqHkC5W0SxXy7DEQr0G1K7XS1xYaWwis0
1Z8k8i3lNX7OCWa6LyCH22dl67K7DQElei/L1Q9uauto68dvmvKzFRobduycqPUCaNrvuKA0+P9i
huaNgnvw0+rMRvubhKD+0a8paRh+SP+817h0mEs38jijeIonOE+vkSxnj8WQU3gB+6kMzI++cFJA
egFdPGP6xoGaRNmuM9vosQ7FMRUcauh98jDQh9vAjS7dkroZchRYRrWkqZ9wVppNTditmERiwgS8
ivJRW7+hqPQ5NqcqvKHulgQn2SzPYnbaC46YIpncg0QzldZ3ELGNfFpUyLJWn4ja0Fk9/zkqTlQU
HiUf+KJJnPjT1HXabMVlNR6nF3SN/NoJvfkxfaOqInC49MFO/A525B/7JEcHRvI9MjBe7B2CF9RZ
KE0u8/MaPkbeOfqpIbjRey3ZFQp2PV4bhE7IsApZGbWEjcohUOf2A4rSGGrqxjw3X8YaJAHi3FwD
C1Az1AU2Vst7zt31ZCm+G08AtVjTV6Lah77o5szbmaeM3NdQAn+J1MQPrxdwyEqumatros+igORA
0d4sH3trF+nPvr+RPpma6JTeoKr5xxBDJ3cYjgfeapFizT1RzqSuGWk+NWHk096LIr7tjt9ijIuL
AbhYTetdZI/dKcPtZCABVavvRubyeYZDAdOI/bfQpX2rh8Ju/MDVRvkLMOVbSoU0tVG0BGAbkifN
FAdovma95ZqkyELELycXeJObc58gV0Y1KuH9IsNsYnklwf6aivPO2Wit6UOgAViBVWdUBHBV9cpY
uqMFrf0CWtQWs8BYzuLgdQOX/cjxPzHVtjNLhZ4iodnbh0LWcpr0so7+8vCeL8dDugaY59KLiUH8
uLFRt0l73sHyebceu4/SHSKhiAVDiF95SD86iMSiSSLbPkCpHZ5eUjBuwMFmtQCsjBR9POlCLUWW
yiT7azdLJANbZtIZKVJce7GtniXeIS1GLJfXOwxPIAAg8MTSZMIEefZadYQUF2kfNLg/iaU6IqVb
jBuMSqJVr40Wff3IaAJrIIijqo1kqOCJ38U/IcKKXBOdcA41QDbdWAXqjil6TYx1fb1dGzF54egJ
y1rTBeHVXixX4oTENzxLsVASBLdDHNiZ7SEZqKsLvfP30ywjsoPzIPYqV06hi73ZIIhl1SfZcW1D
n22LUi6VQgwgQUxhlk485tDrK8KeAlGNVBSVPWi6kxPedDtbpsadk4LFwZg0LpTBDKUVT4iZFuC7
GZDNbEwn5Ki5eziG/2ajnm08dECmIcfAzBkQ9tlqSh36ELXKHdxBL5shxeCNKw/CxmXnJ7mQtE6D
BvMsoRhYKROSfw6DvZNjCAqiehpV1JYCdtQeOH1ZU8bczZTEiGoCHyASIeN9S5QKbeVasf2BA3BH
TKvaCzRl+dkglamoXG49J/ij4XpYZbdksbGonwYgXG4c2TrF66Yb81K7RXItKUdrKRLIQXoFl9y6
STk4cAzwS10Xd7ODVf9870Y8uZZ0p+WxgkZKe4waSOtzRNaedhw3Vf9gUB1RLcy1HHD1/SuS6BX2
ji1HwhuHh7cWpUNiqNqLr0zypvlQvlyiETKkA9rh0fzjyvz0A8SWlGl2EQWUAaYV0fMLHmTkjDdz
DWsJqwAYvB2qVSB63pKApMScqVHQdaOCSug9O5Wvrkr27w0Um8G/hQ9ollR1n9Ykmfp+MRQItt8E
sBZU8PFv6jpOKvkdHKEQh8bo9EaJBFeJoTLV8NI6jq4VMEjrixdvITydE8+SSLMjwG/q923fmyXb
CQtkXSKRQ6B1/XF7QcVybmXP1M/mHQqn5NYWX4iMcCXHZU1MvHtZ2B7ZPuUmvyVPXAfqmtfh9Ndf
wRXD7diEOjLc5sO4cHL+NXyNF/S/PRIilXOtbGZ89TWa1Ffvck5znfnt1apclsM6ne0JDDSQKGlR
hKdCJU7MNI4McZ7enMhV1rn1l2+JxooUshzqZg+x3+TnXcfrnhseZO3zSEqDOfUDGANTxpQKsL1W
I208u/43mLTrfm6asQ/yb3fgYHiF0E8HGeSdLathstk7RiBgMUrQ8TNn+NZEbBrH34FmUMLuMQJj
9qLpWvCI85MJcKJBKwbXKJv+4AZgJ2rrMD6v0gi8R/+5/oyWnnE+bgNgLMWhRLZ0EHmW4+ByP6/L
EoLCbcI1JN3XuvBdFdJ/vZFakhidw1U5PHIijB5ynhyavvnyUAa6cvURZ1+Nor9fyHYxaMHTHRuE
DsuyVyqZsEw1mw6ir6anf6TAiP8T+/WSP0mnkGjjtDZIQoPPX6JNTVzYjTc9MdM3E65KXuq9iv3G
WS2IEdvxkqUEFHPKH0xkIV12OZdJYSmzPnLJ/+gEJogCueSC5Do/M1IQEHK9IzTzhR+csiBiNFFM
oyeNsITrnN8X68iOkU406nBpaD+K4f6uGWJpV50oPVCZdt0RMf7/G32qd1EmP0j8mS604aOmW1Gq
fkUnmEEiL2tLRYmbvpkACKlH8oqncvtzgw7k90J4lx6uSxOyTF52anPst+GHOTedNR2WpOMo0r08
9JZ/laSB28+YI+YaE5dTCHWA92EPwyQmH2vHJv5/oMMoOpaTs1T6H9JKtA9Ubnynct2Vu41qSmAY
t3L/95stj3V9YvJM1dTBfokEGKRt1BF4VF8i9HFrngf6UBC+z2KmAzvTePL7RJjYyg401c8h/esB
p+s3RakXt+xn82CrxToX9nZPA/dzy5DUnNQ+gLnbcJnOtYArK6IPj6QEYplvxeboFy3Uks57Fsxm
TSRQq8QWkuprVpnkHJEXSjrloPwhx04tmUSc8U+4AUQp2G1fVIWov6CuBSF3RnHM4K7nttBoW7GG
25TFG8JR7FPZMY0Ep2RIVNK4qLA7tov7zgFge1oAFfH6i4/TGjs3zs0cG4yIS6MUkn9P8Hv+lknD
aEBi4xS4wt56V5Zr1+Jh1Uu4xFo0oNk5s6qtaYgPSPRpf8ykH3H0WnatAzOpKuXo7jSqDmjbE5S3
r5izWLIIlnrVFsnxR4axkgq0/cbfdBAGTskHOUg//dqqy/ye363zTXADDkVB9R2/+rS8Q90MUo38
FDS/otEHGXBq5aaDdFqEixiWMYWQyS/wqiastgrhy30ZhJsGw9JA86b6DRTA/KFf4QChPnIH7jW1
nNGwydj8xd+cuStvAyA4TWD0ZXYvOmYTuAU1/pqEi6qSIfR7BTUkX2Zqt2mG535NveyIGDKK+VDD
Yrqv/7HYxjM3rtHHi6nHS5A8R4+MSvKQ2/XWTM+U6hEDmuLQI0L3oUv2s6uBGqOlJjU3tEY8y3Vn
bMSqgSY/9BZxveJ3NMuWUBophF6jRKkRpAQeSEnOmSHo9W73bN+tdvGLvOn0WkOUqswebhS+V1SI
wb077THPsdAHh39IJWYL+aRpkriiizRxSzRaFvzx3o1ggQaTWwiF/Va7VOhrbG05Pdx8zc7DfsjR
vip33Bm6SO9T5lXsTZrGtbIKlEcAsDuO/6mRJ1+kXkw/kYN5YlrncUkuuwCmhopQqInFcakFh+Dv
Mv5lFGyw1Ii6xV+aNd3VptCJ/6hgzRssCNapEJsU54HKGJUxOheIsQKZ9X/Awu9Jt4cT9VojJa0a
LzSZcvnk6wYcR1OsE/vreNN62cbDZExR0IiUY2jLH2nn0wNbVivRHN1/5tMFH27/lggKrW34iULS
slpEaEJJH37UtK8/KxYARlX/r0RZcxiwLy40RyQkdrQgt5raH+swRiwCJKEsrLsLaPCq+APaDh2l
cgrQ0ieGgjLTPFc2Ygo7WDLb05EY4I0q8D2XuuEvVdCtYj778diq0byN6wR++Ffjw0hu6Vy/ssB4
UN+mOV5avHkjeey2d7Kisx+khJInYdfYjPuDoDto6FATGaAYD+e0ZKD0kRErlTstO+ZOiOwvGdgO
etkT937zYCN8FJQE1n8OJmIF+R2ohH6+nUnhAd76FNQ1XMjy6zBBcvAUaESa6tZ+xZZjPSFfJIgF
nCYBk482aVm51e88lXAYDnvizpQtznetDW52iLJFdXKo+bFxjlIjqFF4YWZeWBNhsdOC6SVrJHB7
EqU+UOB3fgwiMgh7j9IXbcvNsDXTCbMEsqEMw7AhdAq+L/IodetCpK3ANnZhP73pO/uQzubwvDD6
lHo6LebuF4oCb9MF+iWK9UJjp6CKRBg+sxlufyCH2kgWvYPOLlw2JxR9w7gDDITF94Uj/eIu/1yh
hRwmo/ByllHGleNJerH/WagAg4zTY/kqP+bpjojdjOT5pQVkDukLt7gZfk6w16Tdm90jtimjEyxD
SoM7SnQeQuKccLXJFrbq3FQgzEDYItGt8ZY31zLXGcK/sNISO4GGNVQ+uivUM2MgMoWekAThVgAb
V8J3G26zYHJQjE9mqhjuvFyhERg96QPMVxvJFAsd13EzpwCPjLLDmQBDvfgpbqJTlUaJkpbhgkKd
a9oAFo9TpP2UNbSOYa8YogdHA19NgVe4xk05sYvbPyHGsTmyx+840tTqF+44qlhf3Hg1l+iZ8Dz1
c2eXlt1NW5p/T0o3bI2hOjQJbZhqOaYab4GwKwtncbGy2roxuTwiFai8vjAdezP0+cgIy/Vlw6pR
/vtyKovcoe3sS14eHfPqdDID5qa/MqzlhjI9ncfjrVAsoQ76j5g8TUiiIOlGeReR8LfDRec+Wywh
8AbohoJiQXaSxtTyp82DEQ0HFPngcCDhFmNpDIaFrRQAiWenB2qsoo46F6lRrkNlVzsHnyYNxiTI
tYeA0YfS6l9z0gYm/Jh6VS89hJeA36QVA05tPf+pXwbGkQRBt1RJSSSbUEC7ECEUUcRCqyB+oUo3
CXC4KF1w0SQzkGcGaxmEn/s4eXWEC4/b4JfW7xo8U6xUi17k/vyVw4HDjxyVJDWcACKEnoIhcXXh
yRf8RjMCXjoLlYceFirrTtaQ4FeqPGEMmO8rxhh+dGyLNtynY0HD39YjhiMKqQnXt74Dajvq5oUg
8roQ9XxZB46j+5OY7DmWoeS5/zC0EuQqpb29WT6eRdka60rMpfH6tREcLswo+yjIVhnbTFATYQUs
N2YvraqnpcVAGYSGIoDKg/My1ANfaKFa/XSFsa//0hisXcoBuKrAj1woQQiEr7dA/VcxVZkmN0Gm
3SCnFiNkSq4K3Yr9GdfRtolukx1sNy/u40COKxrz8S5QiBJdVWSzlZhL+9bjVhd6GcteYxsqMpjZ
Q7cZX6qRlG8/HVWoV6Ix2J1qx3q1RbAxpEtQexhnRbPltHR3dgxWcdLRtKXuoGslzQieiimZXexR
Wb6HwUdFsDkMgHoHPAQzjS260h8l/hfGEtES3C9wfkMBA9UWR+Szw/WTnGWRYoD8XrxODUcMmwAE
JbmSFjUSUR2zcmJiba0d2ExYLXPOVeZG8899i6gizEGhiWUftB9q0ozFCgRRQQ+FrE+mOkDMXZWk
K5UzLgSU1bUzhem4EJzrM9sFe4kWIX0CBpTn5rClFb+udC1okpT5WzX7nYbm2ybOKbLDlSoT+IB0
zrEq+1JlNLXvJhE3y2Ffn2VQilfCtMyZMbu8lq80lo78y061R1A8s2p8kfeGO+YRM/MGGA4nLL/7
4KRwdB7um9TG5Tsu6cmJCJwI1IctWNH3uVCat0Rj1+IDa3nhL/Jyks/Em4t5pbx9HGUsQu+HhcpC
6wmu7IdLwnbqZEQO+uKaN2+/FWEQoLIhqeVO5z2Xp50xELxHJeMmNkdue6X8ldyq99wAQa22wt5l
e44YGBnISPd4Rct4TPuu8eHrjPweUNti28CLgpqfj0YyghOJBs//2T+gvss5C7iaIns8bpo2OSRg
jWRHg910bQ9/WZmPDcBODDKpkhwZS2NQuw3PVEI+Fsm+IuKZjT2G+W5yDgc3A2tpfUesENfr7qvz
F4E+eWmfGS50zrBPNDVKInosbWr9ntB201gqZ07BCBrVLbTm5PMi7q9f3kaaWWd13zkxzi77QAjP
nTHSDuXbr/oigx4rgM/CFolZDd8RfQaGib5bgnpHJJgPxTac2Hi1/Sxp1tdwT05UjHZEnuahZUP1
2btUXP8Mobh+50WYmBfP+w0c9cHnPa0RAEupTnh0m1N53p8bTH0D2lsE6P2HGLl3Qm85dr/9kbx9
W7prFHvKLaJlhgGjML9B6N3i0dZstgLaH8wGmU1F5dAoXV1uQa7kyYAvnbulcL4dwN9vdRD0L2Ai
5g0559oUQ6ELBFpAnIDPeQ8LWTSOqSSqdz78Cgb25RBNaYZqCGH6HaFV4jFFCkdn3Dbue2fJJWrH
7+EDbY2sXazOLedpPIy8v/CcY8rCz1AtG4tnGt6a17FWnhjYcDjmf9SrGMtVGgeGvEdFLSNi7YT3
bbShDyAb4bX4eHP2sKUq0fKiJB1PjrJJpOlOh19Bcar0Q8+zpFheDRtq0zeStRF6HT2IVqXM7jug
i1FcpOxvQ2jtDhV15goKtDimhdWyf4uq5Wi8upfZCM8nzCWtzZF4S0/NJrBqCZRmOoDFkMBDiLb+
XNor96af8G4W0cn+RDmNsWThGToCWzeO4i/t80xGQpBl0vrXd1fFbFkJFRh+TvChI7kj+9UOluUU
OwUl6MfyC+zjTCobmdtukGrOtAnfgiP/rjYmVgUc2SxkBaFcKZ7CqlVf/XOBKNRp+IZlanUWjCTq
EvYqCGCBHY3Xx1QzwGcwROtSQr2gQW/vJzGAyju4sJ4p3KlIW3ArWvB8Qw5oux6FdH5suk5Td2rG
z+b1SS08zfL+/BQgaxsjXJSlk98TazphSCDUnLCO/9doRiUMJ6mRF7Qx3b7BjmRanAy7I0B+wq9J
q041bY4Zd+pGtCJuOEXV7FU+821BcNkA7xXBWy8IgAs4ikiMfYOUSL9k6H0erW2FzIdUGVAlN1HH
8N8Chttu61xcCoitQCFN4Aj+4MMC5/2SkfD+rCT6/DAPxQk9arJSjSIs4X8sLq07xdxL6tfxpZf0
PghYJOCxQRYbrNoOdyLGL0cXggW3k0EA6pHk0wdxRTLh5TT9jSh8h9P+fDpYuytdLqK4BKTno3Mv
/cK3BwpjDdHsXvUKmUhVXqLiPj/QiHr4e81SFUrYTosdRfu+ulhZe5iauDiDgrzXZHxzvNeUpKFL
cAL9drzEYvzE8KTZU57jD+iOGlCTHrTvk5PedQasdcToE/ibF95sVGIEcbobECwA1UtQgWIfZcKM
4Z1iyYsGEEUxXjHNpOWdPmxHxsxSX7k5fVOSUoxMP9Ke+P2thRr37b4OhW+nWDQqRUCk7+0cAqA+
wR2QEjYMXXo4yo9Ea4eSYfnsc2nfQAn/woKeTpa+391B+x8XsFAgaeoDzle4kjmPK/MzM9SqOhSe
MW0YmwiK6JO5TnUiRl+mEgZGAbXK6GCznr+A7wwjoze15jNIDAt3Su9UDazweUonuEIGHY3KDX0n
baezW6U4it2nV80Cm5/+Dgmkn/wXVERtDxfOPXlcieFA5RmZ6hhYL833ZxUZ9cZ+IcQeNhDvBpbz
n2JlPKKXynXlrk3LguIPE7LS5Q3JpbHc1HUMXrRHwcF+GRJymdHXQ2u31BRtMGL47OYJOZZgPsk5
VRNf9aGrIyzWQYvDlhIaXTdmXstui3vRWWGr8XnWTeFOmrUYb2RBpDr1hmzB3FXsoRAc9zEKJn1K
l7X2+w5PPRoLcGnb6UWerGjQ2NEMOR7VylRtkwDvjPos2p3HUOClPITnG2ZHhpNem7BrOP63Cuju
es4nd5Ysjh5iHYeGKcPm+9Bjt9W4DrVtOFk9ofGGIRlK8zQ5SY6ToO2JtwqVaUU3avqKjMUBd4eW
dJxg6ivuxWyT+t1GxEISmONxp0dZbefwihKEsriwaL9xo8fTD7iP9IcLhQ0+6pfqJavPOGDbPzX1
oIjk5Ucyo/fmX/sB9r4Uja3r4/O88VWCsTRxmsGyjpboQZx5qlyoFXHG49l2hamvdILJIXgaFoxx
I/PfV5Ps+t3vWr5MITMNBHBoD5XU6hcRe2rkT8aOdFC9YSeqh5y59qjm4Mxses1NmNZBb6Mj72It
zTKRLgHiADI29ulfi4DtFGEvnylDb9yoZ4JGxMhFuIzhxYUcrc929+0ZAA9KSJg8j9r0P2PSFuFt
oyBv3gwR9a8lfdQxWwKzK+Z+ffTmzfDVnK1DLSlODT8Lu2w5Wkxz33k8PCQlTNBQrFuz6z5Azcoc
1DSCZ4o1keuokIcE/IrNce8Jb6Ha7GHqSce7iNcSRAEWkT2shnaf4AEOuPj2zZJ/UABQoFM1GESl
LiJBEGuRS8ZK61tD8Dwmzcl/nohLYxXdQzA+Jfr4pCEi8BEKcJjkGu0bnLodt7zz9rHmpsW6WAW8
mTraqRtm6BcUROK0QJ/yCHS32CEvaVds9FkBGIa48/A3qe/DEQnWOuhRqe/cFqpTeuRFM5/3JUHc
XZeif8RumRr7id/glRtJvYJ8gAfsTq69uJoKNAkpskGCn6n1VX9+RJWoioDdCedS5CVNNuOSpA2v
wTJ1zuEsDXphn+cot4xrmhtrf0b+CvA+5zj+Nv7myaFKAIc096vNWtj6w1DhpT9HKZaWUry/i1ZC
HvaAANzL1CZy/ZKmGjEbD+Qpxhi5Ieh7JNIpMX7VFr3yOH7/Iq3KnK56efrFBWzYewTWEoAqpNxk
CmSCcJ7wtE5bDsFElSe1RlxwXMQt5Tr0p2kIJwoUVR/T3VBmBv69oAVwL2X5Q70ogv4Tc2Jrd8xB
fyO2xuhwFZJ4bzaVO+Ezq8rR+NdPjfhe6EnI362wL+775JTMwhrzB2QX0d8pvM5cQf4AUJU4/yE+
GvYkt+S305y2X4+qJrhA51FPxKwB38GNmwzNBw0Dt9ivggjBUc2hr8WoCdNFaGyNPML+OWLxTOVa
4rm5nMIPLi2quxrUXOz9QYgMoIzOLX10FMOY03nMYVStNLgPxWb6+At0hqNCgRf450Tgzpkw7lF9
B2e66m5NH+XqUFU2MGcJ8IxHG+k+whleOtGDMT2XFDY+2+bXA9Qj5ZacTIjqKN6yQWkgh7CQKhsh
msUf8qjBoE8jSQDx+x3VUfb/4Ix9EsSMv2s3UKlhRFGmE/H7OMseMXc+dvY9lV68ZaoySNHTpTsw
ANh/palAhSit/Fo4se0BoWuBndWmy0CV2UO254rQJYjTUh1FCcixX1GzjKDpUCIeu01nJ0YZo8IZ
c9k9Io5CLe9hTjRrK7+73JiTH3YFkpSZfotOsnOzHyacaFCKxyXvoueoc5ZVV/Kim1d0W05IjdwX
AIhGb3qhbAakAvij/23mGUE/YxFYVjABFUp/Scz/A1DKMfobq0jfpaOwO01GtN5TK0G79XSRO+w4
787YTI5BLsIjNNOM3c2zyo7rp4Eu0AbiBN3PTZS4kYSXmQ7riq81Q4NqezDQD18gSeW+9CRS8fi7
zpBNZ6cRfdRBt8QVX5SvGKj4CekqZUFjSfh0oOzH/qHxJiKIB9jxMF21DdzTYBpOoSV92JAUqowl
gKpdBqnBOuKW5Ol0OyfxzVL2bNVVFrsqynR8Vxr0QfTlqLhKucs20VdVXXPmKnuVlOgkap1kbCNL
DVS+h0GsryMXxSL/vpf1FbAnvpPMrqHLbPCj7FCtcW7MrcqHS6b7dMxt2OYtNx2PJumjsGpsvebR
9k0thITMa1G+uy6IIAKMlSVUbtloHsArnT7Dnnt7EP28v9HD/T3XuLlWfunl4A8zhAPYgZmlr7mA
X+RbMuHyj1hTgJweVi8qCAikgRp8xanw2ziK4onbZ6DQJuNcos0BUe7Iz7pnm2Xs9D7nCiXqYwES
QZN63bnqYhXEj3lRnXMo3mX8ZeZUHfNfRpw95l4D39efTYigalmd32LXfUqLa5jTePJJiL/Fb7o8
VUzqJ6C4D7alpdAvWK+u3nuBkOEBA9tqPs/a4wkpaSVvFd5+3WljIvxQ7IGKxr5zokpe3GmkyayO
FxUWRAHMM0LadDa3XXgXewfurv+0H3A7i728rINQoLVwIqlHPFgUTqB/hUZdjtlWIt8azKqiRWvB
9krkDxqxrAWUAlomL+15DZHvOiszFlWl/59UEhg4j+b1MPCS/rczvRRaccXsW+m7gl27ar5jKcfR
37rcViZmIQK0kvc/QLaZFnswtRlm6++Lese5aw8gNQBBI+hIJ/MVRX2U+KkrL1kBxBEguEgz9t0j
WUvhx6HMCxBUPnQyiT4gvvcxqJWHoaqbtijZfGvdU/slT6LjFe7I7SZSPtZoEi0kgYJDm7ta9Pph
CfDv1kShsOnbgDXS4trNo8lvufxbnAouQWyNndOLNzpadeoh71lCQe34UN824M3L7Q3l0/hd+ogB
9FgWWNXG0yqVCstQ9haetQ76z1sSjM0SUfiPs3bnRQoXU5tuaHLjNue9NurmyfAATAQJNM49fkgs
P/uyR6jm1Z+ZbIBU7jyNnDrPeoU9HmRuXLY4PpQdY4P1W7LT02w9oVl9ERSGPN+Bw1zV3Xnu9JFC
d1i8flms9AXkTsnwTaMjLRptX34aUDabOpwKcy854g1ToYTARro8qagkEQ1ldbc5VVaV6qg9nhGT
F4vCxpMGfZZLNM+Q3zldfK+Ec0jBgPR4appWZL4b1XQjt8f2cwa56lvucYHI+lexk7RLNCjo3qOb
t4BsWkY5HwzsqstnljWjGNpOAruKkhlIZIbBRMRWk1jKqjI3yD5OJUXPi0f7AjTQKscGnoT1Oefz
p1RfyM2qvsgWcgOg/ZbXQI0xMYCfK7c0ediLrb6wvlo6PhEcog/UVBC690JQZWBcOJtBlh9o1BXm
9Xswvnj2Pps50ZUeoQUAKzdudxri/TKhyVceDEjZMMgD9KKCt/gmH7pV8Gl4mGG8x9OeqUWVDm0w
IQeX9h0GQa+57hSa14azw2mWqqBgVD18TAACjP6Az06S8aserK4Cb/rrjDFoqY4IGEBouNdDkNnh
V29kVQ0qix8fFuzJayC0bUNQqALzNWQ3CdY/R+Ur0nUXRrh6QM7MeljvQU8lRndcVTVVuTiUcZRl
xQc577Hh1UyO6RyQz6ZKuCEv++tB7aLxTl4WkuVSQ/4Va0h83pxK+YmivRRYJRvQOMRSViIHrHNn
zJuW1reMKX6yVaPbmVVdjG9X0jCZOIh5v13tFCOpoYoybB56nDvJHnrgA8LU1fcYOfaDO3ETGjwt
ZZSN9fw6Rid/ZM8+ptUQFPDGfCyPVCG1/nPVIuTjhSbxbYT3E2+mb2DEth6o+Hf3iI+JEgaxuiaj
4mBHln9PdDh+D6XwQFTAT01Zfp8xpC5hybbkrpcxZbggy4f6wvarG0TT2kY0LMOlwd/Y1MfiT1Fn
Ygpfc7vHhVi/+I7pI9rgndPrposAMY3Lf/B+cpGeX8B1mV+F+4mHoykzUkG7tiy7l3AKzhcbBW94
5fP4XvQVKmmKNRXUQEuqB9tw1OncIQfYZHgdSyGWP13H78UyJxq8PFVnROsnNEcu8ojQoFAq+KO/
fEqDr2n+VjL7KzpPmqfOpAAXIgBXSpChhOBUZLDJ+8JWFESU7tgZ8QEzbIwIBKt2RYGNCz4cni9o
UiFrBvlQeYAg10FgMtKnRu2fyeP1a8xJFSry9ltlrYRBqsqzWqz+7qLbxJyb7lJYenYdI1fq5LAB
PX1LtkBmTUhuowcfICM1BNPDU6fZmnISduLT46IOIU2u8Bx947FPi5Bkpq7v0Sqn9leBaXtjKIK5
boWzBEs9z1sazMf2qoHveLEAm7OoCRlM3UarvX/aGqx85IrtmQunIlWfoOYMcglcn3Xikn+ZDksh
q8YnDc+0R93Bcsr9bvG/Ayg59+LNXVnWNmDenuq2ztNjQDn0Qi003rvoW0l+nZe09/XWSu4U53sA
8h2s9tPVKc2B4399Z5irf6vZaVNhmn3UNOar8VolcKN6rKoORXD/AZtGdtlq6DwYeUkPKAX5/rcC
k9sTiDc6QwJwn24JDAB7VUHMzybUM/lz36Alwdzm0Pyj008jH9or+sHfRTPQ3h3S1GH51AwPmSsc
F7lxJjDFnqwbDDXTxLwSoOoxRzAmEI9NDcxtfjbB4rGs832pf4/W6HXZeBDoB+rJj7c697qBsHH3
Yh+TjEuwXXMl5br+FWwzit3JtCbs1ewkg/k4aiHKXlCy2p/vbuOSFM+FCi8mwdabKddSiu7i8pY9
msmUjCFnDU8zCVscicvFE4je+PJgLlEY6veVRVTvHYxRPQhU2rghiUUN7B5WNvRu3tLiCPpebZEC
eCNmuMzRejOP0SDCE7Cdeu46epTX5LWuSCN1nExQ1ISkNkUyyCZFhKQXAejEVHXafEhREz7o0KMG
//tLZGS4iR+y5JHl/wf6IG1phwAuHE1v/HfZVySYwkVCPiMv1nrL4s/AcTlvxT/U930xB27UMrfc
4OxA4HQ7WZkF4neTRaXo7gaOAjUBszFSpHW04tBIrebdXwl3Fx7CPjIsgr6gvyK14Q79KCnXmqO3
F1Y1yRr5ep7BLIwTjX8+NZhFdeJK2ONzkLGBRlaAETOgb8pdVxlbeZou0rHOZJTsHLv/2rEBCetk
go1ZJoOl8AT5hxnz+mptOLXJz2nQc5gTghCKRocpQeT8R7R3KvAUfgaWD1wOOjw+rGv9l2xXDGlG
PNVSk++obyktwdYcZN5JuED9RSpUe2IUK+8oGNMy6c7RFx7WrUwiTuZPuJSJ+/0+LF02DkHafV/W
I0KGq8CibZdsUZvbPkqI97vJoYjOr5P4tNZFOaZhS1mK/d2zn6hGrkOvrXwcPVYJGMM11/LB8zMb
slDyZGki13Ig2Tnxf9ZvG7rjy+SKP5xqI+7TCGvBOl81wCm2lDZ9a+2QYyVvMxv+h4qpCg7klOT6
M+sHhD/rZ58va2lIzhxuyUVjofldZShp+uGQd616Wqt38SFMjcPtZnIe7gO7OKfRNFXX47DH4o+U
vjw5vmFi/LPJtYsr52cOfXQZQNwsyY62GFV1MGgR4U2Pi+Dh5LXLn2iFBy2KTb53OY2wwyNOlO47
yYGhvqTnjVPpEUBGfj01RTDmJ0wS5o+7jIEXO0Hf4m8ZuHx9neuc5q/laEqLLmqBibnjbYvsB613
WQ0v4lbaKAwoxBSfA1X5Ef6o/WlR6ecUrJTCpUs69TDE3joefhKzLu1Y2GX4yakhnpD3Z4np9g8r
ww/kcPHTz1Aur5LTyfepNF9SkHJktepm3iyuZjLn/x5EQJcJkYLssolhk8uoMrrK4Tb7j9F4aePm
H5VsbAowq82BzUuE0GvdFgert1/4Y+scGOzQm3fY3Kfe+JI8F/YLuzhWGlFrYa5MVnlRa7chINLf
zU7hhI+AO7hD7eWHJzN+cpnDZqSuf8JOB5DqcXRDqo+wJLXaQlDbBYdmlnRZo4iavO9FQi/GZAaT
WkhKnI7nlI8yoJ1xLevECYKk59AOPuiWqX5YpMHykRnRT66KGkbxk77q4OTwGvc5IFlZSoq9I4WK
BvWwVxISuHednLq32/gA5gmbXWxuDHldh5AJVWts0FHK25LYUGyrpbE8Cm0CNc4QhIUn8M4X+RFM
Huh2A2i3iSs5b8p9TPErJKiW936COA6Ieovz17wf2q2lq5owxd5sVLwyBbOxs8hsZ/okj/8b631J
BxQI63vBRTcUgH8hyvGSN4qkB/BcNm66bXj9/JWUWZDtDb2bLr4dNlXuiPVVREqrZVBqHBmmNabc
eZFj5UX+S8Nszc7c5pVa7Q83jy1BpFXxOTKK+89u6kV70G1Hbbm/FjGi014xdkXuOIh1EZYjVkRn
/LYjstBl8Lurlqv38mv7FbdrHfhF0RP/A+SXifKFKdNRxteLVyBYpvM/WMZuvh/TEws1yvQjnljq
W+9oJt7/lXmzvt/GqKyOwwRGi2yTkXMDXqDDlzRvhoD1s3ugXfYt5TE9DKKvvb8YtQRaoXr2jw/v
R+SbhRVjkRQEOcCWpnDMqYxC6s/z2JdS+GeTDPDJG8J3sthjOx0wd/6GZw4jmQNucnyprZfjCFMC
dab6dFFZsujOT2xfDpJmRvmbQ/fGWuY0ycjXQl027isY4k+Z6CFFWSbhmlymlkiLRgMlwha0AF84
qd5DfDJ3yR3b8Sa82C+7GbJwfZy9hO7wtY1PSskX94AyxWAYGJS1Lte9+MoGZ8z0s4kXyTlQxUKX
bLWFTb386nAAeT3CAPGRagErNGOkc7lsIcyl283udu3EFTzV3n/RUFV4e43+cutOdYy4swQqcZuL
Ik0d33cPAXiHa+q+eHxT5pCgZHi/O9rSvxmMK/7ZfHzsc1sp1Z+lUq0k1dDkrRLkrZ/4dTOqiy4w
9GB88S85ZsjTRv3j798XqS6WPy+rkaGVspKH7Kn+s+9jwJGst64S7ah+CUgpiTN+tjIcWo48pmPB
a1gsYC/jcXanQpvTk7+iEpSZvxekvSKUHpkJkzOG/qywcA4UNojY0uoRRZPrWL3+hCX58EKTxVsX
LRLSWBSsY0zEzw03bUAVpnA7OKR26/oHTqmbmtbPVOHFwT7WYSQiBS9rCedfHc70bOWhD4MndBC9
c3T6H7xNRm3E46GC68e3PiObFarfBGofhhtH7Nfg2whqZi0PzF3Ko6uzJM7gBbwcncS0vo5ovOlW
Glgepyq6lGuesfyOWCpI/vB9Tzn3TyWZJhYVqJOWQ1mEuML2DxtyVkZINrrioJYuI549GyyAOicz
ClPqqtX+2abfp+96rpYLiyST/EgHHnbLBzEJlElvFujifiAwEe8kdsgS/HUyo50KsUC1mkbBojCu
urvru8alcvX+FGFJMOW8eDlG57v8MDQEKw8AZHZslAhPDxxk0UXgapEG8gITaCn9hcXvcLpOA3/M
TU9ZSH36QboSMj9Hsb+y6I+oqB9D6xMxxBlZnxPFYbXetU/uEp80rvaSyHlG35jaOkntmYj6JuL/
CBHCgUp4IjiM2fh/wSu6qA+VCQZILh4Ggml1lsBZrwhPIbsw1YCsuMQKv1dPTl/HzLglYL+fHUpk
2oDxPPxkncCVXZiZqYPXW8Sgctuiu4JkANRivXH/afYZzXG06aTmX+ax5EFFc53BXVw7XqN4ClhB
FLlzrFn9d3umoNOEUQgUJDVOfljDOzVcTLgo+jZinz0qbRRgxAbtRnTUjlK48NpNeCM1QoW4EQii
az3KPhxZUwM6NiWktfSdFu2n9FNll/kSgWuQCBPhtVaVQBS5DBh8Fefk/HdOvGtbMzk4SfKZDDkL
fSxkgY+s4mqsZxm+G3rpgPl/ESt4yQ6ruhH5UuNosHgwFi2qEcEe67jbKiTvd9GgjI1T8nBExATG
iH49Oxr/Z1EZhDUQFAAyCJj+gk+zVZdweG8ZL3VMYG6pzJHxvXZiEG7Tz2/IisDh4RUDM3SC+F/7
B6mVsyN3yEg8kxek4RUZ/a51Mgxzhojd21Dk5AWQnYqdzzkjIpeXxIfhbq2Va8KSw5XKRi5tA1P0
H836nK+BIwB0ItJ+67mNmibI2owHf09Aj7qRpY51YGCaM2J3iFd28TIo1SReKCdb+HypCTToFl4Q
E5lQSnYfBB6Z7DYcuRxrgU/pfvbposbr5bcO+kx9LCb7/IICxUrBSAGuSLEQKhufajuW5ZrODl4f
/IAGNaEtmiivsV3u5bPcJEcgEMqv62x9wQhyfqfhOrbt99hjx71HpxZzopnrUvP+gYwdUuhdNq/O
LhynYdXoVCAxsfCp2UNXJZ4hjrY7Ypveo61J7WwMMmVfIghMOG4i77uk4EYl/vuHZeh94f5CpHBf
ZkN9YtsY53AL/tclabRwG18cp/0RG3ixloCiAzPx7+3reDR86RhzhJPSfKbicPm9rBfQj3h84KhR
2N6v/WA/ELEK0U83wkGUADedT3JcaBeWeIHzaDkla19QQXS8QcgFX+xjoouamZ1UM9vUDjOFo3bG
9DIrIEJrGhhZVEctJ9DAHBph012qNYQLqpqR3eo5Nl3pZoAU9eePO57ZQipJeD/kwmH1Kwj55VNa
OvG+4EpkAGULkmf08rpB2cqJXO1d1HOBvgLc0t8iqInLTLjcRjM65q/KoPkh5lujZW4ZXO7LWx/8
MTIsiUJeBWjV2Xsb8ttFA0hNF4VWU27RFLmm/0qhuAnyMGaUq5zzvHHDjlzk/dXcCt3HIFnuEBkF
Uvf4hxOY0Ivk4IVLTwMZGABAEDJujwWt2Ngvs8/Fp82uAsmXwYjXEi3E6e/xW1d/ZUVNhzURtE8i
Hkq3w1cGtJSaxuCbuFUlLckhgFf4htdOsp6pAuKccbocGjTxiXlUchzJJdrvnIw9S0qrMyhaxBra
eYhmTmdkhAYxIoo+q6hdyntdumP8tb8wIMBTMi9MuFjT0ffzgSbSlrgUK+4gm3e+gIzI9JVE2FIy
EukbgexZzFtaIQXRnzOTUn/TQDa57fIViCgzbw3EZLSHk0b56jYmNk3TBRTrUxmmuQFSry95/nJE
Joz4/uwI90NQ2XzRP5xxjEGMmxZxoX59PJ1EnztV/nSZZhAimRVRL0VLENftEYQwNAz14s3DTnOP
OQy7998gmGwwVbjc5u1aT6WQKAPJ0euGLQ30+z1e1cUoqD13HTzi+dqfvD0G/riDIhHXMciOoBpx
vQvATfiRbtHvRntTvUSXIaG3OjsEGmTjeBuSEjh4mTwSe6GPGDG7WYBIDdcQ3vumQrz/DzBGhpc6
bRMzVRBUzDkPHO73mbTeeA3d/B1dPzCFrA69HocO3SLIxZmHX5CUIqR/rzTw7dKckcyK5vWioiEU
m547/SqZLBnTDhoLYxleJKd5CdjqB2NZaIKnpV+91UK1WdzyI+Dbac424JRBvMlptz4kTbhGcWEL
0zOpl543ojo/uZCiAstnz3v70685FPuDg0+qwdkjJLp8RDdskN5fzg9wzew/OWmZBOULFK1rgsNk
hRiK2pjxiQcVUmZ54to/BLPgxqOwB33dy+IWqv4AXWFQO5DwK/y19PkBLrlr+cJsygkJfuuiQql/
k9RSvHSccVEnRtcMjv4qWe9VZbkYkw6tfQvQxd/Fv1kZP0zYDxSdeTswNGF01zWPtA8/zPw8z2qJ
zd1iWdZxgvqE427/WUhVqGBR5Fd0GoS4rDklWojRrye0Z2hmLBQm5VqU5eBqdGN5shy6PE17c7+v
YDTfLE706Ih8BkFcYn2yw8kp51K6IVkW+eFd6XY7Y3Oibt8wgNPJ3Pfb47JLaRBg8N4Q9mjLR305
4IMrWh5sQgAf43YKoo7YNR3Pkq+afvejWjgZGnQTpHmzTFcBjLAmItL+jd6Tl9WBrUDvrYLUUCcU
QEkn/EKl6MCrBwOKTm8Z65VEYHPnj8U4XxSrDh4K2YDEjnQuhXJykqNpUDsFhagWIQ05CvjBYsLT
78eBeyi04icZEYIJXq6bx24+D2hum2nQdQI5ITSwe1pQAbt/Cu8DNvag5myxZyxVcC+7Z/e7l+cU
cLvN8ID8ZjOfHdd4C3eW76o2XNFE6s6pXfyH+kquJxJJCtGbpqW9sETOOeTH1pajMiewunhSoEQu
8NSGAyQOla7MauWf6VKONloprQORD4BpDYPgmawU9gcEHrVzFY8+SAcsGH5BMwsh3oLvP91kB1i5
9KXWyQc2Seex7C4oAH6QftuM7xOtBBTNPr5RWplQINu+Hkcyvd4KtaSWpMQuB4hGwe4lU6cNNY9m
RME8okwONhC98l+J4/dPld2sRuiD60ECBEB3pQc3xmQyiLiGvIE6UDnv/VH/ba9liSWngorSDaHj
FPry0fU3zIRS1DWUGY/PtgqswCIOD2+x7d3YTsAahWMxTj1To6hvbiSHMXT27BcOMdX5hOb4UXru
aPdgVjhvG4qI0A6Nq1WnLNq+xlT16sIZSlpp80hA3tHOiGc0amUdbG7V0t1pRBPO/BQ2+LgsNAEc
t4igEJwQjIk7of7fb3CqVVK0gbNbwlzYqbaQrfzEfJr9t+xHBLEDoNEhze2/OPKnH3U62y744BAt
87haQgDV7e7yL0o4vJut5W9nF1EzbEsJPrCL6BLNZQGR1M/W1bM7sjD/sCRGJWs39H2mCD4o/XmB
2JAUGEYWfqYegN4GO1f0Xm1+jdUT0KBi3x2u6cRN/YpXCO5MMh9L6a7I/8p8brcozxpqhfyrlQAO
pxHoqIc2Iu5/GJB3K0riQzsZtytCIaIoZh2fzrSH9/yKboOuuT/TOwBWgiTVWse0BphE6fdIyuNH
P11JSbqCQknhco0WFogYo+rVnZlMbaHaCPSxeaQ0cjWNAIQa5W0olXC6GPAolLM13mPazXATL3zf
5VYYV5w2XIqjbnk2nAXGABPUU9iwVHxFrQhF1o9FyFZGmRczX+DuZiv7DM1t4gdPBFv+gmEuksh+
mvLDYO0mcbaijzwsmicsO6m1LNTcf4CociC5aZLRn2qNjS9EcySiGA1aNQDHkyUcaL9KtwGOSuRR
ieAEvjoYBevIVkPkWvPheBxjGa/afqbTzuzMQ94hSJZoqyBwfMaw1VkE4Y4lWn0N7yE7TMcLDbcI
q03O0skbndwSdWrwAfxgMxzRyyb6KPCBww6oZzSTo4sD/TEJEre1eb+z6nXr0mvSdVUdAguhSOP5
lDVusB/imaogbjtrnBnlBes+V3foeSpcg+4zIhXqwPdnKOTV6dAk8xebK9pw184cXG0awrScl4mG
LeipNbaSbczGkyVx2tDTHsAz41D+DCmWYhHmQ4ahyFp31WV/tkCEcTxoouSq42nQUwsmH5a4ikdk
FhbkF6yToR7gR8XwTzFZQk7J1h7U/c72aPJZl6h9lZeOjbnlceNJ3cTAGK4WLcaLYpXWsvLJ9QVs
7bMes9t8hcPMOnmXWtCWcPFb6eKLChJCssZXM4dnAcGWGmTsB5eFSeWtuGZYy24dflbreQnzLtSE
wHi9ZzTNK7JkPi5o9nXtH9S+Eqr3J2uWHnsaT/s/Rsy417HD5S9Kwiq7MFlLTpjeCjqfXyiifsei
KFOF/A14E8SCY+peqQmhNmbO+7jqc9ZR9G6eJBgalW3AVKGSq4xQnDQWc17AoitWFEMwNMWC8Y9P
plly//YNDnJ+4fjlGD88LEeZ7yxSshlN0wb7SWjT1VSm0rhd9ZSaeB97qxtVuZ44Qx96yo0gMXYL
9XHBMB84mO3ZWb6kY2i4w1roFEaWHuBuHOVUPZx/gockLIgEvi2rcmHOpzAqADaPVhc1+jHBvcPD
tmJqgIbe1NQopcqAgKH55XwgljJ/OGifAhcOb96aDUs1VKUH9G+wez95FXyLmQZN4vZ6cVigP1+D
TC5mimZ23tqSY01H1IIrqlgXNcJt7q0btD1pndEI82HfmKhm8kor+mj5ZHycbplTkkkV6+ySrjWY
rY78qA3AqOyU6lFhRTABC9CWTTD4FSXM/LJUxzpeIZKRtfqrH1i9Jny+QqapZqc478o4LBG740gP
7hb8U2sRJAwv/77L/pyev5VIwySu+2jtk/VCe+kqixMSdDOjJ93Jh9NS17CGSEumcV4ySC31lK3S
oPKrMuQOl9IKmVgk5HO7xl9oaeLEqBuHBBgNbCs7PgJRCJ3qmsXGU5HvX0Zgvnhd+uFE6CmihhhB
DcYmRTlY1KFUB093hceTSWDU8CUOxvwZ5C1PRGP1HsKwtPRnXSmleoMwqJWxj7ptb6z2buKjWVx8
J2ttdlx5v6P39VevHADuah/3QzXG+1LVfqeC6wky01jUf/fWCucbXcmDx2Ek0QauJc014J0FFRfj
S0/alB5xTvHvzXuangGSLs0xzm4AuBtmH9MNoCOh7UBjDRvE9DVwJa2+4+28jCTnrN5tVAfTeCAO
FUhpyI7uzXQ34YT+2YzJiJ/oo7k2TJ/nNB2TGZ1cBuHclY2/ccBYYPExtR4DrhrDUQjFhiVX1UyD
HDgbw6yunRjdrDDNIUkzCC9DSgpVAqSrz/7Jj3mj/oXLOx/9m+aa7Z0Q9MJ7YxCl8e5blzufuFdF
T/CEAaObrESV2QotUBqdPsNLf4Shde7ZONghS4FDZg4efq0JEHcijPUZjypuHM8mnX8bmPJ5rBCl
W1/k9TG0pwGi8N0czngGhGXQP/gWn2XgVIZEbwry7SnAoStAKhlVQsJ+zZSoV+597yPQ2ZGLR2ly
z25X4QH9UDbx6zEE9PDCjcqjyzKAQGG7C6yGOvWWouQ7VgRPm/2tOiwUbFi3mlMnrabsZ3Q75VJA
9DabpqHzB22WQSeAG0Y56rrVWZe3WVliX8/DLfGcfYg46WMb28E9jmnmGozDBELi4NYhxS138/NO
ft/I9l06+OlUhyl+hEoMUN3lKp2CWoxsgGyV1RspCcY1SZvsj8q2lE+9NE5uwOJMiN/S/P0lpkS0
WGJxgHc9+kpls4uF5uzq9cJhursnNmneFlbbjWdpzMY4ZYpeiYJvISvu/nzeAx6hqmE+4RGpt6sZ
ixQal4rJtPHxyynGvH9GIX4sdBhxb3qHHeS0OVeMWCZ9I6ZwTAt0ARKXlDzPfFpTbmpNIb2OWzJy
qVGaxNQUN5/rniHZWvZd9Yl8K6CmVBQ5AfyQP4BD5Nxq46Mp6jxvpbjD4CNZbqxJh9nBJFG5UedV
GKvs982Qp8Ry6hvQ/bMR9jO7x7WFR2JknqeQgMaq4qrIrgZocpR0nY2bD9vkpmfao64uBEooJs72
HfNC6bcTviwDxi9iw9Dd5IUcyJ1wUd77OoAoque4OP5aAOwUyo/KhuC8BcEnQbAgAsGEPV2CKcrE
vGKAmyX7Ti8Qd89nejiRr24aLOoiOsLp0cIWbDqhRkUKLvff7cR+V0i9LQT+ocFAgkVfadP/x/O4
ADxg9CBNb7F8SdV//zMcp7LomEpZg4sTGNVYeC6Z9f1um38v6I0y2v4NfMrtU4QmRsEYF9jVOk7N
K7EVp6O9nJHFGXUgl3ldvx8QALrrOgNdbZjTvG1SwAAYPkyPXm6/XIw/L5Uu8NmECdj5OC9QaEGK
rY+MwU7ya4b1636sD4cSSn3SQPLVsNe/0HYkOggqm5GsZ/1ojYELe5PQb9ACrHMtpNmbNWjOsoiU
Y9gUTD/i1p0PpibBbe1DD4sJ7z7/5V/RqUkQYTmp9OnPS31dyEmNR7t49yM6wVS/zx2SbP6BRc3F
2Ot0cgF5RpYneuIBv9eZmIgdvjBpImyh1iKJ1TSZeps3MUTWfS76iH/f/SJuhtSJiBFWOcrYOdH4
r/Nvh1VpQHYnmwSAXU/Zqx+OjTnZ8eBmB45meg+9KgP7bZ/g78buFGNZkWZV/IXVlzx/Bf8xxsDG
E+xJwMgi8UTiQJRFO0xaJk+05n6fhaUhmURa/VnwwAb/6hd3Oy4iuoI5p2kjeZ19V36/5gpWfnv2
AUE4NeMIkAZyr/JH1OUcf4ZOIT7yAczfd9I39KaED54fQkRLDfyLTfBtKg83ZsmA3242aCHpntM+
aVVDIrMCZMEVZUIRY/AHCLtUSOfbmVcrzkPP1zXjvfm12/OrIIHXie+7lUWodV5BcEw4sMRE/bV6
/otO1qmrt+OOIW8lWNuGtHI9ui24dHMaJKOQ2LloP0vmoU3ejZqcaxVKBULuJf69wUKEz/XKx1nX
vsSwaNEe9HF0OmcOzGf+FqBlqSIyjQpHVqK0gas1fr57Kewq2UFykUOOPrQdfqvqgG6VH1SqW9eu
iIeq+UxEHy6NkkUahsftL264dv9NMQDrDnRY8AXlsfKobeLxiYc1vWo+GPK9dIluW/wBWXzvn1bU
t9YJObtXQc9/uFo+sEwiefjCVT2spiF59Ni4QxuA7hGFToe+3WciD+EEAhOoN3oivh/wzyKQZst7
XntdPU1QMO5kJbb4o34Sd77jFC/CHWiSPOENhydo6cT7k8lMr7tvs0OKjXmF1VsxywVj7Mk3QCbN
wVgJdJueM4LKuVR2PG/e7LcZry1ckR+mf9v2mbxm/u0eNyP16RTb9t6J66cxeUPzzcHSUcIBb3kw
+dGYIo4yrR6JITnpU+F06lf4j7XW16GQSSlWJIMu4yqigt6QkR19ZoBiWP4gHrB4sfHoav24Z07h
ZIF0y5/aHB8jXUBVdlrJqkQmspYD6zdY6XDcOaXgAMH6XW4yfUwBu6Cfp56E9kkBBqBr1SIGgbzR
0x/tYwOD4Ch61Lq5znMwS0gpEcO/ImeeG5Q9/UnPzOcaa99KtvLCHpXkoB0OkxfCMei4U0kGw7LC
4IZLKCklBACjtT46OXDB3FNN2JgTNDubu/lXDa7KvDYvH/2skfg2Tb5evfkk3RByi3B6jgwJ9/f9
0NvqPMnY26rgOt8cZ949Xbjaf2XgRcIRbXKHQrcRoNEpZPQgnE6KM4uI8IOGmrJPegm/0XtfblGD
Sapve/jnIyiLQ9dRm61CXTf9q4a/TJKhMtBKd9LfMgqxLHK2HxvAbjFRU4hlM0xBZwn5PbjeKMPA
wKTwGiu+jdPxKTcjic+sMLeXcOv8LpZ9nwVDIU1MZyFGYaf6K1+iqHwoxNwm5gv+VKJs2Sg6eTH7
sQJbB0TkU9ynYdT+l/s2wnL31am8QtsddK5Ordv79mdJfL0XqmB9MfL8R0JqXn18nIRxBdFdRle3
cc1Pk2XOLENl0jk8+vR7ktAP+s7MU0rlOpCE+DsdWE1iP0GW9xyWPAetoah4AOkwlnkCm5IeVq99
VQG1zG8nyXE5gyYdLyo0g6yTFeZWvVi1METU9R3O2OIJcMracXWYsjsuPQgAT0YtAbGYqNTX5N7j
IK/LImRJ4IrMK2PbCsTw3lvW7g/xhDCp1Ia4RtOQ+xb+J3zI3ZqclWEH99czgRmAsW3HEXWOn7gC
53BZoDLHPFaZlMPM/ZcK0Lwrm7g5Y8RiCpOZONkivwnLBBiVnklirY+KZkKGMFdETKbrRBpZIoK4
d9d0Po0518JirWJ6U8hil+QynTbUWx/ZauooSQg9A1QVwk2m7cLmuOmh9g3nPe0Jb50DS+WhxyR7
tgyVEYYjYJcyiUWLthrrbugfoGOGqdhmInM+LWvKgozhcZLuJ7O/qEVOExaX65z/ypq/X0VZUxmP
oMDwCLPINEJmvNGZBbG+4DOk8nCoi9f/3fPTwW5qzlyaaMXdwCRGtNthKystldPrXz/nB7AZZ/2R
oLcf2nGe6hinlm1+9X1haSbE7kexsqZzkC7kA0AihKGwpqyoxdNxYWANaF8GXtJvwt4MnpQPzPg/
7se4UsWtAzCnAKvtC/YH+JPJPYXaV79SL+TiZfiQvqAWR8qjvZfLJWsRGb0dHwiyNDK3qvfVCJhE
L6yA3uetqAVGi9GlMdv2gt/mBg7Wju0GsQ5iWiRnZQTKhbiolaSLPhMi8lA//itoqR33JQNjvgFo
QWkt4lTgUTxMl3DqUa3VIo972jx6MpFcLUNQLII+rRvFGu1zFE3xnQrSZQibuqK5l3jYtJIPbHLr
9No+gQ0flpb8PRFhpod3mV8IWfrGwo4Y1uU0DTQVYrOyRB1TotMjMKWbudSP5BqJerb8BN+ECfoi
edbWHHOH/RFpyWAqKUJf+2puanozzz6WSCttTOtySHk5SBmRArwyY4YQ3AXZCym4btBRaBSILHp/
28jiImRzeTgg7Zm4YsQH05IJxo6ao7Ur4QwDsnOEOObfoAOBQ1rx1Uf2OYO41KdP9nuRbRyBFwwb
EKyYBb6zcJu9qjBjwqonyO+CcGShabGokWmH9tvFi9d1YKsaNWAdpz0xh3N/bPa4JMsdZf+WvOZA
0lHYOqN+v8dvgL0P5gJAjc+XAf5TIbbbh6Bn58/mMA2dGqD20ns9D+jyFhMNKV6rOSSuKJlwsDzo
Xpdysiztx9DUUt3DOOqy1lE6OiJajKIl/dgvj/ladcIfRih4cNleA0Ds57a75NICEwp11TdQFW0A
6H+vSxW6hJJWUNHG1X/qmfjdjiPfJB04psYY0Yje+mSPd27xS7tN4HJ/otwn+H/v0K+Dy3NcI131
4ZOm58nKT/9pDTggg1X21vTCIxhJTb3/oo/o6i675V9IolqD4ds/hUhZpiZHUDLRAeJfdB8KHc7w
bcu4YEP+i7vinQwThDVj03pTL50WIPIIDZm96AsAQ/NTfnRaAYxNscGzAKyTT+3ZUg+XL7zBUsIp
cp3NIV7BzQmUc22J7xmcQbGJ27CoSWUjNZ5Sf1bJ0LmgUfE5wZrxN34Wpzb7TZFnqjKFo7diYH5K
X+/nHkqx59vf9qwTtyOG0ddNN/SmxLZC8QQz2NAQz0PHHGDoWn2Odf3F67QWEGqiN+gltDx+Ucnu
L2X1i7KFs3fJ7VuKumzwvPFlELT5kW1PLPR8ehFmvfTgR8zF5eWdscByl7NpWRqdR59cE3l83png
ZLWTyMvU4TFf1c2cgSjvNuyJR5vJcJk5c0XP4uQyiCCp2qv8Qg8rK7komk5HK8oYWRzemzETJV5r
bMIxgzAfMa9dbsF1R7ynMI6vgB1f9JHc6/fJpJFblDzQaz4Oi40d1XGe8xtgMuSaYBmPCHi49oM+
dqXC2F4LrPnjJP0cmjfwwgDDJE10YyRwQsG8KYhoAXGH/+lM6uxdpEZQMKv1eizMKYsklcSymsoe
DTqEq92wQwL0kYGM69aiMyAetX/5Bv2FmV0uqCKjq5HU7mIWc73rTbAztZ7gvQeUQaTHfMIyOTvw
DMesjpJKhTFfPLNEPyJWcwQQhq2yj4Ih/DZQ16GQvYchbaXZGfhrymGuf6wWYiyi2zvxvFQG8DUj
eniUgVxlA7xYYJID2/66xS4ukl22No24Rd8lR/YJfnGvD+vzY515hIjTnspznkW5mb7qfvdAszKL
GQDgqam2jVmtwE1Nzv8axMH7AHIGy6BmPX08EwrgQE/d07hWA7VnuQPOSaQGwogg8ZIet2ckRjlg
lmqLATIeJ9bv6V4Y2QXzMxbgkafRhk7kwPoeKKl+nBI7yV3ds2mA/KCwekmkOG+Rnu6GRr+91eKG
c6m1krZ1S6gNfBxf8B3TPN+Lk1oe6KMsGlOkClqcJ0BVusJjvYEB+Q7W7qlGvf/1IUruQYhZj60m
xTjHdRiszO3/EmY8q1RaBFxP+mJftgdnSpU6T/x1faImPK89ZqEURKJ3Q8zP3AFXTke5gt9NdpB6
8S0laByo055jcp+5qN18G90IUV0uZJoqHLv5brrHaTEfOyi2s6OyYNbIIl4Xd6QI9QSMPoJsPouH
iL4OVy2IdeURz5uvg4gjkV5F9kRJ4Wb7UKKjv5XhuGcJWwkBPe6/NeLTAZqCps+yhb4GOObOFJAF
ttH49WgSyypeTjGkdm8xB/hKyu7cLlJzXd3NwE+6XYTYEwc5aam44t5uGyc/2cvOAAKnqCqO2IEo
zJ17tdXwE93mj4rS/TC4PnvVbwcP0CoD9rtNUCM9E/6tqyiV5LkCNI3nkZpXoI5cL3a/YSBSDxVZ
PptHwp2Z7xW7l3nC4D0e0KShMcbMC4hrtxd4i+wh2LoYz8RFHtpQGCUcuLO4y7DAseRS5PJHrJn6
xVFmiTKtdiZdS/KTvyH2mBGcVJ7VDs1DhnlqSsq6ImaySWuO960AJXkMDXgd4nyKPXdSVF5YYfyi
K4miq3VJA+/w2TYS2og/hp8/XPaguCFsAl8gMPTzT2ys9Pn7n0OFE3vYj4TOvgOmf+uLrZx+80Os
4BAmv/mSGorVOvodA6UQZUbmVU03hddHg/bZ+tLLpR6g4TXLOESdVH/dFZ8MpNPi1EKa0zfmr54m
H95OokIdC6v+WTjsSLke4NuGzJuLE3pmCbDCNzZmTH/tW3jCX6Av4ure7C8HG4m1QMAQ8TD9LN6o
7qDke6OTvwT8u7MsygyclfvTToL5KUak4NeSu94VHWvV+E3hKuydXqGPFLiFwCYib0YPoBvOV9mU
0/E8Rx1w2LbJYcI3LRU7plDjZfEwtBzjN+JPysoVQGUUjrSXyQfZw92AZIfU12fI5BqJEmWNCMRz
GXQ5Tk5rkh6uMGoiB6RvJoOofMSHNOq9j1P1yYV3FKg1v/gL6IJQdvK8buM6YDX6A5IgkPBWq3DH
FVPdwGgD+C+0JyxiBFFDakwHJMymYDwzbjf/TUmDTm/W2+jeIbAIELiIGhtJtX4CzB1IpO8dLoW9
KWAVsmuSLCkh7oDjZxHA5tI9iWjTH8n3x+2bao6Gu5UXL4yE/3wF1JtLvA5haoKfxFWL8bPQ7iB9
yRvsCVEoH0cIzalSSge2b9ddNuKdEhQthPCN2DWUUfezOIUn8H0kC0ZvE1+lC0stUyYniVQI0yil
VcHrbXCTj1fDyXuqswuc+0pG9jzdQPyDV96r+QnPblJOqeoh6p0HyA63jtfBfuqW2r5j3lRtIyUT
wD3S4yFlR0oXaNffe8txdJsX6ghQgwIIkZlKKhzrCHjZtqECv2dAY7MKiZ4gS/rqCshLSTgBy6+Q
YRGtiV0OsrqaT5P7YAg4FneM5jIkGJAYqGyrC+AR6tCWvHkVub7VtagTQHUFhkuwtBbSINFRBay2
AdxTo/RcVrXZc9vl8rYbWxKx97A8sEIElIvGPswSO5Y/+2K2ZOrqfZzhcNny9VHTX6MXlVI2LJdU
3YM7ybEYFWk1CsAOmuA8J78a3bFu8ZPIuXi36s6wZVKAVuHu4LPMvdGpdTwuhG1byqHgAVIuKwhC
36zorUbtJhK0Coy4gKbIa9z2jHrkGN1mumsckiYSVc/iiRhX9CMce6G1KkHZtGnBVE6X6NgHGFEN
i81AMwhFJwPOEKMXkW7zMG7+VSaugSHyqlsOxFs7TeWvKDqEZZWwdAEc9Vq5CbI0/VDii+Jw7GpG
agiGIYPI0WtKXlpVkwsd3nJGXdVyvmFQFDA/vehC+sAP2ulfD0Ywm5vDbIeNKTwjd3jO7sDWM7Cf
XHlSPFw8eegF6utCAPJBbc8yrnq0JP+CA9s3sOP5GSMlCG/XLH3oZN4NF8JspmLZ9MRqts+fEQmG
o7/kqGkq9IupPYEbDpb6h5oS9mh8kw1jLEEuRg0qOSzjYwUO03grvxf6AhDJCpdgjFk0YIIlCVmY
/MPHiS0UqvbQBotiNbjNBoP17k4pZ9x7+w3YzPsYm0TjQjkDyySSx5byjDD5WPOFRFZ5yHswCSi3
guYQUxHJPl5+JlI5bo4h0ZlRm+1X4TqAtI9x1nA5mkOuVNN0EYaMmLB56bwpAe5IyHBpMNYI73Gi
MAn2goQPmlm2ektHuC09kNGn76OqPgapXPied7ab4t3AkavZIVcZ7l4iqmj847twFMCn72AZ526l
5cioJg3uJV66UON9yBQIY+YBq5KSm32ifIU9qz/SXxamVvXbuB/8n7HyQV6E2dcDTgD4rPKrYLQI
7wsHqkqtCAhZ5fMer8j6d6ynGh/jfWqDvP+ziG2HljDPtpO6HwQbV7iuow8ofvI5cdckY01A+GMA
b/iNIUS/x4ZxBXnABCZmpjzXWEi6iIqLK/2oXPgexKf8zLRz+eiE68jDybcC212i1SX16MYp61Sa
a9V404a7uxX09X6dvuPO7hEJmawcR75kMliR7dbPXXrcOxuD7wi4QPCKKWgCcKXyfiGJySL6JjGM
JUZNhD3f0yLQT/bB9lrVFPDDHuKBAtj8crPaANP6oP88v+Qzw19VvTjtydjGpeuFOzHxRywSkII1
qonphuE4UyNC4uYC7Opk9Znsqfwi1LyiD4YY+04evvgK5t0CEbeJwBzLavpLO9ypXM4cJxWmUy8+
aJWGx1QJnuxivxaHaqmyZUzzmNZytCI3aiNG/wAfIoE4zwH9poU3v+TNvPGeCy9PUed3U+JflFl0
lyhZErmPfgob2NTntoFbnansCJXpSMjd6EQk+UYDnwpp1ekJefUPwZuTzFerHxtVHALkh3A20dzt
/R87JMsUaJWT/Qjf49n7QTpktj4FUGK6E6gFE9fIqkWxygqaiRtpPDAgYUFENA13i7b5gSumqmhz
gH+ZDRTNWqNjg+wEbN3vPvgDFLgq/FWX6zNMuQgIy7u8eZjGQk3Rr+TlvGrmp9KtonsTBEIa8iIs
P94WcbxAMzPn+GQv6603tJuU0WHSDfmxVZpZcZsUrvl30HragJ8cv5ImEj0TRMF0FI9fLPIF0/1u
25wQtMnz1+lX1HSk2gdrk8+1voFVM7m/VO2V3uXF/AD5WiMoCiejSJGrfJ8egJv5gPeizrjM5Akp
H8De5kaVy0pcXdwlMoJyNlD3AYXmbaHgs88XXSRVY005aJwrozwEBkvNMjGWnxpsgM5zITdQmg6n
ipXamvzXJsjbIUkg45tK4Gz575sZwKLUFihpsw1T0q3gLOgMXx/iyyn8nVy9ty7hOmSKQjpJw64j
+VT5Y4G+gtErMzunq7B0hM2Y/Hjc0gGoeXpOrq5NUnrhLHTfjpcWkxcC7EOC0gnZaxIuB/o6nT8O
X8uTwAMPSzLD7Mu/XMmorVvh91kTEkASvSFYoh0czLbPN7rkc0I4dibkn1nG+jUPNCaCqYpB12Q1
rNnJee7qPnK9DWJETBEVNPqJ5C/r9jUxKsgOG494+YnX67M6DjnR9dogPz7OrqJlibNvy3gKQ6J+
3B+7s3DQEhE0RjJx1wg7p38sNC0LYfpYmRtLbPaaclDNOCXvzg7EGX29pm2mwnawgS6i/x4tfuti
AgYATOXGdjSMjhWBULt4uRj8cqhl8JcqnpZrBA37FB6FZJwpyyqMKEbTkGHrabBaAYDDcKB5JdfG
XrpUjPytTvehmLdetcIWpijKMe3Yg0jZ0xxXnsSBf9YTsCn5Wa82bLMno75IYPHTt43Y1oJpKvlq
dj6vr4B+trly5FrsD4O8eT/LFDutHiE+iSbHj+nIPOSuR1A8aHzlPtZiMWL1GuyvMTawlda/23zw
50Mm8sR6q5UXiy5VMFEyOHP0iKtSd+wHyX/KCEVMsRsNx5Z8ANxqvzRvqNwF4ryGQq5921WAb2rr
NtXkAnQWKDOX5Tw3kkNtUR4BCzFBPodXUKjf2KVNa0yBKdr6tW8gCP5uBr+RmG2A1Eahf2yP2XLZ
0ftWIsTdnEUUTpNonUHHvFNSez8ASV2kiYDfo+vnHk9QbjMB4pQMUO+tJ0OOi/6QabLxHoL/GE8B
KvOZEoKPLSTZD/oe1TcC2s5SPCMjHz3Jlo3DFVzMwWDfrMlo2luOp9E+6hnVq1B+eSQ2NC4SYkKF
BkzAKrUIWP58RaeEzQHBO5FaDddPErst5tatLbjC2iO2b30pALmZXHbxr4Gs7at45CR2MWvaRyWg
Kc6FhZIa9MM/IcZPsiI3yF0jHAYsrd8LiCV38Ig/NjVG5Oov6yQDLoc+zYWvuSWfl0H7uCOblKMZ
yVKZgYqYMWJTpUdu/p0e9e1lJ+JqNzQ+5HecWdxNbPL04KIw3DZsw5ss1A6JhHR+6WW71lA61vUS
IO2BGGSjYyAn+JF6IDjJlSxv+qyWPw1RxjEJCZ5/8OX9qtgRHSVoj9HP8KsAgjm0EYR70Hgo6b/b
rNyvoM4omZgOs02qrxkWn8bQyqJqqA+iT5GbSyUvUzQMbZCM8DXpOFhUz3avpI7cOMDRwZchj7EJ
pESOa2QscEpRhNi7yugpjcZXauVx7FYQLL+pwPkZKazxsAij+L7/FFv59yeWPLZEsVNkCdmcbilD
IMyKSZKYWo7wrVsX21c/36ZJ+94C0VlAMv4VGv48bVIQehqwNnbJwNiUxwidNlNOkcf1Q04m7Cqj
LIv30xTW79KSyBXeRBGlL3hn8AXekrMYu28W2vR++oqYNTAiyQYabmvWlq6IY9mJIS8hEpF1VeS4
GMNJAJX+VwjfB/KAeS1xHUssSyIsk/311U++5kZHEcdKUn15Wn7koCuYdvVh8ozJsYnKZIYdyHqP
V37V7hzhdScdWBQAS+yPIsWvzCvPCiqrD4zPyMAbDdtOlnhAlmU1IUYyQGaFajeGez22UHqdRzGw
i/jMn+yPZx4zQJze4tORk3Gd66z9YTU/3Ql7SasP9PP0bZyN4yoj/HXckcWu1GHVZt1FNks6nDzn
Seiwy8PaVSCBFYOyjRQdPy8rwGP3s9M0JMElhIT0WPh3zaYAzSW3ae1y1eCtmPbAi3442clwn0yA
Dvm8Bcu/4rYGmWevigaYRIDEGrwj/bfI0avRpFQsQlsktH8T6G+geSii6bmAESevVUaMjPtC3fP9
o8gXBW9tSf7PlhPWn+PG6pNXz1KH2Zg30qKxt/Fmyqmd4vtp97WSWYaEl6MUOF8LZ988bhRSXz2L
+0x0xoDhB96aBLRTF/4XRKtW0kpPLPbWKyInYLsec6Wb3iH6rQrgV+3moY8ANPHHdwvev/1Os5uq
j9urnsSAe1ADNmrjUBYqU6IBvB/qZY/GinKH6OZGSzK0ZTiYlbTP2wro/eHYo64b3LnkRrpP2oIp
6uY7bqjGbCOK84EeN7HXQ6skOGdbdONEiW1hULC+D7PgOliSiifk68HkniXlwGKlqbTgUG+k12T0
eOliUxwIJNmkDb0/u7lomudXv5jhzH5HPmcoUtVY2Et9TGKZ/NnkJuvkJL+cvmdrmnXqHj8u88Y/
bgs2wgBCAXe8V3FaWdVR3YU+/lP4pMkFclfAjqo/agifQqFk+Xl/IyEHCTAqOLS4dstkeLlJZKK5
4pEz9+jw+YvsZQlwGl9EcCIAU/jvI+z0P7+hz6Ow/OLNu1BM7S1xjzxE1SAG8fqumvw4Gti3LSkW
B5sk58yht+216plaWK+bAV5Ky4kNzOOqK7LyoQpBc1KbNjhPIAwInCOTHYOB7Su7RFFnmCDVNYLQ
OD6VQIbUaQcoKm8RxCE1qNhIbf9VpQjWBhn4DcdS9XKRK2W+J7tHzCXWvSV+DmQGbI4J6KpETz9s
Ps6pvBJ4/8kIvvI7Q3MnPNfLvyFdpF/vXw1JeFCsaBP7oj1+kUgbrQCaYJXaU5d3VAWV4jjQw2+h
Snz/81g4pEQ8NfNBgqZHNf9ILEIbtx9pdej155ZDIOTuMiy+Ie4kwdMKstrZYVASXLYOkXnD2v2w
fZiPq6ascd9Q3oWyKyflyjjrPzFg5SuTv4aW+6FczkO9QrLZtza6fDJIx/4THhZlas4rJoCTnD3p
pAUovXtibCjSsZolwpUpyDiAt9KmVR1X6X99DwaBMW2tnvmR618Gm6kvVx73utaZMRjYJsIi8uO1
v6rb4et7j7Rc5KMGJ26ctotjwD50iGCC/alQO7faZxeC5ARX+9ZNmjw80LiVl1Pzm5nLHphMCER1
ZGVas4UvdWU0SMNYMcHGTLMxWdvLUFO4vh74hlTUl3PeXY4AYWuyb4lKS0LfiuV22CAf3ZrVTzjQ
gmjZ0b6WmtOnfN9ufxVjnzGo6iLFH0s5sQK/tJVf9CRjpXzAcNivTLYwmAXLy/OGj9XMxQtJjNuk
jshGWs8Vj+LCx65Z3cKAF2hwIEZJmv+Agj0JGG+YkysTk23YaV8nU4SK5LQAlBUIk5NvJ20C9gMP
frTnKCNeA7dJ5VN+R04ug2wYcl4HKX5eZMWSl7EcLxd9hMMDNfRoYytb4dVFntjLxbTWZSgtpBX+
v5E1RAsgAywJAqhHZX5ZpppRIyy4kIYpp43dYtz3+cO3/bcjtpRfS2HoZKeO21b5VoTdWXuqDF60
qAzQNCYfjyvRNKipcpp5qik1jJLV/soL1Q/zzO6eHDxhQWbcwk1BWkyEpM2RfjocczhfxkuEGJmh
B4g5A/SogpRwMSoupni7mMEG8nt2ICc18kFuQPqpVS8QetLDOgQyMTd/8Gu0CpsNoxE+COrX5YDF
/6pSlFaHkQOBKzlPQ0lBp7mlijclRUQOX+9qM4jPG/FVf3wf4S5IOu5LuxzeGE/e6ddAHGjKpHuK
iqxfrGJZAr1Mm3ujjAigwAi8TCtEWHLGCpPa5gCIK/kMpkqKKBVoe1gr4XhY3HqUlpkC2sAaJgfb
cf5KvFAqYrT7FQ4G9pmfezDZPQgLeUcG0gat7ODjK/L4b7mINK0x/JmPi8OQOJOAmW5cvAPC/bVD
aoqap4EqLR7+TeVQZ1XKt0Qlwp6LPRJhzv6noA8WeLOqc2KrsVLs3ATVv33aGEmb/HDBPM5u4n2a
eO3IGpKc32+bbSTe7146t+7KHcSCeH9FIry0tcAb76YxCXvvhA8A+ZW/PAHKzmwaEJ9OTvp1DtZB
N6H5Tr+mA+T0VP2M81qFfBYYxBQTFycZMCEO8sfVoqjfGCoTnnfbXKHsdah9qZF7XHawJ7wyuBBY
wqXWv1sRS/1rP5CcUPoQLyLroECDK0OzqMqNYZnzMqlVjG5a7bPKrdJerP+uofljDpC4AGQBOgXd
rHfKYKsBiCDqs2kMDtDColFq2n6Zz5hrsIMisdM8Dvtc3OzFa6VvT+bkvUv1W+G0GSzJJRk4B8j7
GFjXSzs1H+8cFJDh2o9zp0na2+EnpLLjC7clajwzwXl9sSUuAf4igM7Y8Y8JkQDW5gVYHAMOA6qP
Nz/hEO4TPiGOlDkg/U9KiYAHODyElnV9VSry6M7Ql2bcCwaMTXe76db/zzov8Sok+HvWiBOYppjR
8cJ9oSogoR3UC+ZvbffkSY/UiXxUmFMjilzK/DVsVfhmAymXLrva0Umuak3qcfTHXmqNszVZDY5q
PiVRyS8GUI4rhV+BGAWsuXYQ027+p8OehETjAzuxayjFFpuAITUnFexXrTfGMO/+hAL/iyX3Cb4h
9KBbUZwfodWiHltQLgF+6rdgSeJKVjQhO68/I2/GoBHTFy9BLDeafpwnwS1tUH0cwbX2JfEs2XT/
0AZ+JoPn0I1MwXF25VJHati7jFgXVNfvqreTTIN9eQs3O+5FjqNzRzTW92sqj/oqPJ8Bd1XSOQKB
fpg6JZQ0JnUKe4Jp2xA8opcCyE2T+f9mSwS0rLEt0IkEqNVLSfOF1XF3vsMWmLivn5xK4BZmcwi3
MPrkflFMsVSi45+0o9QJR9u4kaDKteHVAzWNY9NGVSmfOleyIrgqDCVBJT0Zo8zWQqMXW+nPeFt5
6pLpIQXzkQUJQffOR6aJ5yhnbF9McME+eWZcnt54mhb+oHK5DMxZz7SSl+3BnkgxATd+zAEHWtpX
8vn6ACIQVe2hLW/aP0zX9OLO+Jg3wxddk6PZE8ho1SMTMpzuYqPMppzJocxhE9cC8861ywnxYkSM
Ivp8EbhTUIZkbjs8tVsnqqJxkj2j/0PaZ1+fwPyJXNsxCgSpyMW8Hy4Mht4YEaFMGxdc7DbmxDKZ
hIiEZO9ioiSqRv+SOkZZdsBQTqtvPo4Xd/2g2BySc2BQqgl4KDs822jUlaYcDhV+AbhDznzgzh9U
FmRWX7G0eES0S6QckPD8ZxfAFoSjwX5k7IT6FK3oX7rXk/dR8aGcBCqqSheF/WHZrW6pklXgykkh
/iuIID7a4lz4D+X8YmZ2rn0Gt3Hn1Q0UZUqpDe+opXugQ3NB2n98aoOrfbt0BVlgw0nErWwCJ7SG
mK+vM1uUpdzoVz75ogZ17fcJ2I7Ry7VBOSjVcB8fdTD0PTwn2hsC+ZKaH0NrNyFU77G7lAbXy4pI
woOvyifNBBeiNZ5AIizUopkYYYC6Sunax508/9Zu1Z3oCq0j5qg4x0QAuGFEeEchK5aDISrYTsPS
5yIkPHa/CysTcVSLSppOjFZuvk8gEiFlBUlhVPZ3TZ37A2CTeMb90xo/0Ddv8T/gf3HviPTEJqhw
2B8jz3QyU51mr9AFnNCYUxEEys/NzpYJdl01K8IiLmVZiupGwbzndgprXhNxSU0FfvS36rQPEhoP
OlhMoyATcE+AWrJlEPJWaXOhpUquHMpSg7QzA59RJD3VlmdPnatpb2Lg0FpWHDoa95cv9x/r3/Gm
Y/0aYDTdGGUukkfNVxG4oom2zfO3mxdhR7DVujuZWL1QXtrOuQg/yQu8wUqIR1ZF27+S+R/zCX0F
q7SB9mQoJKq0euaBg7TNQJPcihtVAwh/jiJ2WF0nzgfCSYYa+htdbo8h89d/+eO2k1jcQZcvMq1I
+sWyboFYg0xFovHCaXh8XN2yLECV2b65wsbrpCjvn9SYlcBjtkxkoyPOt0fqbQ8Z24myOsphFzAl
dySVCvayg/gudxXXt8+ngBhNnZ9qaIRnGe2OZCDtAMHFnO5hdlDY/E2qhOk+qcUB81LkhWNmCIEW
crmV5nOp0PiVEIlfZra6iDkYTgmo3L1HcjJRsV4h2eeeg3QgLj04eX3FBuyN2CImWvzSvhjhfTZt
5GE1bPq3VU92gaF0BhOT/KjM5O9FMDRg9qGsiQCH8BQgEAGbgymAv5ijTqP/h8/ivRHoKXy70fFZ
SnKPPFVSPT3yMTewQdGtd8weoGTKvO5sBhaW3ECDHR13S7BlElBhMrfyP2k1Jip74Itr7B+5DT5J
A7iG4OW+YCkUzqVLtv4iEhyjEvzjVdEtYOucs+bbyy0t3zt2HOChj7+pE5HN8ELh5xhwr09KIs4C
49c+ux22h8ScCIGdIWJv5Z+26omvOau7KzSL2OSLt9vljh7hxzscenclx8odoWgExymccTS9h/Fh
qqlVZZIDsCd42mPRDKtkMF1miTFcrNQzblFxGbpcBjSQ958kO7YpC5xiU/FcQDw67e/HYThHv+1D
2W1EAB/QEYCrXtIGcc8/6V7BSo+hhzZ/WYWyG6j5v2GQWMQ/UhEn0RstxFnomLKDn0njzhVAT+Sr
O7lLDjY4TMA3Icolc/J9fBn/ys4mdjVNMexrBFkl4kJiwe8HuZ+Nnrd9g9XFlzLzyt1ZMrYEnMN/
SM2PaLjaBtOjG0YPo5cQzjXUwFZBB4PfiDm2sZ7Bv6Ii8+wbVFcWBcGvSU6xMIyeVqePTckf90/V
oCN3c02sMJ628kiHbJ+IQN2fY3Sp4JKoROu9lEsIc9G6YtggoW6nGSVkVJPgseIcbi/bwfaX8CGS
eE28PnVY5ju44SRrc93YCaDjCUWwHEal4eLRHe4EnoepeyDnXCqrMp12LUpKxnK44bEb9IHFrwfq
sYbCNoder2D7MFA2p+z564MdCvamK0oQoicHGdX4prCSCpWB4f6Sqz+tN8m7WdF+0vixwe4WjOyd
DBDCRlSjPZOyVkJme9tlpWQEeLz6ry157MEeXqg5KKMbj4JvmFr1l0d5vTfwKvPV+78Qs3OcysiV
IhPRLlCCkT7br6GRzZ6toU4quDQlWZTzmSP7D5G0LYSIeoagC+b06YOJoIAStYiKEI8WMseFbgaY
5J2/4NCS6aHDtasZDJyntOmN6f75dlL86G9gpkt919xhBHDTb5HAEnX0asZsgWAT3itORcbbYvuC
TH4e1x/Zsgs50dKAWjwb8Off5XxtyHV9QV6hO1JFDc/HzLF6eCT5LnygfyqED5VcI1lCvFI0h0nS
u0UVg1v7+Iw2mmGFRdB0lwqXLJPcSzmioPMBeSiOF1xhg/JP0KczfQPibl6odBEFugtGzzOeU3Sh
V5/dd64G9hXUKRmYSy01WqwikTxtPXhg2xI+908KXuCs9i1/tLXbJEwyo70x5ar0N/l0KnHqwtRf
XfzqImJgRkurXGPELdym9oaujy0lW/WlRvVrMyMua0moSzp5QS6QQFPNqlykQUGlJUyjjF/BjmFt
TEpg+akDpVP0hme9On5ayCc8A1Hi1W9eV1Uz7RTfCQlgvfeP9XsCn3PSKuHakeaNUTkQj2a9GZ2B
lssMLIaFbTpfqCBzZO9lNRPhSMRP1kvBKljHSnwKZcZkq+fL78gbl3AxqRtWwahAFP+84/kHrm04
0p5FhwbtUbHEWIwOcsPz3H3WoJt8bosGqUk6qBr8P2jaH33UaUO1PSR0SIX5QjHUgNbPjvVX07AH
ADZDV0E0blzLgExldSMvnP0J8Ca1BoM43ii9REclSlKgkG8qfJecoQSupx+gR7EDwDoj49WGhYbf
NIVIe7WBJ9+uFN6wOhKLUijJzKUNCBD/GBFzwjBtr6ryNkxzZSE7QK//3a3lQZUnMNry4u/6i+2L
q+ghhPNzDW64/5DMgGzK/3xUvyD/O/tlhbxfXtMvyU2rX0F3huMe6WMRwLsyup6kQp/dfAheYx2F
vs6nY8OYdIf0T9OIfuZS+Ct5vmM7iU8Df/oujpxxhGafqx2xjbrH4pUsvyV7Jbw0qea/8GBm79Ma
eGsp2GGThmEeMCpqxkB0KHs9P98/cd6UoAzbV0Y2WC0T+CrEm03LWCpzuhoLF8NmSBY54oQ5CJbK
BQq6FpRnJm+GPNBApBTMd6dDeEqJ9RLy9WwCiuLgjQVeOxsim2GfjAD8NUI0Gajx8p7kqwxMQe5z
ydYc1M4eFJrdTdf2yXIv1n4t8WBxdPx4A9CEmpO8Ot4B7ocw3Q5ECDcFQ/z23JyaI6g4J/qwU+Bl
7bMrUntCARxkdhZvBnKh2V6nb0PhhDD4/1ZImUSD/YsZze+E2+s1MQt1rLjP5Lk6Vtt2tnayyUtx
ZlMZOSK8gX7fcS65xgc7b8C/lqyqHMRDzzFsKk1lblvoEuX2xHrmjZArmtlbUkMllMDVbWxDyLDY
xUCvPeCbsDoOONsP2MgHSvKv2qcvyTMR+igorap5lP7K6nRiCb/0IsvueHtAGDXLWnI0z491Brl1
i3cPi+/OJJnGviO0uJ6iYveUQ6Q/Txdytb3JsxveuBnoU3OT/tAmshpbb5NLT6KnwIQYVYnullO5
oFc7zZtx6AQ9zLt3uaRq+Bk+XWRPtbjX2XV4rfjxFDHj8Oo35a530oozroHcK48N2yM2KvY+UorN
n8L6CUrqVpWyEpUEjEMZiLfsPPvsvrN81hFmbYvzW4KTj1qF/ap/4u/fPT6aIJ3kpht0cYZBaQIj
fljahJpr/FCoUy4lOoLIcucgFHVNMsq3mEmLMH/ZPQpo+6EHvzxQMKbdEj9XQFfDgfhNE04Mo9JF
vOuTzqMXnGXtSuFfi367jCZMlDrXVzAxuGDcVY9//jqKiqEr1dFdHpFJ8JNL+j/wgTxcFxNhEpBW
XuryS0AXk+fgkaXGAzHn+Z1eyQvlT/2zP60c0Wm4Ze194oFVIQNM8pQ/zuo3ICzpwBjH72zS4p+Y
K+GpM/i/kCUXpWMBfV9nnbRuHpY8BMvU33Y0qBFPItW0VXEGYdCky7LFxZfEWKmb1Zg7ASNlqStA
/0zF9l2Rw+Yfy5yXitLPbl1xmNsXwh5HolUOXJnRiQeKo/9HIgFg2utJO+GZX+yRQsVGgqblgIDM
E/tMgHWm4J1HsLhsj5Iq7DIYvitcPfqmjwqOTX8594VTHEgJEmlupwg5yR1/CG05NkRUtB/1nJVu
s4DJidSfmT1DOeNjEj4tOzvRAAUDxJaGpvXxEsRka82wmd3yMBczsO1O807MDDMAkwtWRr1VZOzt
HehwEgS6TvyicKSp+pI2OLq2iVs1d6GXQpBixSR3OpH3iuv7oaZZWBbX3Zyel43tEQ2oU3IO8MDz
AmeZhHKyldpyRYsJPJbQ/K2e+F8ahJvyV3J0vRyVAz/B3S+xWdCDt0lNssvNK+tQ0ZvzPvfOZJf+
s5jLIhntvzyI4uw2aIlQ25eCDctUfgEBuRtaamXqoLisdxZCPF/W/zfu3BEqYkI8ii4xZTZQtRkO
HaESXSg7sCCFwebez8mmaYaaC/8N7heVjRITfN4mHMMLC5rHtnV35R95o6m1AuI+37A8TkoSWOw/
Ksm8iMGgodbOFggda1oyvIT4+RbSeDTgcqdRB1JVZWQttg5R6XSoZI+MI1T9yvqyCGP+4UelsddI
5e0tESgY0kPeWI4zWiKvmoVwORPpzoJ7Zq5wqSanVEX/wA1hHKEomvN8PzM1wDGPFanzfPa/I6en
cAWzVZf9ZVUQJJdlLCgJGzOp3qlBzibEBYRG3QBUuO6oFbiqMgMILA0AUSsxrStUrbaO7e1DznPz
NbE9t8/lQLAoKCWElHDlQ8JYYTrIEW5xOQOJrNFU1oz3XE5Tcf54n+UrncVL8M7mqhzMxQeyG93c
Sh+ryvPddB85LcPPnF6KW32BZjwO/VdG/FHcIWFZ2l+bvhpaR8w5I7EVAjPvJzERkoVOn3zeJUQO
1zNo8czAuZ22fA3CBtjIUxgsKTm+BRaOAz3SXiYcp2YEs0yRR15IwQbCGDdpsS58xrJ2HlgVqMaR
ZGei7OeVjMdPF7AvtQfLS1pAMld0Z/p1wbYRZ0QS05mX35Ff6KDgu8YE4FXL7gOgwWbdYgfCcB5a
Lw8e3NWzRSYHakEesjVTi4e6nUQSC2KWfPnzyZ/UMTjz68vUy1lIGSmjIzZY6mkSk/SXBD09nGR1
XerpEN28qzpEBldjyxVHexvk4CawBla2Qrm7yjbNmgGL1P1bHKiRLq/tzKec2dQhOZBodbXqapUn
EVu8W8MzXMRoMpmH7iH6dSsZK2R+Zo2U+KagTcCTf+q7fEfmQ4ufSV5ChoL+ggzRURvkb3bmGgKq
tAJamjD7D+Zk9067NGrEGBv1UwTAbhJtBmYmvK8A9OjCU2eIvzhaTpGl3UUNcqgAx4hjIAcsL19P
fYj5i1PDGlNKyCMkJcF1kigu7gEONDgY0Wo0jB1TebGTEkHaKR12XcDjwGDea3Agv4+Yt8ZRUdhs
qkKTqjae8EsrTSZlxfULJ2MNA9wtoXCDgbSs5eVSKLS+kPkOv/QrOToEJqmZArfHaBmtHZuw1rMJ
E6+YM1WR3EQwYpg5fcaYHAo7qQwrrsYgP+QFY4KlX4VV8g5x/xP7J9xnE+l7Nu9IC+Gk1xWIAI4r
RF0X8XK1TZrA2cDID2a15gMu07gyr7QPvueqsHBKVkvWJKeUlFhEmUx+uHrkLAruI4lc8Y1OF0/Q
rvHh/miBENwhWSx2G+h9hHkDw+k4ftpPBhzle4P7Z9Ar2s6AfzmSR0HwIEcmU5ivSRZAQ5aLhdvs
uVjWn0GwBuQx23znO3CyqrGE+N5HiHwz+oHjg7n2PmMeXPRc3IUTDtIwydk5s9yEIDgVyOjrjEei
dQmRmv6xODVmfvmNQFkmvpy0HAiHfDiIs3/Q2G84Z3UwvL3snV17tpg/65VPyzaYlC/j+e2TzCnf
m15OJahmPJATo7PtQm3yGHsGQPQHO9eZHBXNPr/+veIQyvW52i3NGtKWbHeiKMV3jv8+TVetlaAc
i048Xr9SXT4yHphHp5fwtZrkzOyLEP3znpWYd82+xiPsS4F8JzjNU6p/MxSdQ3ZKUtFlM6clrFii
6bqhHMZ+iyqMRcRwRmxSiqymF4H3y/oqvqyq/hiGC6sY/rWhJX4vpsIw/Pu1uZr3LQ/rn2Vqg4m4
lZ+9LpqS/e42hV9Fqu73SkebOEhej+c2WgToKthMwa8NP62Wx2wBWdSkTdF7PXPO3KNRB+ftF8ee
U5879NNChhHi2HR8dgWfflU4A8GjZMMQU0M9S4893BvMfkLwVIeaDTDX/hTiieRYYpXUad3bVyv4
3j2wfFoW8eI0N+GCCQY6RhnoTcHX4ZFReEskEjy++oJGtl5mqx5ujPM+nApuKItReEd6TdftAbdS
A9JkqVO9bxZDV7p36p4nhVfOckLTWwCXZ6SfUb5PFBFskI5waSoZajp4Yx77dqXT8EQEwNEkueyH
eqjRa1eEF4L4aK1dn9bGECDHNDduIkdAvwExRrE3GF07kSYzP3Y4wqwvLCLSoTWaU11vaYaWb0d6
I3rYxT5oIX0GwHi6Obmfnqqgvd2O+q+xJ7XIyXCnMnmq5cxN40+ax8ge1nXYZygE418gBMdiFK+A
iUmuvLDheEqQAMC/LRsa9NPbPkVSEzCMn56QL7/UhreqLLFtBQd5efNF2fsh/2RQrgg1tUMHe3PH
Cf0WwkaCi8DeXMwyDybV83g39a0bZODzqBXv4x5HE5kw9+uQPU63GL/ZKKTR85Rc4oaARuVSTD/R
K7z9Y9H+c2FdacKVJTCKy0des6m8wB2y+9Z2AttcR4QVs//qQGUlzMI5Q0556VdxzEpZpv9KMYfI
+8SRXAsU8CQ+aNuyD47MmKYaKJr7KE2Uwa8HsS0d43RUMeZ3mVxV+mH3yvhpAl0FMh2LVNaFb9o0
lyPHPyvBG1wFZXglpdmrnfUbRNmF/M78FQpG7NxtpUPUb6zMp/C+xfswwXQw5n/z8NPlVS2Ji+Sc
6WnGtjg/eCRMQ7zkveBfnPa/lpt0bMme7q1ZTUrQ2GwgCcHOiOUuTOoc4zHAkmreE38JioyKk9YI
sAH9X4FEgeKY6PBFtPAVEAoz7X4usEh6f/OjLwtOVd5eIRRyPoRRu1KOGt5RWcrxl7IZVcUZ6JWh
1ythK0N5HMZBqvTl8S9l2Q+aVdlUYjPsmwDbIWRrf6n5RA3Q+q+HGvxk6pDlkA1U49sqVfPznUQD
u6+vDTbbtoH3Hik8xekR4leiUeiVz+OTzz7pL1esWT9s6jBpZZ9MktOiVJCG5XUzaEIgT9sat73s
dyIj+CSmyH+8+fdLrwtedYjhUfU+e7JfYk01IoredQHETFY8iYGt7KNUiMKdyw6qByeTJC6Tw1KW
FL4XKhEzEr12KiKP+pbcSwPe2lFq/MFOFQW4VvVNmMUEgWCJ4WI1FHm91PFc881jHyKiYGUECVnz
qq4GoRrXEhQiwh8oNGKOz2ngpzoUTAjCFnjE0YkkhXvekmpC0gSAHAh7/dbM1zr7tEEyNIenEHIn
SrGGmYc18abPANGmZakHg/hGixZ3jshn+9yvVslwMczA2Y+h2zey9/78/IQ0I+KC41Mt8axn+lc5
eJY/va0nA3kfPoqZGvhnzkbTFirQHW7I1iVE98IIzJue9BaM/Fx172PxpaicIbpD+1BfZcVrykAL
UfyTyGfdvqHfVfdVgesiX2Pqk/D8o14E0owlNBCJZUsnAU3amBfjBAllu0lmqTLMM/7RW5tFImgq
+iAgsKX+CzJY08I+5bvBEAr69dU05ODQatIV1jLJ1tEckrmSyAIwsmH3+XHJ5TzcTIUcqFpYThos
xYXmQKagdISRcQb8euXj82Ue72sUw3Ju02ZdrDGN0r2V3MhVUvwnXTPefYAwjVepDq1bak97BXBn
WhGAShRIcON2SOyi3MkZfSA3BWYYCi6jYYThZ50YYg8nt4OpsrZJmTJWPTbqUMME8TWUX4luHgbP
UVnVm9p3lFthXjUbQ61veXUAVrEUXkqUA+15Sk6zJW0eDgJ/6tJRhkg90HBKYVw3eLm8w8knDRHL
TOvLYnw/GS2hgjmKI/bxJQntG+QN8KGoMr0PIwekxSHcx9g4INokY2YjOIBR+iD7VMnZsx0HWNwY
/EutKhqW8sRdqVM1pd0gt30zhvhXq7xbVwDdUn0J1X+f8GjTFDrGKy8LwXdFAYGXpxucn2jgSCCy
1k7omcErKSiTLXlIq8N+8Zie8FXzrIIZTued/kweEecD7h2xdkyvkh4zRtoRX5CTu2NOvaK1hVqg
oXewou4dzI7pKiyYmce6ZIyVf3qXe4oOnij6igBqzenfzyFvb0yMOzbyf8FHVCBORRi7erqJFoMR
RkwLpJsJA3o9hMuUVjdlhYZFRGFJWCQMMPm9yjCNyks97p3NE2dAI/EdFxGSWN2QMfIf9TP5Wnl/
fCBgONTQnO5xBcCInfrgckeg/vrGTSoqicprxTNDvlLKLlL8ashrG9AS/DtbK1U/Pij/tJdrJRrs
zOFQvQdol6A//cilDAkilZW0wTM2ci1cW0ebtsWBDJwVGifblPK+i0r/qz0DcX1CBjX5Aue34IYz
xLHADzmDY49MFsOdZ3E7YDJhcjS6y2HUsi9E8TRb8SfRXKT7xTYXokCciYaPaRVS/Sj9YyVpb4Iz
5VBN+DYZdjLVvstd6VtEuldX5Y7kTylHyZNdXp0ztaADic9CqqQVXzLBcwre5ctpExgQ9Mg7Fzxb
9E4umIeOxGtgXRip1c3k6Na4F1/SWRoMeqLsyAWh31u0+57wtVhC2bI26FqoWxH2Tc2SSVasT2SB
XX0W/m9e/IYcw/Oc9qpSHCGyoU/TCLnxaRYRa9P7JjHyOS1NMWSw196WumrWI5rzduQfYIOnnLoi
5jZOpc54WLmFgmE5u4QcwZF4vgg28+u9GqOUoGnJZJ7i5094XOODBzRO254cNmVQpJMbNdXpSrtX
m7XNhDpukpmQ+E2+iDzdc+i87dgn3z9oVXT3ujhZ3b+Zm4/sWqBnJpP2We58e5S6EmbDucg1Gkbs
gWDdb5GDWphX2KtraTrwuzSRhydEzFhg9UNxfOZOa7Svooym4JMRXvEhONpFOUfVujc7DxVwOBlR
SOcUaKQgRWTWJqW0NheZEqeO5GOuUnlyKdInxHaOkDnkJDUSy8mle7SpVE3xp7FhaehiGlX1Frrm
rDWrto9WhtCGU403MvfK1m2uAv5nXcCtXIX0gOeEehS5uiaAAK2A+XEdvVmGkR7ylbFL9OctIxsO
mjx7x7K1b+3/jyDS+RBkkzLjnVBa0j82yHvLIhvVEXRY4lXsovhBdK5x2iXkb2t5i/C5pGNE1x0T
t2UDGRzpM4cb/lJXyX0mE5Q2txy/OUuVhRnnIY6+Jf5LWCAjryROUAMt/mBWecFQG3t6DlunDSR3
tIZXLECFN9GXrYD8xYVWFFHe8SguUvDnbo1HOkIIu7QMtiQYIAcROsOg96mTk0d3i399gskQQC2v
BWvW60P04Gm/fGV/ucW8wZkqGdWXetHsX1UZJt2kiEgUqBI2wK6LApUFD0n9nKCBst/zCZE=
`protect end_protected
