`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DFZ5WgRqjFT9lVyqK6nQpKgB80akrPBjimQzluHFLikgdYrj5bwA2ssN1ElOIV9nrvuu87ubKZBv
lnRe0OSrzA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kC0FQeS1WxNdMHZ6za9mILmkUWaq/YvbftmdmD/YvkxE9qXCzuQ4X/Kcd+x95IK0oLwYQ53mcHtv
EJQQ2fhu6R3T476x8WBoOkJkm/HOADjkpZm+Zg3MJSjn5sPtCsF4Z2/wkUlCmeZLLxI5OsYtWFyN
04svrx7Wq6Y6eU+BZBw=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xI46Pccjo8ThDecbCfZ+2ohSnYQOsnWr2St3oXXHpvwFg0Nu1rUBEPSQt4jcO/raYF0ZQvMZFiHg
KSyOn4d3AwPjS3FPjL+Ky0GBJMLNsYWxYDXZrfSova1B+0HzhVtGQ8xMO0ZRkqPilj00dH5Hg4rE
JlpIxyXjyhpSAWu96sw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bFmZshi0sqkN643qM6zE1i27VisWSU5eY/nwaA2zsxUk3CqZcruFM4aqqI7SbeQ2eR59k2dkeUTC
m4raP91MF7BThgpZc4IkoR8C7KjDTBjNC9NjnSaEn9In4SiO+V3mvFEDMaW8s5fXjZ3hyBENWPaY
9YovoxnXbpPQ5325vf6Yevh9YCoyIasfp0RqxFxjNHdXJhHsp010HvJMvimpw2f5pdp1k55zFvXH
pitA/aB/99CW3J+QubemecW/ILdb7msBsNy0/qeyv4b9K8OPKLNSzredgiYa4fGbHzgphZqw1/a0
AtorqDnV6AITy6RHzZAUsvSRnUvt32AY3w8gQQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GT3YnJzupabpLi+SPy7VFa7UWjQwy7qFFlY58l/uq4gMFprj7TNyCu1vqVseo2VwzEizHzNcK7kH
1GqtX3RH+CceHQiYgdfMZldAK8gWy8GAkdwVj7zmpoUaIt5wYYMP3SDiidy/J3PDwAEN5imFQH5Z
xm8DPpTl//MGSwXokSPmpszqyH1WYwp8K/1j1JkB7HsIBpkoWthkUZZanmOf7weEx5wMxJkQpLz6
VPQXudw3YQYkb0Sy4QvLsAhlnfKh1Vq8HzScK7btRBJvs41joO9hm9fSDvjrFzJ+V2KNNEL4J2Pe
TT3vkjsziFz9KOQXBiVLM0jyNcQUSQjZy4pC4A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y6LshsPD1xF3TdW5KuFKeeUs/lgXWIJ7Je8GJUjsQs+U2qvOsyNMAInwIkk16UW3gxJ5JaFc4m10
mmnHCs3YIOr3JumCuS1jJogRkVTqPd2+o+j8FypFulSA7owquJjLTt5jm6RkpIqqdTzK0bv27ruA
/K5EPDB8CYmS5HhFZgaGGk6Ka0Ip5SB7ivzUfwsRLUw1Z+K3Epp0FNgWB2SoQOWMDTdpQa71cXsd
2OsgR12rpRLx16Ula1xC2MWeKR16MAnz2wagfpVIn/dCyIGHHVYBDYUrii40EP70ddOLlwG5SErt
jE/m+WDVJygvfcEun3Ys/e1u+V1AzDx+vNxUFw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
Uus/h2WhOYqYiBovodvY4reCVXdj8MkqJvk6OurfbPvYT8DjZZLZwSk9W1al8HkKHKI2YzvPoyk7
E0tqf5G5zjBbkC8OGD+gVyXjkqFP/vLWRONyn6sm3AuwYk6xcbp58eDCZF2LuE89NJkJ8WDRicXc
gUYTemHpUc38CpP6K6UysTDE8mrp1IdYLKkerSP5Emlj1x59fU/ngWGe0NF3XacyWvEPgglCx5f2
IZfC4qqhoWIcVz/FGZsO3mJwwqdLUZkE70ZS+eGs9DqgsuKlhIPkGBdq8zc6BQ87msO0MYY2tMSf
pE7VWKWn/UWZbmNENbD+DeLiIEVMiejsPL6lsYq5JNCuuJK9c1B5haoJZslLjosTnIfSZYT0iugL
L9z8HvHQle7srZ5mTEzOTPOE8EVXAt98A0UFSKf/5wlwxxn9vBN8PZuXQ6EDQXHhJXUY1O34XmzH
LwptSFTndPI8KSPwfnUvwHn2VgkI6sLq5KgWS9Gne56fpKrb5ZgBaoWi/JJ/yuGzHNHaIeLlhU74
3OATXl12Hr+A+CRzry4eGSPqsLJOqGAD6QjkZKDYaZcd/rMseK8KA/tO2hx9zhu1BMyjTUUDDgVQ
eU4ltoPS8HZWnPEqp9HY4YGmKXFLX5/L/Ppt8BWLpMvoVTI8twbzoGqXAubZQP8DbjM3QPF0v3nw
VVUIybmVZstWuqC7Rvizbj/9jCMogs8bE91jySiFacV8eF/NA14h3+bZ283JHbDxFZolIINws1Sr
e1qncd3n59ARJqGCAcN6Ahqmgrmmuu47RRrGJ2Rt88/ynRAO8jmK3XO5eZUztwJPIL0YPZAT8QuN
YPOGlG2Lg/ZF//T7quK39ASUxz+zXyr/hwi/nQXAqiVyjjBRWV0tvw1YKKYVOxPn5Y7/OLjAtcZN
vyxlsbsWO8bAcOmDpHJnM6dQ8uKFLd3bRH8fIAtrLXJDlbhX4SaQt6wrl/FoMuNI7PzaXDP/hY34
BohHDE4BOBXEtgxk0gJ8jO/TqVLbaury8WW42i3Rp59DMfJReVQ1qb7OE4VRRStddioyqkmb/0Oa
ZQ3X5oQhg7Q+L9j40rsUShBrYc5MqFRO/SV7n4Ely6/iuuTePvhJWHeonFhTQ1TAQnhH9UZ/skYT
/4sypJr6wQOdKlAbEvu2uZrKJvhZFQ+V/7awKxtpzjKqDCJz7YvQkJdySCvXVBBujceVzxldb4IK
THKFJAeU/VOaBnvwELlo8ORUE3zGQeh2EBCDkdhbLjYFmzkT7ojfVLctgkfEDHAHzKeZvOr9loe/
thQ9Lah2wLNOk9DAjXf4PtEAHUFRERZzv8svk6gI2u/7L7Nj7Nv5aC3tqNBbVV5XKNtqNqz61OC/
NPI/HfVrCu2Q9av+X3PWM/pT0ioE+l/JzyOkUD6/xFpp22KidpoRJKCMyYR6lz9j0ZAG4ntze0/W
pP0/t4u3ymhWUlylDxZ1KOIPC9GVPh3ezg+T6Z9JmIGVOSqgvT++CClff9LReADg7IvL0hdEFKxU
AOQ1V2PPNbTLt8QGDwU7ozs+AomGTpFDCeWRkDgHXLVvDw8XSTkFy1SqZ/KUw18XXs8pg9q+PMNV
kGQATXfTY55cXvp9+1Z+RwqNob0RGyCf1iSRt9p/+aNO8KMdDi/ao8WhLcrEIfaUydmfJ6Oja4l/
I6y52k3KdLBbd2FXynYAsaEelv6UmNCHO2QIIRdFzicYCGAQ11tBt26zzQvIdP4piJoESBoChq0U
cEhTPHxPuHkp/Zxb/v1gSCxj4MGj1kj+8FH2I5KyTwf6IwY/1+koepfup2Mp81mG2hbs3Vy5VF9C
zf1FboUnK5OGxM61dFt+Qx9feJ8Q1Q6BVHr3HOhGdoFQd1ZGXP4nEYTWKWmIJSCNbEPXqrJlPSp5
twYKdYHHSwr55mLQG7+f3mmpHdvjMKC5RkjZV6LRzGXvlvd+/fO4nipIqiiF2IzCDXaX3Vl3KlQz
z4A2/dVOqGXPEW3RkRX44DVgy+IhvBjcVeB8PBKoW23Y/osQEh17gUntzr/feDtzlXFp8XRUPgfu
ApcuoYHR52iAghfiOeTk5cr+KlNRF1d6LXPvxwrUy8loF9fnc9lkvsgvB+hPnUzrSBgFGcWKQA7O
XDu/XnRtUBSFwMQEnzxmNtHIEnnRjgeOq5oXMYgoX40pAqdMW+4wBxTi404mP3xCgLs+sq6w1tC7
JIeDzOmx2ognzEzLOltrpiqSU2GQVYNpCJfY+o38kc0ivz6RNPYOIFCOdE7o2Mw4TNm6uSJVYZoj
9HVE97cM7qMjsvoJYH6hkgrPxRBdT+AUFKjsb7NCx4CByB5PVlQuRbmIfu0dl4M25YVkW7pdT75Q
faejNVZ0MzICCSQs+A1JKHH9g3UpkSHMtdnc2e55n5KL085HkLb2rceex9LyRwG3+exmvBI5sxED
PCzJLP/5+jq9XSxaK3hzA86ZGFs+yJCag3CogAwnw4D98r6zyOEqRPK+JQKFbcvZRddm9V8gdEwJ
/Eu36BtReNrLlHtsBUff6yANfHb3HDJ/Suzr6qyU9gIzmblUTScrMnGTNlIEGD0SSlS53slnvG39
4QN58K0f1Fr6KcxoK2hPbGmKgO8MsTjDgUAO1hQ6vnG58p4bkt9stx+B+A2A0L0fxziX/kHqoxxV
6hbKUqCDnT27Wz4MV/gCxXnE1Z7SJrM3Jm/+bhmVOPb78cDPZx8vLIwdv6YPUPP/lTNz20NT1wrd
+eWgxOAq6RCr/raimIopvhVSbcT6e02UZYNIXg07nPEnk3PhbyCdIcrhwZ9Jvdq4mK1P/wOOkrNf
PIeC2L3o9+7WqP4aZtUkS9oqAbOzbREuB+1201zxf+sUzoL86yoOioBF5h3rv37BsWtw0Ufdu0Ks
Bo8JTLtD3ZZ8Qox/dLGc4bwUoSYjF071etQh/DDJ7GZMphnD2ne5Sr4HRW7uFZqyiFP/ug6Kp5Kh
e3/5Lbd61dad55C1SRZrJARaCqV4aOlfuYvVB4xlBHyd422xstno6u1bhdCuNQBu52FHxwO6IN0a
2106ywYHu3fzx1GuyjI5/Ya0YqBS93Ut4clNmPjNeGAW75JD9BjrX5y7AXz9RswIiUHdSv3ec525
8a1dKXTl98DAZXyAfNGoQd3ULV2EAofa83NM9CxoydHA8m3Ry3WOr68IPwtaWKAHkzIdenTihM/j
/qH32nD/25i1HK2qlvVL8a1rogua/UL4UL+A/Z95uBVEdEDSmv0EA13v4Rz25ruCzduSFSfR+W/3
uPNmnpm1lDmCt7NnqACA+XsjHI80vWaH8guhN42Ega/iRezkNoUupiMfEeD3CZ+BU5tB8htxPuzO
Hafagc/L9sVC/62loWVFu8vOVpyRSscNwOwfsQCz1ztdJ5mBC43fDn0y9NXegH369JcXY6x4QMsb
3Hlq1GUAcwtpwqPoq2BtTtfI1fjsAGdm5gDIfCyoUIUmCquotjUFBw+G/cRVoZBSSy0XTZqm+ZtT
hFvVsCqR0/4seLSyc8Etm7qDdDVVeO88jpBIDCFvn/OnkJOr2HO7Fz04Ur8HyxvXhKQeaPSQJ/mt
tVYQZM6Az112g0Kcspm7UoY8fSNNqebsnHkWaQ0yRt0+iKl0Ier8WKpxx5URJVbI2/LJqM0Z1gvW
IhhppcCxnkX6LAJSuER7U4RYXOWSWxLOfjwp2fi2Zo/RV397AxfIPV/R5DasTPWRNP1CK54XDlbm
fQGb6wvB0LrvNsavQlL1FJ6tcBo2Pyrs/6g1Uu2MMPIuD+x6j7kuPP7lBfqj+9SN3LXwltxqf96O
ehz68S9xPkHyuo17u0BS5h7Wquxo0s2M2G5f8Vec5H/vIapxCq2B0ARYtuMlWdpPFp0DKCu+2ShK
nLJWPLzTOzb+CFNiOpsOnm+efHcNbxeCaDx8N7qzskHvUAiyfwDc+UNYlYOksXHc431jUGCrOHfP
2ReJWWSrW08uUSq9IxU3Inw4F23b4uX3ouXK7Y7VeelFY6UnkauhR8fOzSmmG8PmzBIGma4nh8M4
S3Oscge+T2udMuK8qW7xOqFhswGx4gm9zEQYO1nEP2bDf5gvKVpIupE1O68ZHEeZb1IWLH1LMHSr
7bCgixtATHLhM8VLT9Dj+rQQeq5UjisBbi+ZqZhThIqlw/1TpK9RDV1S9XPSN3YzMeiHmieLJ1rE
w3F6uTscgXDnosoZ4yurWC9ZtXhs+tc0uulRjdcgFULhkc9yRJzNUexhWV8lMYNFUntN8GRLTqKH
k908zpCHcANqjEq/g7OGtj8Qcg/abDa139MoWZCXB89eOixZy0sgbGangSywSqjyvmeT7Oq9ZBDE
CMPg6F2g/CxyLNq2XXQGQQ/Ar9m0EmxWz6eXg4hLyRIsnbZfzgioEdmUxaX2ld5Su+/zRp7AgKRV
9rQB3+kByZwxQq0JWOlr+eKCkefNdFT85hMxBv/RK4D+N6jIt43vaZd21E4TMOjaDYS8zBQKDGr3
7xmZ6LDQGOW66S/M2x1AV+XiqSXQ3JPkD0Ml6+aFXWtEPsbYdcstdW4pYfVoaQxIAnVGA4lNPBQl
3+BEbzU41S5yAE3u7zWPM6ilJzoLHfRQQodFRUc97znxrDwQDaYu3y6J/811OuLN3eXCHDzIUf5j
ZEFi2+U1L8jALHh/8OM7vw3BCGYFX9bPKtyiQSTzYBRC9CJuhLHe/+1ArDNgGA8pLbeRkuPy9n7D
SLyV/QGTA6c5ZLnMVr/ZacyEmyNTkXnEtILwrOCDv/mmS+RWoM2WdxMXLTdT05ZUrzyftHXTT2Xo
SB6jaIgWTdtyNFnbKUx5i1TpFG4FIbZDNh0mWlH9Lrp9Sv+RqMqPkcaZLYLqyP4KorntXXS8lBfc
t5V/aCVAh0VRcLElm/t0/8jC2zRz+1tso4zq5XOtbfIFT/eyo2xWm9kPuxFNR0KrULsWZ9ISVJTT
eWeSIsivY3DMEHbPHEWuiqpR5NyuvrD/80fn+QigH/HPVxeKsDnvWi+I9bwvUSIjTEL15U4hdizM
jUwLp5rLd0ayxdWsYOREt2XWOTmFZH4Gl9ycxbM8bX+F39DfN4mC3wuK0VL9rdj9/vdKKMpCPKZc
WNGAch12/MJ92oTbZCt8UNjWF/0LAFr2JVuscg3y1V/bWG8Og9uAcsXCtX2ZBkHWyNI5p29CONsO
VA7J2WKABj7aUbBXbWuMayBzpidw+/r760GGut/ualHp0+k50YeUO0wbqe+cE5GRu4ted/nTFlew
1Vx1OCrqEaKjJ+r7WlYMNoxtIP+cHRTJNtQ8JpF2Sali7tppYdACx1lSHDV66XZWXUp9uHketmCq
fCH8woZh+fw8tbn+swozrGKAs4Ob8nfYMVLM0cb9vQCMp6wEeGC6O2vPaakZEW4AG0/2vnxT9MTr
BUWpniOwGZMpVyE5XhEgwHevmB40F5L6MnGJuhf9dzLuOvB5amnnV2Ri8w3p9s6nkNhu3j1AEctS
QH6DXryMkpKNAQOctkaTRTAqTEBaplUG6d5u0TgPertpibSxFZ6dgpwO6XD4iDwTqCuQx+ikafAl
9elTSMXXPKb3DabYEQKfReyv7TLJLKWuTccsc+4daBU3d67WsnX/wyj3DvQucZF9qn2Uo3yZwgvb
dzc/leTWVTqbMMNoV7fXDYP6YD2Yv+F9+XoSHR5O997rKnGFDHA6FdEC8bZDuvzSu768836JsYuY
p6KEOZb1UViOD5BENorNlOstDIYK5VBMwzmH/fynGVLHsRPkxxeHGzTxHT6ikh/ttPm0+yJpaY8s
9gAuoU1tuDWUhwnyGFc2PhBz+I+m8U6IZY5VfCN3rBv61eIgW4sUYOK+0yZtPmIq/OAZFDdwi3YN
VegFxwQnaHPrAvH/9+BKn5qipfqFHwpj4FzOnGagUCUFCb5ComDeSgMlx6kB+/XzqAtzamexxONv
FwGa3r4apzFzF1Enn5sXAkvcBZg/nIKnVFH47jBp/kIG79FzEZH0v61F8Q99WdRWWPMZlaY4YpuT
z8lLPKa5apa2eMfhC97OvDPww4e/BCTDbZKUbTgsK2mJDXkpzDXMsEVIqTkzI7ecoSiJw2VdYMZq
akJv7Zg3UpOX+T28PHdEzYFkU469AtADY0hlNdGQgapcUyKPxtjccvTNvCSIdylh1vU1zKvkShin
pluNe/pDcnXJFlCZDcvXxGTbAqEQQ5GfJfOi2Bjk7XCsX8JFmt3HD1YLv3EZkONQxXCHcXajPnoc
1IxPHyRnBytmbuPp+WyVbVr3cdnk3CtvCDRpmZB/6HZriNGXFrQ2x6tAc50POyIukcAuMf25QkML
FmHWkWxSItD1sibPEQJlUCofuwhMP0AV6w9g5uqDIjal2Z8mMAApJU7zk+T6aiTTgBKGkGQKVYOY
zwsPWmGtfkFDBL0odu0Jj89CQtcjdIPbidRQtgTzNEx6u1ARWCfA3XBaylm0JUNwv54WLU9URIwO
M0Undn/NLcISyMCY8PKHyxWKp2h7QSRaR3IGv/tXG6NWk50l3NvIHeQlLFN/92OC7mvu/G5e+owq
p8b9GnV4xOWAEYMiLZKkcfD0btGgjLJGgHm+M+J3pAGVZYA6Di+VCM1xWp8b0MFMyIRejeVIYlsX
ZgrA3gYrWHGXfLif0XZ25laddyGY2QeKVMdpclVX3LCE9uG2zMazrw4y3vwl00vAzRO0QgF5xP7E
G7/Cq122a142mu8gmKM81AFWRoYwmfYSaZE1CkZPsCEBLjw+vRMftXyt+kXnTFlXebUlksW//ENj
eLB4OaG4Vv6DmFqPjdUjydTIja5mz1Tx3jFHeXAHWvnUHcSh2kDak2e2pCwVOEIsPw7/pwPBHWlu
mCgHRryejG18Zb57Khn0bBWIS0qvURN6zG2mf6K1v8mZiT2/K0X1v36C9czsyqvhn0TiM++aMsvM
TkmmtXe35UjJfRrAFXYd/Kh7GNrqzYe5Kezq44O3f3g54XX+tU0jkdAb0a/J6cerfyDJhkh8rk8/
mdHMOP+MnYYxmPPBBSaBzUJ3ApGIHykXoH0+K1hxp9I1Zf5DbDlIHkkn8HZtbYPHhAOdvfziXC1f
y5cNW2dWoUdmBwmser48CyWa34YbABQVDKxi9s3WnmCKf73lplktMTqvz5cES4IWry9JuQX4cYD7
w67GQ20+gEsjnASybFQwX/6d7azgr9ef97xBSNkSR8v5Kxj/UpI3rPQC3yr8okPuDZSPn1j+HejW
T5HR8J0I6ayxU7rqmANkZ6bbMLxRb0wv6Kdp3EgI/SnrNabAvwVLLkXdAri8JcMg7eDVkPcSfZh2
fCvvWThvGto/ODNnQVkGr4YFeV4MWvvXsZmdOBXEmzbDOMAJ7sMVuZXnCLYcqK8bp3hTusxrInnK
ODXQdlUi+KNXmvHsx5kkIYL/bAUzDRhPJzCJT23pUMiZuL/qppez0fW8MvZrQnAT8j28Qd4cR1eE
Pf4SrIX3kP8czqyKW6C7gV+7lFa4SIGFqkpDPigQKA7KJqW3FR6RSVTa6N0TItPb2698ML3hvRJA
yWFvbCRcHUhywleQhLL5eaDxNwG5QRLmcY0rGYsFWMxyL/gksQ6hQFKlUiUnKIHL25d5hnanKbeJ
r30jyB1UuyUmB1j43cdFvhIbyVr8unc4jvFJ7QHTUMZSux7yLVeBYmta01Fa9ee5xcTtJSkZUbdl
UOePiUvHrGXHKxW5zKoIlZR1+dUL3nj5jIR6CE3Vb2/RMqjqgVGiwYESCGuLGLhKxub6APP3sw7v
yEPVCRwmcR0oHT81LX1x79rht50ThzHPfmpTVC7UsRYuVLwWNP2TgNd9Jmr8/VdJ+qRfutJgoz+N
9KooP5bqH3QXgsRTNBpdRlNxEY62iO+B4Plm+PXUey6pJrWrbM23s8t14sYmvRE15yi+ZrqsUnbW
VAukmV6rNx0pDakcjAmTle/sGA1D8MFOeVVWOme6RhT4R8XeXCzxNSrqjOB+fs+7Aolz3xPAoPc5
GvNWHA4HuGBzsdPZ2tori2R2NZ5FFiWznPsQfVvYVj/F2K6W+3sAJxrt/U3vjo8kYPgKDe+s3VRP
17KCHKcpFT4OHnvLZkN9lW3tYbjClhrvgpPmmlV8cRpWLHWPcNOOuQbNteU164E2L4KM1vlpEtsn
kg5u390k59DL6HGF/pqX3nhT4+X/BQXwv8C19xUkO7W3byP+RnEy2ykyda6btjNBs+EyIwn0suxl
GQ+O+lz6fMEe1vFc4a2GFo7i3JLq8/Cu8GjIzyvSKJeWXwqR9H1ktkvS07vH8gaTriN3UlPGr1a2
qWyUs4J8uUw0wV/lmm6j7/5Rrh98D0OFgHRaWoJMoyRxr2W8hwiCgn2n1PmUBnsbYcfgztNllTha
xg4TsNETCI5CMvnj0G9MCdgMwyUr53Ttsow5IJXwJJhv+N5ZmZL4EI3Cvwg704/ghjvnntDZPvzu
T1gW+IX7ZFwTbXwReHDXpRknXA4AzML6up4KyOA6dk/xKFXbzgPyGOng/y52eSfFOndDfriU2dV9
CGRXICeFiHIrdaM0iqYlFbPNpIgciVnkwQMV1DWOEH5oJmzZo+ZYzjtYgT7ChrpV0tbGYcyIaMAZ
hIfRMTd6py5WyivYN9Xf14mIINzO2EhM8qHu6AKZTD5WNwLE6bCndTmYho6ewHYachiqQAOzlXuL
i2U9H01fjpjafD0FqJvZvMzVL0vreOvyPupTwj55oZMCksIF0RaneVMQj0NiAyvY78NNWEl0bU4R
9svWGDkdG/CXCqBnIDPS7kj88gijT8lOmVe5FmjykCXjXKBglA+3glZhFm9nWNoV0FdiH0d45vau
ut9Qj5bgRA5fhPNif+2/QH9vxz7q8CmqBPoX0Ixvq/xxvlAVo8zKrucFMpqXKWdeDr6s+A84f3IO
3ohh8vyQJjeNfEJTQeHnFp+6eOpmkqGQJn6cdYechFd30lnATMQr93BK/f/KJ9qfjJRpV4Hj7gCt
1p3zSWOP2JXxgzZhDtX4DIRNLN99Hg38e4uLr3iA4bKy0PfE7TijDI9iw1aO+deKnfrSFtrKuP/K
MJk6FqbQ++7fGIHxWZ5rzJnmKsFkRgbVPMZwM16D/Pui7b+iZHBTCrun0ekwjItODyVHxZebkrvU
FZjdzSZieiFnkoAl4N0TQ0MQ4Z++qqMNiao/SskvxaYt6CSgkKkujNXRVzdemh+AAlrMzbcMU/TM
P+rRGVYHqVhzVldcXZHj2wm3e5wZAMv6A5NCedZmkIu7YnH/2KhtSXOe8H7r9gKWUKPAg4fifle/
ICYTWi3eLV4NIXianAzX25AAVo16EffSCUaf6KU5EiJy74IU5esMzTS1YNdByT17ShI126y7kewx
Z2p40P0/c7SuX2H0IpyXD7UV44hZqt7NFBhPpyP5wIOCipqlUG/pKZ5T5aieYAinliwmDM1rIchg
OoishVCcTGE9LZDCF5VtOC4+5snEl2JImH3zH8LTHjhM9+17kAuit6uNaF9/vppwFVIRibtXaspn
r8jaR2ZZqW/dsLOOOnb1CDgj9kzH4QPKXCyprVh0NW/u7lBs13D8DoaTYn3CZzrEqdqx8/opIRl+
MkXmAjaGj6oBo0Ky1DxlRxq5Hg1Gn7kdSCgD7/hj9fD9obL0LD+fP8KzdBqej+0Y0XExFzgPSOVl
DT2y804KrE7por3bYI/cU2x73czEESsTOhUkdBEsOxyQ6o0RQ371ChPV+fPU+4bLPheU9bxG5nzU
LcuyT/pTiX7DhrcQvmRR19CHsUxlQT/v0/G0Zy5q72OkEqXC6pmFVWvebFdT7BhN2244txQS9FbK
aYZuqhgJzdtfwaEgE0G5BaDM9xDWxdZiTEddwMZJTOlZKpnIVE6cxeLUObD/QqR9aBc36i1jWolX
PMSczey3h5zgyR+/9bEuebLeAqh03cjRj6NYh3EZS/KyPjuQ2G43vphEstWN+cRW+knikiHLyCuX
WN6ai92A0x58BJPyeST4IZIzraPDdxbmmd1BRORk+jYD1bv0qagmqf6Xyc73opXGDSoq9WeOXfEm
+ALEl6i//dgc4P9bF4j7lhVpdBHXEgueiVDusPZIgkdCYwiUNY+o1vi2sftSdK6RTIWfYDZGYQFq
5j/Iwmg/wlB06rrAn6Fy500Y8cJULLYtLDek73NalQQbSJSCwLWAJ+oJH7IHz5L59rHnELyHDGbb
/4T5JvjEXezHDJCkHZXbBactmHod7nawmzrXhBe3wxLQYl+NQCvaMae+1a0OLwmVrY6OlhloO4c+
Qs2ptsuaDYvznEwoIqNEAFdByHctFXZBRuY/VljbQIV1MMFFszjhMRmsLMAuFY1UtQ1cmDVh88wc
B6XugWuSvEUUAYQ0NRDbGbE2baazyAoxTqkuYjGKlwcYvmJrkLg7NrqGO6RHcGh4lU8DIt0Qo77y
Nb922+6VFBQvCacdKsYoOhen6CgFV/P1YChzYVb/TVLMOJaYjQlIbF160Au8Jayf90a1O8m7hLzH
DXINTt/AnkJjZf3Xc7nBPbMU+sJHUWzKZlmlJJfB3kdBL8KfVyDpalYBruPeC2TSWx/whT58KP5V
BWZQtK6hzHzD++Y73+BYTWizYdRwaz+Nr3+dXO5M4K9UD+F1Z7ABsH2mmtI15xdUxyaqE4w8aljx
oO76dR770qssbIpTKHRXgLnvqFl1aGTSbqoQdy6MleelyDUURSw3y35XCZPLybNRz0McYlnIzKWj
d1HFQnVgTPJsLE4OkZp0cIKVeJqqoYFM583sD6QIqQGqodYxZHExXG3fewamigR3Dcc1cTBO78l9
VM8jg3tHi0WJk3I43HB9da2vYyVrj6G3y8/WTs2h+RGJ8eRYa0ewiJ7VwZXSZF8V9QKjD2VFaT0w
u2YUfLZdWmal3+hN1RmFlzgQLwxDITvBZijcJ48MLsUTdybtOBx2JvAgLOyUeVWm65iKg0daG96K
i6MOyQ9AonaUf4kOt7EzJGuiH5SYtkQYzEvGN5vqfSA58cHJOf3LdyQ5HkWlVbFQmiEKuotZzRhv
u9y/+NBB1+0s1SOAdBLUb8D4Z6Tbrl6K0uSJY92pAi6dhs5DnVCXpY11C7xHrElWZZnfHU/TJUit
Vshv+yQYgbn+a4TGOvvi4rssBqbqvCOdnCZOExpsj2n3379gqYxnYMwKlf0bkSAksDt+tf7NxgYD
dIyqOaNQS9Jglpt2bxrJMHFsnJTEwIkwHaSAK/v0WjKKuaccykIsvNoKtKJ+Ag85zmF/Vo3D7Q2k
nbbPoIZvQO1l8tEGA3FUNJB0xvkKNfokoViFKssOqmFKPgPWf1zufGXBNuGZykoK2C4gH7d9jqvx
60Qay3gvF1oxk0lJSsr8l4q97FEcq2lHel8URGRy/7EM1cBgBeJcPdURDabbqboUDeKEBLqxZkGQ
cH/ehOaOR1o6Um8SuLSworyVXttDYsGPs73IJsMUMP0PqlYB8ofURRjvL56UWi5abmPtWr4FGn+F
u48qM5JnUsakruadzqL28S789mbKQ0J3DEAgTYhjqgckL0DQdXd74es5uPRvCiBCdeoUqTkaMt/I
n14vG4tzhPrIK5CDNBykvdCxDFbOYm/HZRTMNEVFf6Pl38yjNBW7XoWD8t2YVUA9cDAXtPegCrRb
lnXNa3b+wh2bIfQyH0YB/mYsf3t++7Yk51fNJ27x+T3N8GC1bto9KFyzbJDZf+2effqWSGT3jpln
tOu95YuU9rSZycX1/CEOjHK4u9qcP+rgLqcha5FfrTncW0363+ghhFndVhj5ZH3sJFBBMQ8RS7KX
JuuUROat83z01Pl4TfwHUB/sSXGWFrAP4fwODYYcRUd9SpdzLuxdFUOcEy3EPApzyKIfKzNM50f9
2eDCaaEKN6yTG4SSAgyyRzwoqn5cBX75gWg5r6yauuaDe8ZrlRV3aBn1FW4WbFeVnhRk/QIfLH0y
zMuH5XVfoQmuc+YLTjJDiD5JICtxxMkOrJ37EeMHQvwQWrNejZ8tMZfHE3DAIx8skAKQU+GMQR75
wwxkGXWpZorqDwM1m/JBBeh4PQNPo6yPlGPspvM8J1pdL4MF6LML9/LlhO3V54saVeVvSs4M3nBs
V1YzTso+CVCJ9xjXoTObuUPUc+KyjqQIKCECe9332EHHitS6XxvNp6sm9v5FjyPmZgwaTgDEmMld
P4MKIQlNIxXxscXA8/bmkzohgQBOMYxwJIE/ELFT2+qD+bYFv9NJrFXdH5zDYY5WS3SHKbFC/ckh
gs4BUXiXHaVasXKKvLhxykK+OB+ICdUANp6OKyo5Xn9WAiliBB9V55CYJv1YfP4No4q6YpxPxaVY
rS6Ud/BbCIqp4rIrAiGhcxc3/DXkEB2YzZiTbmq+npR1HdFdtq38TcX+bL1z2nPao5eb+Rx5LPym
Py6Hz5GLXBLBCtQaVFT5a4mgcbqVXWGV/cRMYjAI3lAUcFj/84t8gko/eG3qDFL55rHF3D3dzEjH
M7u3fSe7R0MuRPC6Bep6F1m+ozy1e+3H631J+VqTk2v0BPrCrUTqVi16CwNWTm5tuwRCH9nE8tew
grHOhKHKG7ZVeVJymRF5HUXwLdzSH3Kmk3L/Rab2RxLIaBo7XoB5Mcl6lsbHIV0TtTrOgtSyqx88
z54VmFcbjJRhYLF6sYH4lcCsRi3f8RAC+BAZJnUCB7B1lQro4pHlskR49QJeJrSb+9H0kdCZP8+g
tNBLdOHE1azp3Ea4cHiwFbfAlz9kWWyPYZcug9jSTLH9FBVyQav6pvPwOkDUvjLKurBuP+j8pc6c
jUy4pbuhH3n7T2qWMi97KgyqsPZ+m5rAEQ4N5wM5u5dM6PHMYXblQ4VBd9+eNNRViohbeRgku8sT
v6jpD/UAGpELcBzFt5ItVB11n0ePht2671WCZUaZsaCk1s+MDXsk4rzNKgE+/MovKBjtQSab7CIQ
tZDmyi/Isx7gAz8ZZMjqN2kmj3GRtPH8cp4WnwOCgfVAOtFHUTFX45Qoz6QhtueK7iQUVzPtP1jG
6Dr+su+bA2h4qY4pC87SQ6mXa/cldb/c7U4yPCHDRXZLY6+/vZpq5y2PeaokLpuGWOSDKOZR/3rx
G97jozjfHNpwcDP5O9Rbj2QWNaK0XWTjxRzkZylA/KVrxI/HNdW7mLK8Edv27UoNAYRkmgwGNKC9
Q+/Zz14Ytn7esb0gryTxv4ln38Et34dZ2g1fnUE6xE4n57/4DH0kMTdpTIoyB+QqZan9wnfe/37m
AXKCSMO/CUaW5l49fwikcrLnSwTFunZ3z28bQrKat5Cf/P8MbocUiHD9kc8I64eu3ttzk0gjg4Ct
LyBl2+e8if7PK6xyryAbewq1np68MvaonEaUBUzxxP48iSdbKGbtDoJxcfHiyeRDhSyBh4mOFF2D
8bRncIk/Qq+lCtaz/OiAkuA1JeGNh73SV2AOI3SmVKRqIlmZQe6bSK53ePSJSYaOfX1nplMWv8fm
AIVyspEP/xM4Y6hgTz83/l7z5XXfvXEb8M+xqEZyoDlZgAxpy3IeHFQnLerewar/9ZI4SvQegdo0
DsjQI3DKkO2LJFy5xks5s03uinSWIGZ1l+col/wv+l5vQcH9p7XyDSVjNw3faI+PJI0Mz+D9nc+v
A6rs73sdJFtz/r8vpTXYSFobRtGyUBZ/o2hgTult57WClqGEVDP5o1KLQKR4Hn7S/Ftc1N1jKaY9
Zk3g0n+PauKqoA75Js1HsZoINUs12L48GPnfYk9URrMdkSyvhq6KZMweqnF+xP1OuCtlgYDnGyWs
dEqhz8HjaakBPUcZZXRdJm472DnTOgB124E5v4k8MI4Lddskum+Odne63QLoiRTdwE5dV4cTs13d
/ntLD6jrjfYH0wikSmv57NzQBplAxW+RbrlWdfZWlCn4dptpArzLm1ME14AtVS7Mf0INI832vUxc
LoAuxDx0gW6EMuLlSf/6wqY01sXRu2xWfmcsn8fQWjeIRbSL5IzXZ0anNoVSIUwnYcKgOtB/xoqO
ZQkMMyZVA4NH+vo6HlBaeqfKP3WHq4KMD0cH2MdkSaz5oJQadXQD8uLi/pr78CdK6VDuEMValdjH
LbsunhKCqfasQiQ/iC6pAVGl8JBMFdVdYWpo4pFfdgvEh25hlKvSJ5Wo/5z5kiB4vualXr74vr94
Y/qbh6jbjWbpCkt0kFyB/5p+4lrBlI5PUce+Rxxjuhslky9USWWM6dbXaS4PcJCJ60uUvXAfTNAV
2fIbL2Yv4mjEjKR77CXI7fsByhTcyLKwlGH5UDIziT6vHKxPdH/ejrbrfG4f5foz+LiRdCFmNA7L
Jm4HbBvAyb8Jk1+jnz7MVGndmb0Ky8r6wEYNmka4aEBOOXAwcNTq1Ao7ljxpvko+rpzqJgcbm0rv
4L22zkN+8Je3ZMLWLgj3+e3uhWkkmjtqb+sMvjMq7zTPCm1425GIMvP/czpIzZl/kPDOkceMKT4O
3uh+GxzKOq6CID+QtTVjMnBxkYAYzpocF8sFsHMqXQpUqNnzm75CrD9aR8zlWtAAd66LfiSpK4JK
Lgbn++bo6kYiVWeYMG8WD/dDsF4ac5KDAfhIioHqPvwZM6dG6Kxs+dd8AHXOvQPdQktTh+ownlJc
gsJDlLFokKTixdCtBODXCDajifl748vH5xMAGW8/uOsTiwHkZF79r3pNQWKJMQkA+lou7Vx6X1w/
Jsj9cxRysO0MNBsuJRO7Hamu6RmoR8v/qMSngsJqf/5PtRSVo3j0V+84c1NKbaWj73QBdS1++vhj
Td9A9zrBPdKjttdlU3tFSg1xzoCT0iotxUZvS6awxcGC9JtmxLe3aQ/0VHB4qlCnB5LqgvRKBBul
7/fBZrBwHqyB5aVKL8qqa3+1JtdkHb8//x0EwKTbRh3edfEHpw1jGSvDJZU8jA01v5M5DxjuglYQ
5D8D/pgW9W0lpDJXOFgzuUH2U6k/kgwYRmCx4o+MLMKy+4Idya8KVc6qwYSOpHEyDTP3mXcQN6Kn
aQs+NsJNTMtUhxe0LXUrWi5YYK4enJnESBu3DSE/SHsh8uykSCj1E1h5d0ywfaW7KmOGtZwHhilB
EKjEBJ8qBp978sCw3YryCcfIB+BMVVGKWdZQ+7bq932D8SYQzpxiqhlL9hK5iP8+s5T2QrqO33vs
r54UcQ+ke4Hp6k+FH2iag3s8rxhfNyarCQj0i8swBozmKn4Qlg+jc1rI+8LxI9CXU6mseGlB3gbT
AUhovUrKyjd2Mdao/o9xqR1jWjepH3mc+DrNkK4mCWhzM7t40Si3WlXeDYaQJJlXH9HoaMzSyxSL
4xjFitn/Rr0zONeJRxdYRk63qr+t9rWXFH8xCGCVhmi7CDZv5NAMFaIJL6MrRMQAX1MKMj4OiBkc
iBAzbiOF6yKhzFm/VEJAqaII1JlJ65VI+0+zvHqz8UnIGKr/OKcPc17qePZ6vX2vOQL2ILrpDQ1I
mceAfhiRfhJsOlzNJI1WU2pDg2it+bYR/fa1sylXAcmoHY+kPuyqyRPUMy8xi4sT2Kz2haencEtu
fw+itzOcRwUV8xDs9d1KVbx+rusvD3ffna+yfc4l/6zJ0ebWsijhxEWc7zTSne1UqN9sD7rL0yRP
Jw115CgBFTVhTAZQuYiJ/5n/3lFtMKUJRnBXT/VkhWcPBVnuPA4mPoA6LFwh4HS9kSUr/ADnT2fG
O0gQyGBqjuK8kGvXeHquvufij1QmRGj9yaxUvho6SQfWwUinwegKW5cGA2U/hLhkU8rmaGBUne/4
loWNVcbGZRVBJGAYLXVGLAInRrA2WVn7lNOUkSQHmUsEMuOVEhFUWR4vCWJHPWN0/Q/koWRNT2BX
2ZLh9TQVNTFeI0FkwlhJQv6bXMnb2i/dY4luShH+u1VIZ0CZ1w7cntf6wJIkQZ6ehfFrk8GU6gYw
S5w7oeXouamvXcPtp3x49HonZmh8cy10sc6Utk0DpYiAWWmd0/rAkj8b+DdHqx9XxAajqWjJmgwT
EVmuatDpo7TL2ita1wOWwMaDX9ID8za+2jrPybt6AYCRvAA4q1vxzhQWlJLtwBNm1hyDNChE49Z3
avW0pG51ISZ0rPFBdVogoXjYjKCesOxCDRqEynhRU/28wiU09UV9HcSTu8HMCyh+UcthrFp0Ef+/
2j762GThZ+OrD5bj9+GjQqU0uP7ULQlWNoQV0STMF2eqkxXvf0SzFzrDJlJpHuKCRX7oQ7OBhYsN
GMMVZxyo2rtlP4odoLjGaDqdOCKbu4L++dg6rv8tbc6ZsWvPuZgLe7C4f4f2vohI6yT2CzSDSsh7
tJbID/ZeA8qdp1+0gpHF9TFFv0CMEV8IyzsUhi7UzLJLw+myCsLXk8hukC9DY/QiIsmbxJ08CY/1
GPKKhOZOZyE8ErOnpuwfEyyqDmdz4KdNW0RP2+6LGIlgQFh3HL5XJ99pA/HAh2kg1ZDaocGUjtv5
WVKH2k7Ueqeb2pjy2ebW+FDNdlsKnkOdF7EK0e2ODQrAA7E4Pz9ZL6Bp0tX6TTGFbUbfZoRAGANA
NFZCuAHj4WUEjrhEmbUxP4C4T+22vndl7Rqh2weTM4QJbhP2vnstGmrxB35lFmnGO3bIxggX4+qv
pPos22sGRNRHz/mbPXKc4qw0Z5ATwSf1bY7AxFnxyWSNCfY/0UWLIiMqtD9eJTUVh7eA3roThg78
J/t00JBq6BIbGCnk4OgM3N5m7niGAM8v1AedongENZfqJLVi4d4YkHiYWDL/DZKC5W6Pbo7k9pa6
gxx2hT6tvV6nz+3yRe7tM1OcY08kyQ3BgUAQYlKLuSUClH7mtpMPb5b9RSsvKrPlcmqQBI2+EAPq
VGiGYp2W06uZoHxogsfoAa/4eRUVPPOWyKb2tyfnwtw5wxAVQSlAOnCxA6ifXadg7ZR+9JWYyoAy
MCMDMugBKMjVwnRhnU8PtoT/RJNKct8ocCEXehcTleKHPbCwnvkPlV/Lz5Td0iD1S9NTr5Ucvi0A
z8klNgDfr/xYGWWfLZXysq4b/Qq1aArN6ou33xVtQhv5Yk6ofhOoooP/m5iQsnG26PraoOlM6pal
dDQWUrFEpX4WKDZqHYIhZR5wlxmhUGeRF5P2TeWa5njfVc7GLk2DsigMNIRLnQ/FSgXiHiCKe5p6
46R5gpEqaHPxlVrPGzZMTGx2dhr1bsTNDhSu0Tt54hPUhBRfe6J5rfPHyTi6jEwOvLE50XEqm0Xs
BsYW1PP+PZIA3P3pcq4NGBXd2X+pzxEkb5qroVgJgJux6ewJuM4qTO5uK1l2MytWVdaYR47GYYrL
VUBuj3xZwPWVhEE9iTFxw13GldcOnWd5IK2m+5t927PWnvhZuzsFlkjqJZznXCnWU675S2GrswxZ
+InYl2eIX0/52uS8RJifXvQ/3cypem2D8ml27gXrRLf6jKMEmyWjPXFpdw7wRs2EbqKjTc8/ey5o
aFbqqOu+j9eXvXUBDV9slwrRpxCf4LIiJEnNyY7R8loBvDO0Ie6WnHaFnA7ZCmuWmD23xxYqLzfY
eechOVHonx089aU41vawtxQCr3iVZ8AvNohvjUME0h/kWiT00+0kKXh3DOhwof0XAQ5rkHFYF6Jq
FXvFQFMEHJPg4QsycCbUSqVtMab5AFyqLkNThakmM/H94johAEhekMWO4HDwNYhZcMsr6qhiYZTT
qn0SERK7cf8t4THp1rqMnR9dj+Oh6gm+7mIeCp9qSWr0L1o2JKqIAe+EUD//LLGPHva66otyGQnT
/rPvrz3mYXVVCJeha2eNF94zP+4rasZhSjoJXM6Im+aYLJOS7tzo6P3SnBN4vOK0US+R5ry/pCU9
bCKZXP/kRSGcHOuKI1be+3/KmbV2E3goZgjqEU5sPuuawmOQ/l2U+s0XiciJDdW8Nff7kNDlDOVP
x5IyywmJQD6tu7Y7U1WkAsu3Q0U++srAfMBcUWWdfNetQJs986i4wE8vGSF46Jxh9+hDaYomXnD+
DXlYc6tDBUokQvDpPqublk8CIyLIwrW40xuEUKcwfS1d9CzlAAfO5mtCePsNmr+HlzJaHH/f4ZpW
je48GEgS5KOFP5x5BwKcwL48zB0OeL8nJ+qLyD5yP6agMyns0r/sZIRua8MyIHzOt73Nz3OUE+or
TxdAmnghJDo0rUN9bdwyfrMoaTk8FN0WCcjDusuOfXM4JV6Nhme0a8rd/W/jEi8XEGnjBsFtv2t/
m8073KkDtg+hOWD4Hfn8bWe2x+bp8FbYTzrqe9W/ScWso/cDgfShd8nLAdeXH3Vcto2lljxs+xu3
swP3UwnZeRWXDxiNqPVyjoDuAtRc++D+Xd9Yz9DNBIl71H4RS9UrrcLM8qBAHEaRe5+Ui+wV8EBY
HQMGGhCS3564ZuQXRjuApCPkdIv8m/NBowrCNpOzjOvUNEJ4TeG/zR+9p5J0q0t15v2X1E5bBkpu
EGoYSVV0G2AjdvqOLxs83FwJoEVdSPFEAIjVxZs/ZqCPKnSDTeVv7/rvk7PgnfNMwEONtOuDxDsH
XE0uQ69ABlmAkRsSqpUebGjpsFeyDUqHTmc0VXkMFUKoFwR5u5/ERP3aY7rpAVJ47lqAU2oPO2k2
m9RNo5jvVkZMJRVlKtcGHIqrMrez9TCaqcfLo8g6KzItmEhOA94z33ashyKfe2dHVnKZ0ceGiBsJ
HC1blI9MJZ8HtVCgK06dFkFg1OR1meE40AWqFxFATq5bU6Rbq0jmRHI01Ks3MHLiGxwV5RSKSzPR
XCwWtGUjDphxWrHn0+ZF4W/erjn5rzHdOavCuMQWbpuP7zngzFDSiL4aMVPi58T3P+e8ACBZ+XLL
DEPbabjsXg6yEqyKO8wpzZF3Uru+Z3WjUbACVRr43q/oTEcgs5FbpawwVSvfL43JntPnWC/LU/ZY
znAzejqZIVJyiVy04mmBkqH5i5+hSmJfCbT9FmqZ0VMNFxnXGjqFvsk37Ax+cZ30zm4NtvcCT4U9
ZKFDyLqpV01aNV/0NsuNRxpHCoM5FkYdT/gYsKMlrPdA1HJ0m3mqcgQJl8AnqQMsDEHYX5bVROkG
HpLW1aJYQphQhRzfeL06Vb28BRkJRIcQx3/tuQoVmlvKK6A5fg4g0VLL45jdllnFurEFZeqaAvuc
W4Uc+GPQxIa9bI5ebz1Mp4lipd/meQC+b1Z1c0TyRvpywqFlNK64/DdFfwENnBw5g01q3XLBu3/u
G959Dlq6ocAIVdwJ4oGHhDkCs0HJL+s1uvZptEFCk7Rk4Y/YWE3OOfJS4TruOFXh6cn8ImYCerNC
k5QzS8EHjplVSoQuUf5fo7lZxvcHfc6YwR9WIxZh3BA0Vmsk3CCLwGyQlF0cWL+wgFyePB3XU90d
MZrLFBxb/EA/LR5aKVPy3wZOxFahaAqVpirbFMs3JPPQXZ2mZXe8yRAJBWETWxpXyH2u4wMT9HtF
whkn2pko7z2g0iMShLh40Qz98Mu0gV3Gogpwu8T2xrq401ESs8fNkoUZzdRWM9sNZiONbQ4iFRs1
SI6ZgxVrFvKYbfIgF3B1JjgdMXi1U+5w9Bqm6stcaLJd+drwIVRRLokBMVIFkGRxdRE34utR+gw8
Rxi+87LXv4R/LHOyh6IQ2dv6Lyhf0V2VyPI7bETUJGlV7CDR/tziA9crrY5KW5GCr1C3o2GA3QD7
1gGostP0Ij4M0tiy5qvnToWxDJyQ/4/JCwmSrDv2WIiXHVEtw6A860gBv0+jmoCouXqavkAcsWDd
C1DMVaILGBpdfIWLUujOyzqhTVczHBJmeCUAaa9P271FWFdn8TqMPZw7rgYyAwtbiTlXY2lOrZ0q
uR1oq1i7ClIQtWRZDIBPfKrw65oajIU3qdgffrQZ1Of/7hzfe1oyMxgeu8xR6ICBDsGGIHHyYqAN
gUS9LpVWtUX8YjCdczc6cj1624YNkz2F8zuAdj5QtZgSWYspv9U1/KU+ARm3VKdzlmSyuV1N7/0B
9DBJbuXO4nFBNkwXxyc3DZzL/gpVkcJZD3IScrj8WjjQ2FTIX8u3lo5sF9UvwwU1qS2nay59DUGr
y4rDn5O4ZZSJXR2GFzU6GqWUjCkHBzhCUC8VOuCFnMU8DHfJ94DoMSIBDuZYF0QPeiPhJ0urDxJ8
vIxP62kQSqDUJ05o7jAYNI6fZLeDDcVPY6/qp/+LQ1FDwTbXIwXk+U9xAVt9a7ODOx0mPCfMiGG/
3lJivrwaAC7pKGDDgMseASvMRtEUgs3FBBih/pL1z1rQI/5nsrThqURetsrgjVWZ/hYbvNvy9uXR
6+gpxJbtslUyK6uMlv519ei99TJ3sOxxNSCJc7/6LK+LaI95CYD1Q6mQROH3zBgASx3df9dTPzwl
gb5P81iw+TjH7/HkTEO1bbYIM/C77S06AzVT4lra7/bm1gm79bHH9+udMJ1Yw52it5XpuZeXMyPT
MnYY37rhZoUfeCpjnw7aJ3D1CiH8qK/RNm+nhO+XpuRjCsZ/K7dj11L7YeFxpbCI2Y198/GNp53R
QTwRr4Zd6Re6e/k7hRFsZu30QFfmg2w/Pbbl0ipGS7g5wRlWHP2rwCOuMj/G5iF3T4h0uDwg27yv
ubI4Hkow+0wphoBF8gMbd9dhdYkWkG9VelOnLtZm+ZxmWgjI2jOVp9N80hWnEGncuzOtbZJcoQHG
CoLxtCJ1TnurywxmNv976mSWVbCXqk6+DeoVdvaxsMyR2/7ZyXIAkbKM+VCBeBg6z8c/8wmiH9/C
MvNrdWBOVC/dRZi4K92EEqGTuomPchPHe15BvDVIwlkrDgQrVL9iPCOoJZxFi2MAMx6KdcG/Gobg
OBB0Vs0RsLMDWb9yRt4mRPoHvn9/DzK6ZxuMF5N0+bVLbuir4BPL9tsiOi/sLzMPKVq0UYa2Hwtj
7RvQLZfXDiLchTtuv9ZAALVyZNhTXQxrxcL/qkORn7T5Sm69+DjnMInPphoXxhXBC3VgTaJ/DpIm
gEOdOib/n7fOi40b3AbcjwSO4INVyIE1JhoDn1zgeVrBUZR3Fu05LA1Ee/QoFQDOWP0N7Gaw68xQ
UMrdie0XN6VJCuUyYf725qhTlUWSS4zO77ZslBvktav8eBCcRpFxE+YjyqzdVocyYIh9M5CRYfK0
0NT6qFUQ0AbJrfvvOw3XlDGSf3Hw6H08C2ZhV4vGCKUnu/cvmsRXBMxpFDsDT1LbJgXPPDOTNFeS
Iik4G87Kr5lieC2JIvDxaQcClpHN0rjyeZKizBr6bUj7dWQWRjSNWfYeUg/Au6tKqYGkti43rD5M
IRKlcwbvEmNXg2zMP97OA5c7KoU/qZsKzGFDiQiq1vu64nYB0OialODAIfZWlyHNw1kVYgvRF5IC
JVnISg04vKb1iCdmTtvUEMdFdlDDVZSSeoxgZ6LkdIsZP5DLEoumNPSg6gLcg+YWOmkpdSiG95Fw
NeehhjC/14RT01QIWEz7WQyVl3NiWvMJ4KQDg7DPgc495mV0Z4tXzP01UI00Ejt6woOkfXAhKasa
+6NHm1e0eQU1JveMt6IQXZbZ7UWZDb+R9vnM2eCAmqvVrDUu+RcvDmb/n0i4hMusBD0SMqkMF6aP
IK8z0RsicDHe+P5sujfxGRwjDPfVWPIeYOq0ODvJIm2LtTrN2APEfso/9DF5UZ+iZJXhvEHpviO1
CrLHfCsssIGQNtu32hUE7G642dyYsT+GJ3lHPbdeIjelp+z6AnVG2oXuSs5LnCjvc33aKN5N+qUN
Vq+4iKpLubed4ZJvqJTlXsuViSwYgWVvjHqvM61KhmCZc02A1qRs+NxORZWPCtXZ2HX9h0ABcaYb
0axoWNVfb8XHn6kdecpHSW14PzUpox3+HTuo9cAOgrp5u3Qj/aM7y6gRODXiSD/Ua3rJmglaiXSF
j4yVHd6VePrlc0rsfNMVXuMrKkEm7lasW3W04pQ2Ou1gs3koAhB3eIBUN0Okiv2fw6oVtJnMA4nn
3oldm6YtDS5K5NQwyMxvmS12nmr6GglUW8HYEUmFZo9IImyVzEjAFt08qZYIMEXiF/TGZB+ALsg1
0QU60e0o+LdJeknuEURd53VL5G2iT1duYlTpqDMuiB5xaNwdpYwkscL0Y40KQ2RGWtHVux8pn/OA
aD8YZWRN/81unan83LAJJHa5kmO7MUJ5LdjEd4wEG2zfYztOuBk2LkgHGD8kgAlUCRYh+0NjXtZC
yqa0BtItAT1TQ0KkhvNwkBBYDterln69Un4JlPNg/Zo+roXOwLfgkS9CSpLQrb1yE3yUH+jivr9q
T0088mt9N9wKIyT7gCaDjLtVQuJAK61D9QUDN734i/ksnb63iGzkYbHlw4Pr9rhylyThg8WmwwRS
8kyL9iogL2P3AO+NWs+aQuKNyiFPkDure+Uoxdmb7CnB5swnOQ8j8G6DrzdWP2mKNCEYeI/9csct
6PLxatatFcb0fFcVCX1Yjit61FykgEpGL8vYU16MY+9MbTu8S4NjRzutoTGUuYCkQNYk2+XBl1AS
B9u+JCv7TJCc0r4CpkMWyJczvg08ArusGemJozB1BtyataqF9aBfDMIfIzUs3jvW9G+Ruy5K7VgG
Cn0A9LrKb22Jg1JvMD0F18nYFByTJyD9Y4cnycDLKoo6VXpi5eRhkYwLZXBVFrmsDkQsE2mtEhWi
bCTpCY2dAVFyyvqLVrMTlfWK2oruJWXGGhIJQ9ehvEcdySnWqNsUgIXkVZO/DReeFENJrsh6krOn
KOt05E2N/385ZzlYpGuPhlYHL/sIwnxqoJRX1k5bcJtq9UvVKPBU1IEuSDXNDYArJ9mPPe4nu0EB
aeyJKV/QmwuRnyMICztSX86/Qh2sfY1NBpf5ZcpnTJ4feQ61nE2dmbP4cSYBWjHalc+/G1BBSHwx
Wx6Ibrh/MK2Up5ZvvFLdFALZrnGLWlT5LZeKgkYS1Upi5Q6uy/Auxb0TFF/whrR6w3MfzTpMrKY0
hJr49BCPzt4pcYDnlCieGQdYIHVEWrpQEUSAfQ3ZQCZpX5hj0v3FYtj4VlwtWEr/wnnsHblNMO/Q
9eley7Rth8Dur7+bOVajAHppdvFD4zciyEg7xI8HjbiP/eJE54VNecyseykh3/k0T3pDRfm3VKE1
crYeziTD9s2bqlybMgtNVhjg924Z102I9/ZAzsuY8DeI7Cbt+KZ91xBUSivCAgxil412fbhr2Ifa
EMQonW7ivixuQLvhYh/cK33Rm6RVTM5+GUGNZJnvJPPvNhQXu2nhlmesuuMAcfIfzDTvZvAKSjox
SBIGVHzEdfgb+7bMGGucVfHUlW4IdD5vATV2BSzx/mLKYrqdsi4XZkz7SykTfatvE3KW45IgKOIr
y3+e7ZBbrmAZgMgfveD/v8RFV2EUKvkwi83bIt+gq8GViRNOZhgqhkHGjd5fc1x5NDRrifIv9D2U
jirdGY5ZpPyn7DlQXc+v/bXOM67jzVbuSC4D71e/YrQ4oSPMu1AxhDi+nbfb1aJxFRDyb+X4dowk
COiv2iMemKL2+bI3IJW+DRuViDVe0oenXL8y1OJtxkv4FxIHKWYKoJmRQwByWfO+WWH22xL5CAin
2Ob7R/TFkCivylRYi5tmwn7AzsOZaemRd3IW05ud6CVNM9sZfmZ1Lc4om/btxYIWTI8AQdoEYjaP
0nz1OCG++b2iI/PDT6zLj+L/z/UVFovNNGFUaSoJtHGGpu+hKCXeu0gy7KZE3x9C7tUbhYcfNmVq
hyQVkkPTziOU/d7VtdKlQld/HksWWP0yUqFIxDLlZVNtLBoKaL6gkZhkjBpUlLkgClUHUdjIdPy8
oLub4O0UwOdBkXwKnUNPrjWNIjkpFsAzeu5+Pmk3uq/Ukz5C1yLExlLw9Wroe5vyCODOrRXItGyB
Bhh1zB60T81kxdNh04Nzwlxn82889nKEWqUgfvcjsDPQCY2ye/sfbWZke3u/Eb55BdUArzgGFipq
c6gBxdtR7++W2vKeHqGjEbgUDT5g9rzR1ydC7QWEpuYLcW6ls+9TC5haC9uouEMu55GXVuKIdFdK
ZR5mOhh8p+C5JTEaZNa0X25ketfK+ADh/2WIllSlnqcHO89YcsCYXX663RMXmTfxeSVOSLEYeWxf
IVYp/jGf5T4tGP11Vew15ghU9bekBuQqAD81JDTP1Cpo5Q2K9vYwipqRMsFUjhLlcR85id4lB23n
YbAJ4MsVg+anfpKmsyXQBfkbFjk2xD0orFpnreBD1Vsa/v+frnpyTqMgztulffhRO0oFsJPH/8KL
0qdhjj5D1BirwnuOZ0f2lWtEkSIY/SiFi1BuhgBKgUPuifcdInEXJ0kHZzEgKEAQJ6NRxBEZcuvT
r8zUuZAqpA5BumlP+pVdmIQFL0aCRcS/uQ2QpevV5OY5KbZWrmkWTGabpNA5KEWOT6A8pAma3B6U
1MmQQzC3Ai1ef0HAXHUbrvdqTXQFf9wkRNcS0l1dtzgE3KsAotMkU3IwtGyC9Bk406+IFQAR8N27
mvdc2GtkTP8VvjLbRhKKd1+YoUt7dhdL/8QLV4GdboXEg8u5yrFkV5HicAiqQjrsydg34+Y+D22o
7cJGPqEXaIR5B4BKFsrjoR7cqJpy+Gc9MVYHEo678FPXQIhDxkj5yHMPYNCYJT5Kl71AN67k/rRj
30R5fRUkQX1t4T1jRfRxLOWyG6av850YyhafbD++UUmYnprfFEfQv3Bx5ldEel++TMikmwVxGeNp
4/IJj4niTg5n34tm0RRZY94ldOnTDbMD6rglUQqNpiYs0WvkOUOSS8EkQzg8EItK0IgdvSK0QX+8
Po1LPOJlAVrUSlkzXYCwVJFzMm3n/qJkqI9Jnk37PzJGtFKdDc2X3VuhGmlvqUPn/RAVXBfFJGa/
bO7oSwmPbvJBT53HkwRiwgMiyW5m+gfhLRAfge+W9akG35Kg0y5u8O0esTc+COCn1M68b9O6jH9l
V6EYLAYMuBcEfkZ4cPweBeOtOZnRSy/D90jsJ6GBF3i0Lj8ps04lrLi4QkTFkrQZQBgGu0qP8lfJ
xR6oHzIVd1UGcNtn3CDcLUmUIg1Qp7KPg98yi+9dmNG5auyr4GUXBSMpHbEcNoSetvbTzMrU9ZJ/
houi+b8g9YmrK+yCuTxaiebBrxgn4TWhyEqj6yKsUmp2DE1wAnYKdyfLmNndsANmZ2CgOqU7Khyu
Mye5Z6R49/qjNIQ+ROgdoJjD5a9jwRCOBuKqaEPyGkM0WQWfznEhCfjzx9CEiz9qhhjTnjYeKQjp
OczaKNI88kqcVwy9mT/H1P99b7ZvaMUiEAT5RWiJWvm17m5D6G8de+9gNiwddUuF0fz8/0Xf1wD4
C3HW5EJ7IXoo1yg+8/e4iyarG0boHzSlNd8sn4xaaWHT+ovwceg+D1nyYm6tMbsWt3C+jxiizzcs
ab3kDk2F73fcly3DweWYQ2dVKyq5Ho8X9jIBXSCIPV11b3PETmWAl2y8ZyMD+ppSrwu471Neb6Ta
JVzx0FA7MZi1kvsDckYfHyoF7ER0TBV9cUO9HCPvcmQT+B7R2BtGNITl+joA5UE6P6yczqKfSWgS
tM9OUui0B50c/jUwW/BYdn6K6RMvDtaDlrG/Tq3gO2rfaU7pJUPphiaPx8z5owgwhoruA8ci5oUn
su9jcydXSfwaHAPpNos0U9JBc4TtpoumCW2ivuoa0Z+rm/LZGRJ9nPmu9CEl/GC5PPR/U3vuWevY
ylCteqXNVgncszLoMweaEd+Va/l5vMBCHSzzZJe7DQqQRutd01myVsGVQlHufOM3dem1m+3/+yuh
dElmoBo05v7PZN3Z7r3r0xXjK7avK6TWSYw+Bg6z1NWM3FvzNVyK6mhypXVyUdi+sA/9fwfO03FE
yi1P8K2HHdWjcxum1BiRmBuETLNK3nfvMJ00raEqzHZvrHJrzyXjwrotjmmF9tcIOvt5xnglfA1G
reT4M0RHCUu7Z3hX4xofpDrHnu04iMRqRcp+oPGq14Th88MvS4Rg9FJHGK5fRiwNNPTjodqzWjhD
pU9m6+V9/xvJ8e6NvvS+opQ71R5NwNV4VtXlyvEsJ4cOJce+9CYH9IQjzooFUyEgCxYrkMeQRvzY
uYPk/L7pIJAz+ippotu9se9TWrbFFFcyHEnZrOm9zAFls6NcM1+v6XcO3d7A0YrZUZ9Os9+ayt4g
bao9gglZzyBqlBBabWUqF8UfFSZPosDNyJWGSwKRdH2tfb8qloIQF6N8Q/Dzo1odebFlJx7OE97U
lyKaHa15E89191OSuwYAi4gzKHkPJ0g7aLeMvgJZ0zS9xJWVFkvvv8O5D2ZVuzQP7eR/faWYa9Nn
Jb8a37nRKDievWTBsVala8YhhhGh+7FT0lepzauq0lxEPuJpPjWokpcmXIxWLCiIaeeklCCkyHLI
kr5HRaRcBHj/hPfySeif5lMCMl/fjoh3NrWZ/6gQ7PSGWTqUmWp3V5JP6yqirXpbY06LV4ksmWZ+
omeqL0DIk65MG6s8VEez0/Ez2cOzgQc0qgC5n6xa8C2AHRNha15CE44mDbkcu/SgRl5SPpUFcg5o
aZ9u/1pp7k6pfx2xCtALX40EFvZBWTIFVQM/3wNBgqsr2V3XfexaQdqILFjYex9ks5diFz0ANiRC
Ma6qvTiQjgu4niVZA5f8RQ45eYLvuviV8iXz0BZHFAt4J6l1++c7PDYKmObAjiUrqE3PHeR0oeej
SdJKWuJlV0MDimC84WxIV+J8TWTzpaGl15dObXb0QLuDIdxVbdyWZT2PkbjksQerXyxsMkv2t/2I
l4iKJ35h1jzuvD2NrohqvC0csYXmbJLgCCyus3u9SZk77LD18HFfOw1CWw13CWStAUH4Bm5PNCVk
sXM4+nz875mWnf1luX8ruVupnh9PQe5r5xLz6lrmI6ZhUHTInA51oY4KJAUHQW77oSHmPw8+rOjZ
Q0xde3tYfc7RsbY93Q1ZcBT+f6lHQubHJYSu1Z4PBbfa6ZBNVJmwY4LaSUl+YracRRynzPVNBZcj
P3+6maUTOdN48Z+HTnvqATE4zfc53Q8Y7Uys0L8jyiNNPmpG6htgMwQMXRbfhY0VG27ji/K1lZdS
G4OtbH8ZnnB1NoK+xqL0VUFDfN7gFgE9nBBRtoq4bscEXifNzVq+Iu+5GqlwAWF6f4Ad0/ovA11F
Ij4dgkKvJrza64w+gim42qmopgTSM+XXjwG8eYtVH10X9XK3KtNToGynN3n6q6JqDyLGLFw9Hc9A
KtC60vf1shAtTLIjd0FCurON1strR4Dkt3O8IR7gjd+5GJTnwYvsT/vm9yLMsioin8WR91CenvWa
c+JGQTL2O+yjYVg+Wah/qCnF8bb9tdYoh8XJM2l7quy8LmmKAdV7mgcMFnB7u8KubKs7TI2nTg0J
b7i+LCTZPZzHOf/bIMYRqwVeOWf3Uh/beRIWPvnmmH+XBYGGGAeZRtCpf7wemXo43UphXFdu3JtM
ANs0iANswv96TDZGjMOBny6a/w3VPh9VM361OBT2BuAMrIzgwzdB7CzC6BW3lvAa8AxD2St8d/nC
LXBnWo3M898mgLdk5HPQv6VSio6bNI3hqn8bZqKXpm80WEL+CGuTkXNoZCPk2NzmwTcAc2jotZNU
bJfF0Tu4DB22JPeF9iXF4aaO0mv/OueZtAtRhx+R8AXCOz9w9mb6UgqUP4INpkweqIDvkutIMphL
8mEEcZ5kXqQgwSad1A1cWfDqrfTMlKYAJ0HLUic0BC1KmLOjTx5k6pFh9lZxEmWN6W3wIwDUmbg+
AlRiZL/63yI4faFoaEAu1ZY2NJO5nzBA2nsaXWoJEAC+tcg6ui4NzEe/TFt+yedOxV5PR9wettJZ
RU93UMHvdYg0wgqT6soviHp9Kb+ywNaUZbGN2tBlzeoWs9zyiektoJfk0GC+jRseE8ShIOuSF8fF
tlhSsvGgYKaq7o5cD+uP3c4uuODFAFbUw8YXXYfcl3TSI89SWoKIJDl5KZqbd8G+wXbcb5mZUS95
3ZJIQsLrj2fX/0ergaH/JdtDWE86KZksnQQmylkXNA7jvjnwEFVtOGxU/ZJGhd1T8TnH1UcgDaiS
sEGlmYiHo38L/G70/eSTH6K1urfmkWyy9Rv81vSObB8TCbwbXDPq42njDQkYcAm+6sIhbMTgEyF/
YKjX0unBH4wjLKIOaHGhaPA5y100VJZsWbdfdeKV2UfG9e/yccYE9GDdPTLBydJy7EG5haBvA619
gGwesx3XxDEyrxBw/PuW/XIuoSn7lYzK45fNaO44wrlprdvPc3T/PlQ0mAzHZhhAFXDjoyJMe7Z2
06ZZ6ZaMt65lBjlsk+rFvDBtL1KfHepYBwuKNcJ5ifknV1AFmAbq4S50aHen13Pi8fBDowK+Xkv+
VXcKso4Cq/CZOaUihwRQAGTF3pri841SkhtHbDN9Hgx05ciuZmBoAe48Qou0DadgVZSP1hWKYoS4
RUrO2VrgqFyVYglO0Z3NNAb8f3nFPcRbpgKH86Ua2z9Xor5RtL1vhlSyF5UbZ4oSCzXhtCFXkaCG
+vKL2bYxLTm7FDf8g+/KGOCF7bmZ0DvvG3qG5NWuZoH9XWht0+HlfttxOtzgoc5gFEOlVSrpEYvc
5Jjg1jsYZ+BCfFWpzxsF8OY1FNDKJE81Qo+0fKeCj3QJDdCsFm0uQLAMa7CgVxdhmziXQdLcqwjd
/96FzucIXfNToOkn+ONGzVNyWlYUwjVrQP/tkMnhaTIrRUG8rB5uIshmBESfeCLP6knc9TXOHFrk
k/AuKEH8tEX0AJq8fgvyhQSLGkgN6Yx1WpfMap3GEgkuD1idAOGN4Kx6Deww/Xn/qr+UPKL8l4Xy
U1reiQTbwY6iQpW875sLiG+Ps61bzyFn1eyol6Mn9q5vWW4UFlQ29k8t/38jH2/upwxj+HXM9baO
1w4WFdIK+CTPvoF63fovLHa38ihC95GH7nPEsTMwWFevD8lDAAN8YsmrWYhdv3OwdQBL+/Vnh0sf
+HGClqJtoEJZMKvZ3dxbUpNM4wzP0uMs3DQA0/jl4bk/ehjuJEFSYclS4EISRM6oQszPec/ZsJ8P
gOTh3zUdS/LBgelJ2mRs2hA1GY72O9OdhCqPeLpGsTOgtxNSedAHLBbr/GhV4zz92kMSXOwUjol/
uE1SdKkDPXCjBd5tMbvbwI6u/f/05xQVj6zWBMdplxCnBSNh067xAEduHIxNnWoiMViXeKyGHnDE
o1GSZoccFJ07/pyMgwT8A30AEHubD5s+3IE0Wn0iCWuYzy/q6uncIB+x8l7yvoRu+BQTUCt8PaT5
p+itFTbb9nTcMODgR0qM0zEmjzGuFFDC6xqLuCutGT61bejBFqEfpl4SSwx/AIne381g4zp0cfQ+
gPvqt/Xe9ooSxmBpqg4cNgcxKLgo35FoMEyqoLw37o8+fPxV1MhNmHu8zf474figNo8tlpOH7c4A
RhmHYgmZV3XibnOkUQt3ADztUhHLrZkjQKCyEQej72KCViPSvXkoAfK+Yxc4cnriL9ZWdSxBMaP0
Z73R8d6JdZGbE4RYNWXLGsNBOXCfbSdjsLJXYW6ziuUsSYdI/nUQIfX2+m/2JI0pPFa8c5CrBqpc
wAMOBuTVVLBdMTbdmlz2rYnohrzMzlB+qw4nMyTAsj4SJ5d0/APb23q2ROJpKn9VNeJzfut+EsQO
aRnBmYaerF/jzXUPgCyCIc+XibwvjalDjuzO2WWHa0qduDLMRuGkM+FUlixoB3S5ZQO80vIz3ScR
+EN/yTcyOQKJk6r1Jtsea66nZwqWYxUozDk075gmwDxo7HpAlEeVTfNAVu78QGt3sU0sRvDIt6gG
XuaH1ckw50wPK3XOp2REwY2hU/yJQ3jaR+ty7pdUUBRUqhGnwljRoW85ywnahyNLUX9/22JNCKDb
CEsNuyYbE5S1MPz9oe/1zD9r3aHfbBHv+j8G66HkWNC93VO2fsVoim7db1WzOpadfpM2ysyje/OM
/nyTDgvaBqhT5OuXSOqX2/MFhxXvdGnM+W4rjmhPEN3xXfTOnv2eS75i2RXHhtvTU1R0J0P4p2cb
EAY/ynKVGXiCQKfzurW5mbqWeZzzc+8k85Yj1hGgqY0eVq1URe2o7xfQpUgk4krsa7NkRfddJp8v
Y7J0ju5B1dQViz3r/lkGAe4wmTPfOWe1Vow31NHAtNaX2JdeFY/Q9d55ubvcGPAilrz7YBc9W58H
IHQSPATOWhM7Fp7TNW5+0m+V1BmZSQkXTImDEOol2O+f5rXJ3R2f0tadlDqCTU1G/oQSo+SPN6uP
F6aWHNMvhmD48SGSJr+qAxxqqlwtMk5SZupAkXO6XTw9PX2cQirwpmjwfXRlkjhFuirekeucMuPL
OLqHEkoQrxDHBf3zhaASFY1Ji31F6oUaeG2IKzJQveriIh4TIFY8mFYai+8Z/qGw5mC0lYumBJUs
F55SrbHP1bSmY8LkSE0vDmAG/Sz/rpMLk5KNxmMN70pcoQJZfEh8adMeDLjbv+0rFUATzY0B6Tl8
9DDW3hm27rKZJfrUdlCR00Xp7HJyWHvvkzV/57e7SFXV3p2lohDHqVmjg5CNvEr+/Ns0IZ9bhdbB
z2JE65aidHrELwP/Jeynkkbb8vUkYYMTTpD2P+0NUCHfFnYHRs1jh26Oyw5sorWsXk8TdXXUSLfp
w6jDIGIubqJGRrbiWU1Fz4a5ic39J0eqygM0HFN8GxYbxWdQZdIbtoTfVanrB5o9YIRyRrDzGmyi
//iUeQO9DShqZfgsO4sCUQCTc+Pn9CDtJlce4T6DynKFiy+vy/skkoYMjuFNeCPD5El/45KAuRiu
BC9kcO2rHvxD4tf5nQPpd1LLfiSdoj4d+6EoFawYnzUZ+mTqE2Z+G1P4oXVsyRzOAZty+40f9ken
pvjIw2FUIfXfuNGowRUSmNVwqb+J3a2K/WnhbSD5yG3WvRh3Z7GPCZx5BbA1Cw3OAl5VIxLCmYU1
hRgTmCiM8v6Vwp8w9XW8j53T/wUp4wKYbgREcVJEc4Xg40HUUNsm1FAAh+LLibNSD25u1sQCQ3GK
UIRgK7VLaFAQncUN3i17+3ZB2ilMp27RY7w29pY2gCcJma0dgFU/1bVHtG8cV9YTrjOr+mG8p1R3
mTXL0hk6oabBX1BOKgYf2aC5aOnK7m6rmFC21fDOBpjXy1NCMvinxY3iTpT1sHGnBU7jwRK9VJy3
B6708HO6gfgmhQIOE915rqcpsGdMfo3v6PsiN1pESCbr1F819eMKfYfq7qDc+exxYp980S3Ao8SQ
ruTXpYhIFwgmCi98HS1oZZHN9ZEAfyYIcWUin827Cgn7CyUXmbeEbJmDDA6SMW+yCjU64jaBV1SJ
NHyVdfzt2pbTVrZMLxOEQ0JzQSPzWnux9VF3XsRPmqbMhYafN+5t080P7Glu8QZN3pJN5JI0nku9
6FgD7fMb3WOKb9IEJxFAcBnuXbs6IZ3j2I9vsZENyF1oHezEQ8Hi9MXolWDcnbPJ3iLJjc13zJ93
Hq8iVRgxVBpjtFUeziDzcRm6V45GXJn5ora4wsI+m5Z8KMhU3e7Xo+IknIWVKQN+y4rDKkUGHY6t
igErrVEQHAYaAa7VAdP4yYRSUpnF2YmBg9639OmhhnZdT/V8fn9o8wyRtGjS4MC4cxPb8O0lG7eF
ZKVMiIIglWvFes2gEViRGmEaXZbd3koTqd0DMz0t6YImF4O53uJI1nHSu4TUQlzrl11ju1sJQnYE
HTKfxvREA9WaKJfsqq6ojAqwJJOSyMcIRDr2RL0HsTqJTpDWub2QtfZ/7JADXne4YZOK8yAymR9l
zSNwl1IT79fgo1ux4TNtBZxYuc9kiGDkc3UbOmqpQqm5FZCBY4gPvPEOJhUTvkp18y1/7DWZ3BQn
6QjHS3+ZGD1EVVrjeaZYQN3ru+mmzCKHtRJu6yt6KKCEOfm2za4PxGaXggzZcFg9kkVqPoF+g5Um
r0o5K0lZFrLKmQG3WJFKJgtb2McUT2crc4WhhRO7foLBZEkTfBFRtN92HPb+q/hFBVoSTdgzPC2S
S/ce3EGmp/ZNNoNDE9Sidk8/ITdFUg1xIP0yX3CBapgijC/39gJ6/0sb0O5nt3U2zjFeF7AhTZT3
cTWXPvsb3DdPqZdbn+C+LANx68ogZXnnisINRJHTTuzq64sgHmaLEW5n+mj5RD5uW9M1uaaW5jL8
LT0QWdKbi8i8w7/y9FQdxlKFLYoiEHJ6X/TaaGff3GoNZiWH3hOMlUhKh4Gu4JNdlXcAiCITceEp
ND2I+L2VGn2R3bPI4vPqaeMy6NmHtPhunh4Ibx8pXYfz48mWR+KKNzmLzYVPQ7D9uaF+G7SUJBbL
G1CsBkSlOBuL+XJa9Skq6NdRzjwepxtamdkWEdg5Fdf61PZSKwbvSimnE8J9Lf7CIeub2WDtY+Sd
TZaZgC/+Aq9KP8gdZ3DM4FHQSIOOMG9w5JBcbwEXLXUx4KrQ6VkpFOYPFT48a/XGuywe8Zc8TaDb
m5gtT4l7FBPsUvd1TyVpr3svCWEkhwCbK+Zq73UF4xJMLnlLzkHh94AsKYDiLS106kpMOHKiEG08
ds1S7HsAXpeGXcHHPAtmRO3T9fOi1M3xff2hDuyxY6Vr+/t3zmLzyL4XG6z8jMTPjSwNM8Y9hGVg
7R+hciOOSZmWJ81hDXmnWaA0CZO/3Sco4cq6ovIRjExqz31cA2Sdrqo8X/Vo84T0skwKkAQ64l0G
kv6vDgV1LXPohmml4e/nzLZkVwvxOQtVQDfZZXJKsBYaCqrLBUoCVMpmRR7lRvwCc5Hqx1YD4BLj
UNdn12fgXRLxXfwxQYfKTvZYcn8tn8BNT9I7hIPLeTenML0bQDxJwFbJ2xJW284Bklufuk7u/yt9
w+Hio7tnBUe2tuWvSfe+tW5JO5J9wTPrcjtuG4UqJcjKbb8iBbqtSbJ82qPyuVHonaeaP+HVCjuL
Iey8DUY8Ugwl0UkxBZAt2y6eif5u6wss2JI4+YdvKgQzYxQ7U69JWGJPrAnzXUPKSO3S4ei3QnrM
yly/Al14tBccwCBMPswu0sWCI52iVaGHF8GAmwZvYvdYqxh2aZY+V3ERrnnI9TpfGCkBGspNjfy8
VELtOueM155ryHoDtZrUnGVaicH4DHuXUSp+GwcUTcTHU1+XoozfL9XktTSrcrk9kf+hYIri6wz1
2qbxIPvF63aidY7av6IzoFmn1XMN9rqkVc0rwYzmVwu1/4Sf5AXZCTELN2xbjjpyolX8+8qZxSu3
Lmz0u59NZO07ofvhmp5GwJ4WTu3pKAqc1T1I4rBOXknHcKfV061Dmfk7AuVfC2gjkNWP9ms+PVHI
eWQPAN2CoFieIxa1fguDyA+kqfINcl4vBHTY8XL5c2OVeYoUdzMWxY6pszWLGwG+FHEGyEjdRNLQ
8AuQaCJewVruPuhVkv3KAhi3mu1oYJAtxD8rS1YOBe2m4iUBM9r2sDmlVdmGItK9+pLvIMYaxwbs
3jenRj169XaVssTAh/JoQ/Mg2lEIGCws/2lbSh6x+tV8gTYTQklDe1FXy+HeHWfQizZLfHeHFi/D
n4YXz7j6bHGNcYVpQSH0eViAiC06+WjFc/QCDZnAPtUDMUASvnh/XC80F1rEHa23bo0r4bCcrwgB
xpxYqV3opmhLj6eOOxviqQreUMd1EgqQe8IqHfMs2w9IRZk1RZhFdLrjzM7J6VIKviR30LH0CIv4
vITXqOHR2WZO+kB+1VXeRIOVb1wxKEEMyAozBsci9J9I5ktEKTkayzgahRkvQKSrG3WKAilLxEJD
nF86JM/+L7joi8qZsfubghasEq4iHSk57O16rhweWdba7bcxOSNLnKgT4f78ont+T2tnX0ywuQq8
Qv018o3575DTqYpAtxCgY1KicOwidyKKJ9TSEwqdzEZPWAPqsyPixe6kpnm+V7KT3UO+eXtg/szu
h+CVcutxP0gz4tTF5hMEHNF0Yfm9P77K6xQm/3/swSSpqr9Uy3dvm6dHv0+g4evrEFIP+TJCB6h6
0eelg+zKUauOHtKgcSX8YWHXo1kt8UHo6ZrWJQXNi9PHjudSlBsa8RYX/pp5plyeGAG1ZAkD13ne
1ej4pcgVMFe4ESXOk3DG4LfhgiuMKHSGO3g4H91AHJS9G7feBexNW8tZD6L7P/quRVjxgM7ZICY1
YkeulsxrfRGpwf0bZXX/1YXdIHCytF3ix6QLkpCSUOYfJ1BTtgvtIfw1KEvMRwutMrXPqP5WZhyQ
5+m5h0KUmD2x6xGAZ3NyNl9Uzfu4neYwqo61aqwFEh/SeXhOXT6vaEVctluSX8fDXv1Qoq/VYfDz
3r/g9UkY3fGFHIn02827MCAtWswU+cROGb3XJBjQhAGs7saXVWvNso1fykOIEavRVl+fS0Rjzst8
+g0Gvz+489FsUsBevowQ1MPLYjvfm3DWcJ6Vk9BEn7DjNjXGSO+BenMfsmDfVhjjcgKoUB/g+jSW
mCrh6HCwi2ZBwfhvKYaOYOhTNYxJrss7Bf1T5xQvLV3C7gp2kWftwZ73VR3F+VZzNE0AU7skPzH5
mXQz0lZAJwx6GITPzfhJVyZbEKcQwTmchrpheYJ2Azcs9FjjevCpP3sIaai/QrLrb9HqfTLDLGs2
Tzedx4tnzlmKefNaPz6J98Ss+3/leX+l+cLgxn0hL8PPhshU1TPEmDEbNl6Zil8oNlOKDB4eLYKP
vXD1hICm1n6J9PnRDcAkSJK1X5U+SV0FAPRM0AixQ5qO/B5fSZLb1knSOXb6mhHUjpIUGR9s6OWE
jcBkYhD3mrR65cc9+jJS05Oj6gvDW0G3Usj0+oqh8UqHa6ygLhbEPz28soHXXwMOaPQqSlITil5q
ehSsqAee3jWzT2jrvO+7uOTtbqxyyfCHpqbNFyIi2AFCmpbn+irJ9m2SrgdLc7jKB0suVXmBNgTi
TYA3aoFANOZ+TnLY4weuGtkFRc1YDKa9vZdZdT18U05gov4kfNV7TIH0MRvhLZYaBHD6qvqkGx0p
e9VkBa5pg4030PiheARV8f/0J6hHHQamugwnX6C1kZHq8JI47deiYJRt0JugkkNEWC8AxH+MDNhG
JU+m3XjhyrFFes+6JYDKglmh0WfoBXBfJlyna2W7uBBChfda/5CcPSiMXZFhfk3nehsAKKR4zlAF
4xJmfuOouaL2LjUBWDR2ZpVFQ1b3eh1pLUoTGKyd0UGO8+RnEHZnUOCZw5Z6+jRZZGmRL933WcVg
EJNqYfyr2K5ly6qTgx5osy2b6HLwSYgbI314hwx77LHh98dg0pTFH05JTk2lEZ61OWaZWGL/tNFX
IBqCEXs2BAnVbJfl27h1wiXZ36ryYtwX8CHQWt3dUTfks0hTrOKRbkhYQrF7C1xHlAvO9ode490B
nZ10nphHwIltToV51/yGUEPmwzCAXsW6wU+Th3xce7OB3cFoFtqu7uDJN75y0NIYaNSl3ZVu1TsQ
/vCpUpyFnctrJfdlscmvBL8m5QYKRnpsCw0voVK3WFYe1qfzy6biHgNeecmSpyRannjgyxidUkr3
YuhmLfTlD7c33pa/si4Rbnmq3R6NvRailaIaLa975NWqrk/PX1v+ixbnhVwFpzooFEl9A5h8kzkG
dS/XLYO+JWXZ8/busxjPUu62xF1OlYwcEkDbeiYjBFkciGijgGDa9VPNcbjuK0tvomLhaXOAcd9a
WXOJE8X1J6uCxu7g3B+OZnuCfDKEXi9MGzPOV1XE6A/WG1pJ9PS3nuZLJQI/Cw0ko1M6jC038jA8
6+Rfx2nMvmr6Drh/+TAOSoW/zo6OYRDybepKxtwDCPjSldUBcSLjbDB8xuUeakmUt51WDkqnEeOO
yRbgbNJybNKtDou42LUP46aUIq2MvOaMk1nUcZbJ8siTdO+5OA7fZDGKCQD4hAC3gxANiZME/i05
0fCHZYuGnCQC2rk+sp4fphkEOITnWdJsSNpnDPVhg0wfCfUZ2ZiuVmGbrQ50z6pIzB0YA3CU3Re8
Px1fy56S1DIU95nfiIdl0BUN5Lff8WtOekBVHHQL+JGd79LQx6IalQeW+o9xvNlWl4spVb1iyuqc
ySJsA8ri4RfSIPwvf6ubeQRe/cpjC1nkFEYV6BlPZl5aeWJIM/iRg9u5DypMd5lppwLs6UuNiuH1
x0RI3iDG5/tUN8a8tizTxnEctBEwxuVErOlYtEgR5mDyh1T1Fk2gsaYgOL5fpOXaj2LwBbKKZa2y
o7KlsgdGtxxco8Uh3eLmsU1e6LkHdcpYFiIUp77H+bujseA7AYI8x9M8V4JJCP6Vwv90c2W4sPWF
f587qkfgWstg0o7jWRiHGIhIL+FzxbOlnXNuF58tIrbPv6p6OGz3unypCbHGlkGlwLSoNcdd8TUC
IuVRwrK5bZVGxaz5+1o16U4fieuGrOM59JCGosKYlAZKUl+AlS5Q1SFhsQoB+oaQfdgnMYwkr4RG
bkfHiE67rszUwAObuyWsECRczH1A25Ud4XHdJXfE5y2b8GVzPBhfaoD/AfS9qPyrZssWIPtkL8ev
cSKzjLn8g86WQ+LxJ0FEu43cETQjA4omZE0ptffwvsJJhYp1AAlCFbtR1oCk2oEbVXALYkDosWHP
RxdJOKIVo/xQOMe/+caqF44yNojmhzN7WpJz6WpdDqWwPcc0wIicG0MzYsA0vHXn6FU4rzXJeUwk
QB/QOarVQuVlvrjHDJ3nu8Sbcp4vQIfXaeSoVvzO+/uphybyP3mRMKFMe4M1ZJ5JdMgtEKSNO6jl
qLTPQBzGcrHVPdmCi1miGWsPh4Sp9YJX3+veut0pkFXxMzsE4W9WvrIasXjkoUsK9wyueoL8gcOy
uF4YqXwX6Aljp9028OGXRW5hJas6JU+d6Lrsmd+AZ19jHFpcR2RhPbTC60fvApyxiodF9xfHONGD
pRQdJC0tnYdx0YQJpggRzZjc/wg/LdhcN4spiuhFqx5wV1PvCW8rKAcJJ2/0PC7/UWqltlSky+Uk
Me4ckAYVFW282wo30aPd/RYyv0UnpaCgtP0+sq5YBaIf/IjGSS8fEE6sEXQnamF8e5M8ZoqvDrAg
28RtXXK1PHsvcGQSPWtURtqjSldCfrTVjHby2Cg3DTFYDorAVMk1LkTgfOBAM5uDb+VNDDb3zsim
wYBuSY5LqLxXJS1IHWyJNcVHZLoyngLoP/9Fbdh4LxUjKHoHDrcgjhgwVofIH+2mfqKoq+nMqfdw
YzpaPMBfZ2wb8yXhUAZDlJEFge8rgdSz2lcgqN6onK5dxhDVuck9C0qN5jSWwZ2E0AzwnuzdlTf2
XpjaDJD3viVB62h4m0z5D5g1qSqqGhC4lzd07DOZOpYf1wWyPyIBDXa3Tz5PducQ6l3a9v0oj9UG
RcTDQwnbd92oCutnkMb2xlexBWmqaa/H/A/oOl5OycEUIpG/K8gQPbgUY5UIaM8LSTSn5c5c9Y5m
bpLVAcQ5nLfGCKeqqHP2WjZYU/gQCWdFBm7IZT63+3N4MM5ZLc9h7VgQihtBbaEqDSaBXaUusJRw
1Wu+eB0sMaGHu260MCBDe5OvML6KtoiYVj/lLMclfR3CcuI8rDnixE7+6E9uN1Dwfm9bpz1gLCpI
h/Ul7GDYuwpG7/kFvy6FtgDdQvLo4RyYLn8KTKkO23WNsVkVoJApeOVgjK4/KC2GRlIzVQ0kg9j+
wFbymyP8hUem2m/JOjxY3J9SHOPvdJdFbL4k/SzwQ/lPwawN2ozr5HRnEWhaAocUHT6uLfZk68w/
xvWv7U+bQV6Lv65Fuyy2UAxqHd/gqtgWGfe7Rgivd+CvUQo+zkYkgOgTNuLDZOJIiXh4P8W4bku1
w/aZU3VQHYdIMPPr9WUomwsKT1nq2L5Grms4nu1tZZALlX0Qg0EIOBNc6fqAH5Mz6uavrktJGaT9
J8cf+wpY1Urg5g15JeA6eRoG4LGOFhFLDJU7uq0CMm9KhlgNIKN1LJ22M/tpZk9uVZD5CSmutMp4
K3AW2wrlH9abcqC/XJNH6qrd5gbHN+m+MmlLv1xFSCSUUNVte/s416A4uqbeqh0XkLNQXyfWJdUU
XterRmFLS8+W7grx/NYRZLZ0RxiLO/AdmRWfh9F+rduVXGdjxF41F3jehKYLO/trOhKecsngXWew
FBp/aFFuPTL7/ZW9UaUBqANG5W8gAZbkouIxDAuE39T/HWQBsMwanLiVZV88EzJ7W4Qh1sUDmCfH
3HAaA71ajwmVr3HJx13FE8Q0PSRLytK1FhQkf8H3GS/U2V+NbF3AxbezDkycJhTQSRuJszD0uYTi
zVX3UwrYWrBerol0BvhDDrJrSHaoGRGq6XZ6+dMXA0lLDdvPuysiKbTB9CSFDqRco1qffSL6HU+W
nrkpGkA2YTU4X/Xqf7xg7FHlUlUgp9ck94UgY/5iPafa/QlQ0CkZEX4U67fneXk+VxCpOaf5Bbyj
/rqUcvrQK51hQ3uwV7m/7Qn0Cx7N64ZZgrX5cD2i8Q5EDFA8T7sFz1X5HMSTE6v/a1AP147xQhNy
xJAU7ldVrvpt/ROE7Wtxk5MQtlxUjBdCEdkBfOv3C+h5Klnz/B220KArK0jiIWKrlM/aA21gOuqP
2XRn3nVKauciw7qCHQmawsgYqEfvKtzUSBY+ktPcaQ4bAZwfoS1PGJGiddn3qp9ped1KxDm0ufjy
gFaBzr3jat6C+StvIDG6nhs3y1ocNfFaUjUt7PdSgb0oasgDfmit5Os9L1g94i98VcJYPAPVRsq5
C2FZ+ZJapm+1FOuWN4G8Bb4tXFSB5KqiEHup9vWwO26Dlw1RfQoHG36Xe+AZnsgFU7K3wBWRXfRk
eEPnvGqBDI/4WWnU5PkR99+uTuzeH4pLLVU9PrMZICWX1X+zv3+h8Y8cBpPZHv0d7+rQngByCiyj
zJI2wccdor9Md/jEFND6nwZuVbCTeZoyRncvWZU2c8VZol2zpCe7kjXm5UV152u0g3015B2lQJwL
G6ltW/awWV57wVmZ+s9aLD7OE1dIHlK8aTRy7VGnLLK0sNcve89YqrUsPGIhpIAigxmRTPsOL137
170GFRS/lSB946iN8RFd3RHcOhgVIIjxDhtgnmURgeA1DbBUFiOt7AglyHfY897q1Zy5lT/ithcj
BNVIYkC8Is38iuhc9p/eobiCbsnSU//yF5FiU8ev52WHdg5J852GX1r/u5BrYGXQefRDtVUOxsHa
7zqKHAvB12Jb59Gl/rqlNba0ykiJb5F4Bi+1HuGDQsp4278b6VXoA0NvGEZWpDmXLIyso61sSbRa
E1Zl5J8W4akME5olh6HXpT7YSuBeMHnIy1MQWADk02tk8O7DHVgfMHcuBwyQOocZXzpdt0qc9iT9
vigvBZTSXf+pxCqHqR/BUJTRp7TS0iIc69opLf3ZiKj12ymQ4pRwWQR1h3rJZXAECYPP4iIK27E/
yL+pBwL4A8va2v6GOmmpriJOj/V4XFfB7UckV4FAH+Sfxe/9OTyJI/ttVfYn05RfYTTibpGA86es
5MKAgmWWh4FK72Nb3xolJ+dk+82E4X4wyFb1+0kZNaQLdtxikUIalC2G1cuyqW1Hf90ko72qsZza
bpvdOkdgbi+pnDerz7f8c+GOS/bWBpIsnF5EJ6pwfY0Y0YStI/Ozsit/bsBolaZxjHwZfq7bY+wZ
Rrbthm8LlHlXVQ+fhHR8lrPMKwCqTqRcS726yKz7qe+FyEq57dut8YY+aAz8FIFdSTjY9IOfhq2D
aPmWoM+2aTfiQkbi01SnSxd2cm+ac4VjJrlf0Cr+s+A7XXTBiltFj4+EGEPfhy1/4Up7hF2UjSd6
eVtA6OaL5h4RMQ+fk45it1RVQxd4DCPZX6m6NuQm329JlwzuDgOnpcC5uxJZUbnOFFowsvfcOqTY
yeod+O/0vO/ShWmt2sSs7+lR2kgYI8AJDK1dj3vhH7s2b20r1U8Rsp6C6TH+IJGOR+nb3S+tKLmJ
N8haWZcbPQNKu9ZakJ4Tvbf8L9f2wiVkIPvWvUiJyd4FEcgYYj6KDRfy+d5cYsoV+OCeXW01GxLV
4FYSMluo+WXZspQNB+P149yAM3FeSceutVHTPrF5OB/XWiNxjMSAgAgaz41bApE2pogajcGtNUtJ
CM4oF2A2MuWOoq+fOD7begKdSjdM3dL17jVGcOOmUFjM3xwOXFZM19R7AkCnjxmr3jbjFsKzeO/N
e8/79/3pPuYv9ALKnmGvWd1OW8TFgUc+21DLFCMZ4HdDzqJW/U/Hjl7Xj2Z9rTk1plfLP2L7S5nS
tbpX+Jw8Q80dGuPnHJBbWoA/8dvn7un/wf6zWl4dpj6mMTsoGhSGty905vyWvygNvXTsNNTfQDm0
vUj8lH4O1ClB9ghEKfjdIKewZbpo5rSCzZFET3vsYd6Zo3WYkDYDTMeZyxwTsXszrTIvC9tMfm7L
C4suJMNO8DctCipHGYOICFwKkadmny29LhsCzdxhhEgsMBwUcxT0iS9P69XZG5nCTYVo8J7K5jKd
w+9Zyvf51BqFhM5Ry+2j/8yRBprELSLb6jBOP1oxzpfyzA9Je5n5ShrwIgQan5f02IzXaNCMv/f1
ADpI8Wms3tGzQcy1PJac4DWr0EQjOm3NNXGOY15BCdNim6EIt4BexCll84zdv33YIYSlAGqsx6T1
nq5Ogto8Uw4Jor5jPo8Nr5XPm+zu30baTO2NzSCEBqOd+MvDT6l/VfUae95R99ikhtWl3NgAtAxe
CE3lYa9YrZZMtmvjQ9WppMPS1IDI+ACPhU/5CpO77P/1UxfEdxUZu1Y9c7fZuM0Ngw46FHRRoUH4
rUN2ycBbhsRquEs8afgmet1VnsiuPZ25AYSSZmxsxAy2LlE2QwiKIzEuiTiqROCp/IKy7fdWLTlh
QW4V0G+61oDG4o2c0u5IZYL7mJBeTVPc/4B0BtsB5H7yV0bGgtbCmn4oTizgFYIfbUb7rILbuc+9
AonaSdvi7oWmZf7psFT+xAQtSPTl8K78IjnIOz2mQyT4QxwlFCgotug+W8eg6hygH9PTpbfcibPy
r7hK+FDxNk2ft1NL2QnqBmeQxL6BKsuMsXMC+MBBlep/QyGQkETJPw+o4IkfGXbsm7vrlA9mE6Zh
4pt9U4pHnG+Iu+9LLhVzv9M3G5R6OMwk5I69i1zyRQkoODpIdQV3K9W03NnBoTRH32nsZmIOkAUA
SxfO+cpmqo0/882pVVYhNwo4RHIlHZOOgkAjNw9Yjt1/wwA3zAH881R2jZmg42M5lfPOhp8pZrkL
3jirEfk/RgIPiSOMJ38x3vszxjAUo4W/vKnb+q9gnh2CUZP6YGMOLZMzAQZMPrOqn/Ks8ZnM1tAg
yGlfr4hJG2vVYMYWFe7Cy0nLk2HrV9gtgZi5vICXqmxkCJIH5dHpQDLqY54uyIWa+NVZ4wPZzkOX
8vKxlz8H8ifNxCev3m/XHNMUIs1QgGrdKFtwgCciyokU4g1urdBnqoVGjM+5rYf4KCCmVwNqHzoa
cxfZawkaR2v8Y+qWlws8gbg/B0+2VOYyorKfHJl4Ofdpia4dpdIybOeggSv9YqaH+fITbIoOWkr7
AC7FLwcOXqgl3b6xIAvJbJo4fnf8DgxDxESZJht9paLTkKhcqfUs900KK/3K11NhUqDVCfXdc1ek
26Fab7wPtbalU79GnQ8FSQDXtjZay8s9VHYLrTQI5cGfn10lDQy5qHk+2UKfjRPHgiM/C1wRLH1M
CdlsewOTPJ8BjO488kXcXdJrQpX9oNgEAKyUdv7vn7xapueYd/Aq26GRzlwmRLpo8jrcNl96fzpT
kLzNWyC5BJ+GLd1hI5IyzsaAXXZuPiGk20XzvLff25eofLngCIZ4K0EJd6Piwsku0lx1YnqDOBO8
RU8/vXgrlb/8LBhLuVXwNS5B++0qxPMTKW11ZMz5TF7Tf+mhcCqnu0Xi8dLKE9No1MLsThI7NLR2
8iT4OIQC0O+8I017QswaOddD+nikycAHqj6QUCllHtAiCu9D+v0TRDNKr4VnGJ/92ijJjDgnKmC3
IBfdVytu/IKKaNwY6hN3MPT/xi2U8ih/kCD4XKPOtgfEM0r/T8MaqneghX5LUB8YsBM5KaRfyDga
EBrkPYY7QaYlkzlYfs78AIPgtlYpnIDC35AEp5pBDIec08nwnXp5C9gBtamVFOMZsrL858HnACyH
MZiLZ9AiNGncBgQFo+msau7vvgbq/Hiny9/83kJDLi6IE66N2kuzj4gi3w/f9LAdmEVCtK8e/NKu
hY7gIhhYqUdcqJezPbLO9vjyR2D++LblVVUZbIspnGJ65RHv21dmIiIbhQJ43KZUK/A96zxfB1wP
y+CCWl1toibT6lQkoB/y3nl1l7HWzzGv5zj0hXsubWRJKTvE9vKWlC31WwrYJ0HByRvcNoFVoO3W
uQBmarOLqjYUEek84JpXv31Ze0cfpXRQtdkPz2qJdmbhQZVK11mnYGr7SKznYOBwOthRLfsuNw+Y
mkGi8W5SbX1WFbuk1I79bCJu7m51VtMbbBCTBHqDNtKOVaYl0SCKQz3LkXQwSYrkMR3KRqj4TgkG
nuny4/libJYxPsJPvljjgeIM9An9QhyohUgJODd7XKkH1T25mG21T3UNEWx9Qe1JGVHndUbBPIHc
ByDWReYxVqw/ofWitRiW+Ayh9V+IOfYg8lLteyk42cC2gVUYRN0NhWHyHPI6gFgnaOk7N68x+ncM
thvSw4rmkbj1d6klXLurY5/k+kMDFYO+9MrtcTF5a2Gi26MD13hnJ2RDPTin4LfX8g20RwnwRu/M
unN7B9NrCP0LGpTr9IItFakFHzdwF8ZRMEebSN2kMoSIQHFqxoddxP4YdqA73a2sGDPVPfIxgrcv
J/w1Jcu1GY+tu1qQB6jGY9L791yTyLXpJ1kKuuqIeT+ygZQCcQ4Clil/jPCG3xN1y6e0gK/hX7jV
Mroh35fP2NmxO7Efzeyc8xyEPo9rMmRSYFZYyHNMdaQtKwHBwqfYjWOWDJpwiR5jA93AMT8ffKaH
S/BpS/ZfRCNVcN9C3InUxMPZN4roC0zBHC8h0GDFsQmIj/ZvTNRS4xHkA17y45ZWalGpmlIVKJM7
LKZV4mkc0fuRXuwplZnAfZgunHNGj/WH9AHIffpx74L2eb8T2QDvn2TpdDZN6egfvkyuDpXP3uaa
fP+sCvgXxvAZB/pQrdhckTI67kG/pYGOw4wWuV6LzJ0Lo+y2d09oQqUVKTF5+eLmMuu1O34+SHYM
9WdkSy/LRHBJxozH2MHXQ/6CbzbXH2I9ggHthObUmqJ65roQSxZf3+fD65LN7ZCOldPRsDXZBHEy
/uaWYkk758/5L1rNNz1XWEnmpO7ogYGbeRyqvYi4C/s4cFZIORBcFEhKgS478OyMQNKnjiA/h4h0
/T7Z0crM4QSVN8d9lA7BF0GEx39rKyDEsDzQ5QBo07QK2QbtWYtSUoctkTRbFbCg9/hQHRCVPQiO
Lu6gmKLatDFg69GhFVXzpv2FApWo45Q8UMvoka6jf0SAoNboC2LVKGcyd6SA8o9rUKWNPnZrj+rT
ykoglUUhHk5vC1mrXGMaiOU0y5bRfd0wvjI4lqdzs26z6+c9fTaqHCHljUkw5rFzQABus0FSi0pY
LCqMbi7UJyCtj/0mtk3cChIJQRYm7kgeUZmu9fei6Sp6DGCSH0G91RG6gIp4yqM1+RP54ChStLUi
djLrDAjWku8W1zft8N4XwtFLYTxzK+D8810NCBC+xw1mnTdsMwYqXrF5ySEVDD9RnUVGmzeRI6p9
xzjMZlz8pF5LeZJEaEE8K0yHdpSdt9izOSAEUbnUNQhEjPsf5KTGsl8QnYjnSwKBjoTMmgtwWS/1
YREmMk56Dl2HzF0hod7NLmOdsmmRWwlORc33TZv7bCcut6PYPSDN1wF/3njovfUIaPHWqIBgbi94
JZJKW11cH19OvSGHgfogYjH2Z9nRu5vbd5pvogaCDAyQ5IWpRX3fodkBOU983uRpZF8uNMlRr77p
2gqFOENOloAdSi5iavaVJCRQKYsIZSspjqIn3K9w31d3H1DWYnI9v+rn+EuquDVNX5+N/YexfOta
+phoKrlPGGJSTDkMSJBnCxQ9icB6Mj/G3KtNeo9SPBwsvlCDbSjvlixpUVNoGunuHQaTISnaxqBO
fz1O6lwA52O8xbet4F1fPbSHQabf8h43hFnu7vuDGjwXvCI0fBQKUYKm6qdOELhLRL3FIvWdA8hI
X4PerGKHUuIzup/fE8od+pAzZTluBI0t1wfSX8RgLbHKlfp2NxrsmSwI5uEuqnsgsoYsXGa+2G9t
Z/XAYMdMX0oUQSgXy/+bHX65I856pevzkmEzjx+g+LFPuXYDyhQ9Uy19G7SKMlhdt+MhQxB6HGFd
SBCU+v+xbLE2b56PpzZsa0wHwIfTauxblYQCmqFze5MGFQC8OfL4ZtDVTYHw+5z9/MosPnTJ7oQx
JI7mvIeO5cSNuCpeWnR9GAs+6v5gzdMPTuLICmER3TYZ37MA4r5WDOsf+81B2+B0pwrFDCHygkAK
9cTL3AO6tEcwIAQtfonlBCtyOddresa8Zidw8Y8XENia/TfBdVhWvrOwfFxbzsNEIOqF3YHB80px
Kt2YinX35ptmdpFok3J9UQFzOGvb5OYyaGuvnAsxG+yFgwbUiVLHZ9iyrgnJ/KjQrxKDh0MzG8Wb
L00BLyOiF/wQiNPzmq65ue5iG/CEgTIH36nXASBBSofM6a8tZQ1gfGG05V+ZCBRQDRhpMjrogPAa
vEEyU20ddHjWxIGlA9PXbTyuW78+H54d4sdmmnDGxcHL86Zod5/YcaNrgNo9rFj4vtM95LlE9X/y
T2/3353gUCtLD2YhEKYyEjokUmBNqgJU+ki47ZyR+mXFrHGIIiJNJfG9+10rAoR5TUspjx+zIoo6
sROpWhECGRTtAAndhMuibeyvaViCXHiloVVXIIoHEtIdnlX1kcLMG0FfjTo1x1T+DK5q6A8hEtTh
+HR8QNjhRO3DL4gSwhE3Q6JUkhvJqxOzLEjQVU07Fk0NUvvIEDvyW+CavQQRVK+zZ9LIF6xbN9yi
qhjBcKH4FsorUtIm7hRKUiwVztst5hA8kZlmp1msDtMbnWE8KEE1q2hdxaaRyeaNZhzGmzP+Eu78
sENn7OP32UgJBbraj20oMXozMgff1oprqlroo+HCViFKpYJPotAYmPORUxdGr3NA1N0bOHxAuLvA
wRvLuS8VOzXMta6W3yqXnvFe7m2CpFlVs0/W8741D8dV7OBFQ8FfoBJJjih1vm3WDuD+21IcwUjJ
kAwi0wrNM+IdULN5x+5vj3GYrs9sJvpe5j/IvA4eHk6Hg2QVuxSW8buXi3H1dEkdmyMIMBJcMkAJ
sljT9rdnLKz9oLjo2dYvUHQLKD+l7b2dmtUO3JKVJR134V7/YpZtFwnnTMiXtLEiLD79b8+f1Ce7
LwWUbSeOtKilckDgNuxeRY/cpiqFawGwvISASHafFIizTxrqZAI2nAIJrYUz36wE2eJRkBz5AnVs
BKwTZfRmFr2VNnRSqzN3wK4keFGCFlMD1sBrKLfbumU98kbUoP/k+wgeSc9Xr75olkOxaDzFVumH
XUff3Y43DJLknASr/UxdD8MjaMMz14ChL2ZMmdVsEKkifqxHy2tFnNFW+6+NTT51fHTMU73//iC1
TAvqowmFS1MIzQrUAlX5NdSZtp7t0+vwdXGLL+Q9IvWRQ60njSIDo7CUq/E6eOzpqEeNX6Zwat0I
XIW6eKW+8DXBeVJDPsOxznGH9N1FucGF+qliDkckfK2DsC6/A5lZfDuCC/78FMTWj3A585HQag3A
MFU6Mj6o2VjkZQE2NRU5uHq+Hqgbx4ZPYRpDl67oEAmZXcCtBPmXJz25Q7nk4Vcm5TC42rhdF7av
++c32WjnGeucNgMqCM97UJqo63/rq1lGm06u/F4jAJvhYoxkORRfoDD7p2mBlJl9DRWNTm23cglC
Iow49rnPJG1QQMdBNE5F3cdi69KbnDWCFz6nnBoOmA7Sr6opeB+iluI9YOOUmI5GE/Q4iN+WyWwk
b/kiG6mYHWEIa4A+Zi1ugiW3khc8jA3SW4L6yGTegkQKc0jqTYeXo/GogPUtOUKyzRDPfy69AUSd
cHQPrMFqDPOgj8RdVRwsTvAdnmW1JXFq7yu1B83BCgIXanBcPZ8QgNnG77mOoJBEqErgLM2GnsmO
xsalWTBWEofK+kV8RwYGSpepKg1/TVyegAUEAdYewuw2ul2glUJTPzYP1A4yQFlmisyAAgKdwuYu
KPmaizx1L29cr0+oK3sYeE9V/6mtHslnqxG6IBNxanej5REXsb1IpYE6lAwB4qP/Q0Z7jZVoRQiI
A0dSeNKSZKcPUKe4EETyKr0l+KrNXvVjMRpKNnW33H9dUiNNueSHRqmhlFIlyq42nnR0kWaMjmVU
eefFO5tD1EiWpUf0ZLHJtDAwD/SU+WbI2KSFedFGsHOkIUIckD5Lm/2PVOQvGXWTcm9Yi5IKUFJu
GQAWMR42deE8clgwfMM087/+k3kJSoZJCyh8pA7gODoZkeQyCuiGV6yiEfHKUnCOnP5LsPMj+h+Y
YvaNvOrtQrPb9AAmw/mDi9tQuYC933CCxg8sXpN1XzYXw7B8VzpvurDk6cd12Fznl+iFoxg803TA
1XElC7ri5/oj0HMMYt78HzrD9CQXr9Lx5G3i/ICDlQfNRiUmyY7q8q300mZgpCyyGZk7SU908dRa
qHhEeThRBl6E/2O6ap1cP/sXSLFtw55nI5J8sabYB5w8nzLiojjc5kBxGaIhqaas7/DEa4ZOhivZ
/E/aSsQPzHr4Y5zHJxB/D4YLJHENqMCbGb69LT0VBaLqs7UynrCzLoYx2ohEr6FPq54HR2KkTfBL
aEGDyt9v0YICpR+SK0zoB2nvdoJUY6YV/x32SjAyhbC8elOJ/UDfBTxddsJurZzSQQFH1V+oxmd7
rcBfePMhVt9HaU1zlunZKaRnGBabfMQXsEQUDZNjFH/53fnQX5vm0+ieP9tb6PAx2fW0C4wjJ4z8
sywhVGyPEXEUQmvX7Z+e6m+wFybU8u1WwidvUbdudZrEyB2eMhYwodphIescGxrvAk9PDgf6ZD7R
tREBBZ8I4AbhWYASBiKFwq7suf7E3YSnC69fsFcGpH2rHacwnFQ94HXmrie6Cf0bAgyRThhvoVH+
YVX2JTB2J73tNRnW9FaMUyEW2UyhGItCTVGToerFKblZ1PHtAw0bfTuIp/bL1oUeqYsB3acH4Qcl
tR0bvBGy9vwPR/BNaL+NW0dFwuWxRFF0W6v2BAxXiJT4rgDfh9PpS6vARFxI0A3l0efJyjDrFXQh
c/Gf3sI264c3tRDfmmwN9c2eejla2YPt1diNQ76WGWxhkTOhPrLvYhC485BLlVZrP1nNx4tTAvlO
54BUe8DnaKi0zcfyoQXoA8etVZOaL0ioY59myzCnw3vOonQKzTFXfYrClo/hZyKWiGMmuOg8Kvk0
JXzRK8EVwAWOfdMizIJxGYLjjXOW8fTKVyiXHV0zQqPTnXU99TAWSmkeATIu783M3Dj/xPqR6P7f
XQ1GSExVRa2eVpv0Z0erHZT/HJSpjRJnhghF4fio5V2tVzGvSr1a+kHtb5PjdLwnlYdqjtKx3Cih
4luAPztWucmiDmapaYHCuRK7x7CoOw3r29cmJXCLJ7YfzO79YcmCTQNygE8kM+IT1WcimmtPoPW5
5/4FQvT2dCzYTZ00l5ACXSyPKI4t0VhV4GHunjFaER64mdbMuHka1pzHljBPfA29Ir7WWJlTtAZO
Jbgt/AQyMMbXQUaJwNS1Jvg5SjQcAP3qEC2g3vPvXENek8net2uIOJTn9V2IIGZUKk7T1PzQqZkk
P4C/UaboL0hBIZV5P4aBrT267wIARqwH3PLbouO11b4TwPYiUcQS2igzbOFkYzewwS5QZaHzLlxF
wseJIbxWwgVBhERk1iF08rn7smVjTHxr3w8siR37FYb3N6TCFKFlBSTn3MfDYsFIS072Q69vpJCL
kRxbKsvd7AS3ng/eVLY3Z8z9Av3xz9zT+ixF4bP+Ua9eTmDHgjiXFOJX2Xle3LuDjQ73ZQ65AsoG
ttNzc6CzYKc/G7USVvciBCKgtItYsslC9UnyNonee347lTBmraFi13mv5/F7enmH7tnOpLJCtZ7h
zmTgMVxKpUI64BC2P+sb/A7Drk4/D5tRMolCRnPhDwPy0WdaKlEy+7EkS+goKMzKMfZ6qTkdfwzg
Gl2TJtIEFn2XZs2P93Qb1RrEfsKf7Idpw5KiHjnwYQYEWlkcywYaXyO9+qk62ibAZrB/6IExhz1R
FrmlCIotb3FAmE5O8LXqOflEggKyGkN9RnQdJW0HIgZj/hFLU9GPgOPJ0GeQK24t6x/zDGwc6weQ
/U3Eany0FGqRjGek5lAqL+gnQT2JDWLd3mgion+1mD6HwV2bJRALKsuiUMkTwH2bMU6jDR/nikel
Co+rF5p3/ypGl26+lRjlho1yHY7xQmKrfR1cuIg4N76jf1g9maZLlUPZoUk0TXy8mukovMjvfhjU
TAU3NJlwZZnYJDbsaB4rn02b3FGqRvajPwSg1IFXjI7jg8J8ZiwSG3FC9bW3stE0wf1p5Z4cjuH2
yyLoavZ78mx2qTiMzGqxMkuNVTFrxHkLzBV8xj2AYgc+CnFC8+barb1sN68FKGJbpUowxmlHVcd1
T4sWSZPeBRYEEqigBg9mgluUBkw+iy0M+/Lv0lwLGmAP+A9lA/Wyw47Xyg2KCUPiu64h40ffNc8g
VMr0NmaKlM0cdTJDr0Nxwm6XYrE9si8/KRQrh8OyLu9CdAvNB3YJG3XkYkLInsOKK+LcmybjfG52
sp4j9apLOJMXpdQWrkqn5hixm0vhdJNGb/MsN9m5VA6wd8spf5dQ8pSihFGlEXRkg/N5YdsxIH11
83NChn0dlQTHOkqWJDisA5BlMVJ5/spFTclw69pzrUugMJzC0H/OPZpPnR98rRzl/BMJvUNzVAqK
qDbOctzF/4fqYrr6hEBkA7tBodmCMEesSoERwc+dUixU1yJPijui9S0At+pB5B1e60nEcYqIbtte
zmZ1QDZ/y41k8U9Bkm+oLoLopXPP6bVRTVKhn5bqsBd4VDNaGsZGXvqnwdBQvmwg8IJDwj7+Dt3a
kTvgQ1K/gmcLlES2le3GZg2aXrZJMWbkpCJrEki3SQG5FeZzkRjCwDhap0t+DMd1ewK8tGjFwubE
5h2dumz1KvRgs+IE/aMRJQCnXHQV0QnACgs9jj4vewAZsHX8lUknljlX7cZSY7SMKFLDpU1CblGQ
fcgF+dUSss5NUOD9NjqhZPJWaktL9bZy721pOKDIqwhjYE3ikFYwdvsXdD4oFB9D4esp50Or1/n2
McKlqiAjo0fJBfktfeqo7tXwQZ6zDQ4O/bEiwcic9VWusaZNr9QWpX9lXw2HxeQLuMZ45MoLmTvc
bqMBHNbxcT/FTu519DnKDAahgucMkmjG+CJ/ksRuDTWN5G1QK/2HblecOodtb4a0s9WMA41qZrRZ
ADEm45YvGUG3+mJZosn/EXOSLK8F32x8xcepf6fyap/JC6dWeaVBfDmRfCu97+FgXfewi0cL+pJv
hVgJ95lShr+L+0Eg8DZcqbdyvT1hRPyh1GwDCdvwMSRWjLSiUNwovFxcs4B3rIaUXGMHLl2rRGsA
cOHtfih5GljYfoa+b8FlWgJhfuNugyU+w5SpkZUI52k1xNoBiTvLDVAnv7rn5BztTUuyKw2iy71U
YOwZ0lWGvLb6rnC0V8bKdVOCuGpkstweDtB19aMCXIC248mYVUBkKm9kcHy0SnfYxHpeW+5WH/CH
RuPRcX58Xx4T5G4jHdfJg3ts3qGDp1Yw1fCuIlMmslM+7w+X05UIuIaFShD9bQPMgTss5TAMMqdN
la8viN6tFuLzE3WaoUuH10Mwm7kY8S7vXcHEbd76SKWKPvNZv3+d9Fzu2YgAUcIwgod1tABxcZ++
6OSV/wr4g21dODRPraHQgUhGG3ZQWEjhPgMBChdSGlR0yo1r097QXZwe1Gm6kvPxyLqzDdoc/bMH
/Beh4VoFIUGDtfePbv46l2i1Zqm1tj0HbWxl570MvoEOKWE9EoVhv9AV4+XC01Bxd8IuZJ7bftz6
lX1QThjBy8vGfALZpCLwrrzmpqpvBwssjWlG5dGCIzoCRJ/iDJwkjO7b7k9Ghizrc8K7sReu239I
4zXyAXRqNMjcgs9WewpRs2747ftDB+QRHIyGH2S1kIUvBcLHGcQBEKraKTNR0x/0CVgn6W6PciGx
4OEZ4an/Yj0eB1WBzJb/Y2Z9lZ+l9UQF60P23ylIwQM00SwssdoqxRIZSGc2EEhoC1k/FShp68yU
BfuaGU9Eid8QJo7Le1cw1xAYf4b+/wnKWJrl5rExqZQjNUcVgmvjCdnN2etrlXcir1mCAyknoBKV
F0+VbncXUrllkLjWCzs6F7Zor5mCBothpdg+4S7D0eW8jnTe3JMEsJUFrxXxyaoJ6PVKwZKV+Klt
5k7L5RDTTo/3AQpjW2CvDEjexyI+tyNASIK0DJctoKtS+gWeVDUKicubYlm/SUhHq2TX1O+aZxNQ
uRlxD1MFkXRxYgBkUrYiI8IyyTWcTFiZhSsBQfj79jIKgpXLOQS2WjpYoV7/qWWT22cRPsPT8PjA
VGX2bp3lFG18bNUgzc47lEPSMJL9SE55PgxADul+SX2u+gHr8Zn4DG/HMSeBRGKZ9zNoUb0vOGPs
MEYS+mqrf5WQSb/Zb31Ak0ZBNRq/7YS8zw9bO4LxB+Nv9/MjlpfV/2+NZDrIaeOLWdINPOuIpakV
kKwReU5Bb2bbtp5qigH4RzqKga49LbHTDbZDc7nvz5mhKV16qjqhuNxv8YAGmiw7C5/j8EIyjexK
lp3UAHKu4nfSgwbEMVmlZWa4Ybw64urWuHOKMMwq8Nd4RvflnUQNQKtc6U0xkruSVXRNS5huIHDc
jCmuL66mLdttZfEu76ohKYt/YfJsS7kE+cOUURxC00Irts66H58wPV5ri70q+Y4EUtjF4BmqrL2q
WJVo4OFCsecL7DWZj+9emstp/PP/xWvnrWCEfdCyCgLhIOMOfJb/MIlfWOeXxtU5kZDMt7PuZm8c
TBJD1L5Fup3q92iZGhbo29O67pya75X3/ZAFyK1Iv+CHLjJQv0YWzPMlo6ET3OU4hBKclSt5XabQ
uIgGZ0uLdBmsnsz3fRa9rRhNUvrF/dD6HCM/BDPUYKzElQsKX1fElXtSQN47IYjDF+W133LmTm8k
o3jqHEIV3EYJLlO3T5n2iXjUXOMQTQlvJpX75BIZvDrvDcTYRkU96wkH5IZPDNnR95P62+MQN35H
Ku0A0r1UuK3iJAePuj8v38oZwS3hr2MLoEZ9bPkTz0VsI92xCGOXFJbIHBG+8z/UafNN8dRsZRnv
qPJfr4ksKWPaOnPQpRMBZJ6REvfjUaeeLAytXkZ/0BsXVvSpp/nwsoDJ7STIGWQuNs/1Q7jHfdup
YYDeWYPT6kBcGXPcd6bz1bzH94jFFKlzgBG9TcXozgCX5oF6HBgMgy8vp2VhNutRukWIYoOuCfzd
8oW1B9OVucRI7R7UzmV6J/G59r8xT5sttu/Du2dEym3HdVpfwzDFIK9RvVRcMCdjCm30uqEnn4ki
I+XzSh0+We13WyRjP4K4MvNnXidUNdGb4fAX69B80W7cb81W++bOlvvq2MZafps7zNF7yVq86Tyt
90BQ8EY3CnFBImBuy9/wwfOpOGlntFvbyf5ByAH8lTEFzc/DhSBz2sk03l4BiosqIY63gCXSegkV
jNGeUnLMQHYx8jgsRV28YSdGtRDGqYnP7m8MfWr+ZmmgGxPhutD5JVjY6VvTg9lr8r+zwjF25hv9
2QeJTyUutCoY/4gA0Lgjl0YnaF6o4L0Mt/Zk69ZCsG8nBl83KqCCi9Xrf+PD9W/GqrrhWMnoGNYz
HyOuE2ZZ4DBRdBbzCwfx9B4UBorSS5oGsVXMoaCjXQaFdZU1p4JaVGevzKakridCFCLJTI1CQECY
K3NB/N5rCZQnz4ldP5zUFPRUd7w6z3aFEV/EPuHqGP2RihhNF07wAOvfJhj1mWwl9j/aGrnb0+0X
pwVrCoeyu/FpfNWrpP6Nkun8Cs/ecBznMXmqh/CvZ8d2z1cY+Mnet8ECmL9wksWd+VNzovoWQTTU
wi1MIbsLu6AJ1qULUQXdN6oxvAVARKmVloGqhsMBIqyGUtKlmJxARqeck3JTbetOkUXOi/VRcaqx
zvPDuJyvVfzWM8gL1uRA4lQXepoml2Y+RDN6Aahr0RaqFRhdakvxSJ6PEGuJGUZFE9jOnp3wBDBT
iI8UU7d1bNgAnyOYufsqymkMvBKM2hLknXhyLr66w1QqB0tjhx70YCBWZwmLcHAi8xFrU3Ugk3zd
SlWY1vLT52oNmwi7b2DV8cqZPyV7oeuomrqanjl+p0j3WzIXWNJvRRa84jQL/8vNC9pWbM9KSyRk
Drggzmr3aF/Fupy+QzhMQaXkTxocmpuhIif3sQua747uIuSV39Ok/s9arr/siZUTyuBy13XsNYSU
tkTIIfGi9m0E7wthYN1OCVzQMeqO4AvySI+qkAuQtO1ZHdVEzUVuFwW72nXMcdWIi3B9TPBrc62C
gMBasL0AMwofFl12X2gWqSu8uzpJbvpsHryScMhDtZEfEFrXgWAAFk/7IsqlInRFB4zi1H06D0A9
9TTS1V9zD1WiGiZujN8HY4dQDbNGIJQqn/HxIzw+bjwFQDK1yHN2zbHbxvxpz0ETDSX+/c7itKNQ
e1KNgpEv7o/OBsnTxCcYtmzAcgksD1iFTAB9vx1pHOwQK/+RXZ+qiDm+A5YFYTDYUSqc4tAy7Ff8
dHfkG3WLu4idi61y6R67VLKTsVE74ICWiYRhZSIR66/eD894nrBs62SVwDb4wRQFWxa+KFprmnpR
dEHTmKRO5p2Ejbs7niirjnkePRH70tnKYmky9eZMnTmSEFdZZ0q1DcI4IIzKA/HH0fgFdNZkjUx0
BCfJymumFq4VaQOeTesvV0My7g/C5I1GNcIzVsvCFunwLyrUlIF1kr39lzD8rGyQXQoRDe3mFi1Q
EgyGwrIRubx7BCVV/xar8/sopflWf38YO/staFwRNGL+v/nmf6x6FxvxPxoRHQMLmFEBBqTFMPT2
C5UOF2eaQLvKtmRXz56tsbxFlF3A2lW6hIwmiRnsdK8TPqbPTrWVzaZ5+FIj6fdl5f4mbnmbs1dn
woN/oK2vsNsg6q+VIoem+nzrBhPu2O+GeONUpoaEFixpXN9cp2kGdqhsTkPS4ncD4qHDbmc2N7/D
5HTtouaVRpyWLvLpu2EIYqAyvvRPDBm92d0CaI3hhstdfAQA29SFW4QP7HGxDaXm7Sv1C2tVgy7R
I5kCAZCIz4ozVTExT8xb/Ul7veqrXuRLidMh6SeD/X9QKgS22LRI94ad+mEQyDikEEbGVSZPZFfr
fe1ci8n1azZk7j90iSKOUp7gNdiFIUvUb2MUZpkhm/DVWXT2hpqPIQMWPh5ecP42Jpy6wmDukrm/
dyRG15T9EQIcerYn0v/Mf/no5eLkkjoDNXkiOCJB2giKn/BZo9fKfGVhC7HWrms+uvYvpXcl8yXF
8nkk+1Q6gfgkwiXSdeiHe2Zjt8re6nBGN1JnhFOJHAPedyjB0tRG0ehHwnU+KSFGRTH7onxa4oBo
iZy7mpn4XivqCITRW1kM1LQz2QjY6D9J5jXolZApkgcpXQSmq6UqG/j+ACgeDRC2kIsnDrdiCG9C
DSxNRQUdtNy3EoqVXsVngmPgZcIlZOQbDgkDcuMPqaul5ymqFTKkZ2Y2JELJQAAOs9eOy14SOlpo
OeXKRvydBzKIWQ88896jA/yreF7AmmINRwGGOPG8hNE4vYnH/uNH5xvsN9bBUEgfGJfuKVX95Yz8
ERF1ReaHc5B+7dKVjAbxNvE9zK7689QbhhPxqbmeKSTwlsJIqzQ9A/K1zmVtIjlaSWeDU/w31cJP
Ubrm2zuA694f9b02+GpNKfAWIYTgGadV9XReYrk7fAYgfSGip+HXnuzOG2FDpNGituXppICi+oRp
TUMVnqs9JKMO2cABxSbGhUtJ7tP/jNeZdz1skLK2DneHIwbcers/9u9IURFjWzqJJNBwGw6Zbb7i
kvgOfl5+RKc3H9QQz4OBUkUAr+NlkI5Sd9WHM55j/f7dFP1h493Pfzru7s6mql+wWb7ka1RlH4Jb
+9x4P0049ZgfzP/tIT90n1fS1OzFrkahg843gGx2vPwSvIUg0NI3MviVhjmnbluKY0EChPZEO5gj
1KfCNWep2Mi+SjyRnLPklH5sdlJZhvZGYVUxXoSVrrw+k1XGfRp5YpC+uYBMz3ltnl7wLAvjPqf3
lVaAbaqu2PGiwYRUaeKuo95gPVGPlNuCQlhzprTf2LNwuPK094IQQPa35sQZdWZZoKzT4L2OU/UN
C43PgyNW9DHTNseW98l5Eyg0xxl26YDmSsPnr3omb7fu61/J1zxla7kZXcl2f4AtygbKEomc8jwu
VQL8mat1f0sxWm5uLtvsMFKIjt3jqNj3P24Ma0wwIqshOgA6d3ufZy1nwYtyXwhRj/+UXGxCa7NE
5iZCPN7NpBTIDbRJsUXoxoTjo9wMhNQ/jqOBkDI5GaxKZ1RnxJIOoPeDlpHPqALp2eYp4TYCkDq8
HfdXNi235/pnprRZVott2xMyaSFx5UaZ9HXctCS8BjNHWrbjQHh3lyPIDtZTTtfrYwNP2/YE4KAj
IurnLwQOaUuJCu7VFD1ELGFgT1GWEnSlE2RzxWtpCDC1Pzm34dNZb4TO0L7XaNRjqIPdmKDl92IW
SE5oln8fGJikhtx7gGW0VCdIdqUPe6att0tNmOuZo/dyUaxnV0P9GAZn5jOXHTDJtpk8udSTBtaM
EQmwdFzSspkPTFTkvHgC8LSIq5vVaKQfXrbBBgPPUtc0mgHIZzGPzYIqNmVGWSC2W9SFtXgSF1G6
Ec9j2uqT+Rtca4NMKq1PZyg/4O0esVpV+BNf89r/6n3vxea3L5mgWgwHVDHYSMfqAJPnvs114J8m
wXIa6990zpxrCsBQXE7E9VT+sKmtFxgTCuzG+TZ0B4eNd+roowSiBOVUa5UBHeNRwnec9AejsEJB
IsRmhNcAz72iqFNjHmJJIljeEfqqAIfuTg0QxmCfE5/hkEOmhkxyPfmwwlusvaVGGJ0pQt2shwgv
pRhjlgUi1TRA0Zk+ualzo0SEhKH8y6SGRTVtKuUza/p9carFS9MqC1EOHncdBf6ZupVanyLKs8va
Sx/jROdCw+3+zceD+w2icIT16IdxVb075qKEyIqEORUqcbz/GdPNQ1wOtiUpdMKr1Q2CjmO/EHlV
2cFy7YHvYu/8sk05tdimq+S8XHZ+9UPl6fT0/Yw7zh1kgH3N75KvEZY8uEkI9XOPTZpIVnPw/kjh
32xNB0jq+z3CVC7fd3ksj04IfFFz3fAGz0L2XxMXEKCpwy1mKrAQSZolHohCTjUPloXvXQ3BRmwe
L149LYGfibYx3eqhlGwFGod6BAYCBETtuO985h9etoYKiU1QJbidvBbXDszXYcmlhVdct6goGotr
mQphB9UiLHwLRavMCjt2bll1ytQzsiJnHsd0uX3JzKB1qCe3gCO7W46FeMhNxSKfoNsBiC78u02E
NV+8YG+VihTHafIYkORy2M0A2MZqCRrYqeflqU7qwsc5NSX/10alsgbpbJ5yigJHopNs3esTlhL6
SqcMqNC+VipFUtvWztyXA0dsfk3xCd8onZlVhox8efrB6QERleiKM/OgCjsvoiKVSkNFDdUWCTIw
oRlnS86dsZfVBCTl/nDNL2UzntdawiMpBi+rnbQyPMFAUbVSuPyO4i6kBdWBOQ+bhkEBSiKP/qhb
Wh6RiNLBNgmYK4pjCqnz2l3el6U0SNd3YWjkU0GhVHI/Zm2FXVklOttTKw0/AlMK0UqvC7p/nngp
sCM+ttHBGwwO3wkPEAllyHggKqhUes0n61Vu3eBsKhfoSS9rcq3Zo2wM1f/1OW8SX2t+yRtGonZU
/+6pqUhQQPw90q52T4qwRcN0aihEQ/o8/DNoxr9BgbUDIzS0qsy7tEWSn+AZ844F96byLeeZ2kGe
aB/JI7IUWVsftGIs8z4P/8XqVy9WaH725UMmJ2m+382s80632WwTZptYJINbMAsEnG2feGqUFvcM
rvAeBVMN7tFnYn4ZDyrZxYgpQgt//02iOd/iWyq/HUvqA5NdhP64j63OTh54VK4G1PSrQX1wDPTZ
AkELIyUgUa6IgCdGxA/zSuK82a/2KzaKYQfBY4oMBQSHGvzLDhYJO9a3CV8YXmMBhQiGruR3fNTK
273hVDjIDcNRK4yjX/+Db9goTzoZESuL05QNuvD6t3Bk16mtrBErVEt3wjEgoaScd+fqvYOkmaGd
xumgWD9WVTJQVQqjRfSFkDxRU5Jjfj+2Qz20PTCJ96GSoxMpilIo/RH+lhihT67/5DZJUDL6jDrC
xYig1yOW9q8CUkIMlrJSWrjxge2MHj1KBVj+l8MUQM2v8zlHVr4zo6mH8AwVwsGt5N8JJUe+CAfd
/vG38ZZlTGpyl04czNyvh51mg/zwM1CX5X2Q01je/aJUdsXlr8URt11fspJkAad/kqEjTjssPj9S
Q8TXKu3O2Rm8MYi5Vs5+jvGu5DagPmAautcqX23z6quWBdwOMkIRj9prfVzLzL2SyToZRK9uXqdZ
pYfTdn+axmkCZ8PvhXdScNP3hWrFwNGNg8YFulnNrPbLnS2cHf3T6SinPlCmheE9LgzaNq+Q0hnW
VqQRq4a+PKejSJQxrFgoZziiVnoXlTBuC6L7aOVVBU77KCIOYbzF2fgLlpilCQ1yTnJslUI6xirU
y8FzDA+rQOgzYsqgOb0pFHCImlkZN/u9Nmnqv/wynHM//CXd3KrYskPdmpCjG2JPD1sVciBqCoEg
fl+9Rduw8AboW8eeJzAW2affxj+bsTtX7BnMf1ByFscQIYeZHEDklpFNtNZzykYwfyL5mDU/1jKT
cYGdaWfKnCIjkMbcJq7GPnH18oHxCTvpRFT4ycClkN5e1Aq25e3daHvayPphblP05tHOqEEO8Tg6
XjJNEvfDGofYl+2d087W+AL3BMgNhZY4c8os+3wvlvfmg5HgUucUrHgDX0AE7BoG7OXv3yTP10Wp
i8mTxLmbeVrloKnqGDkum4FOWovW93GqZJT+rqwR6wHOxIzIThwfW0L0+nrcA1QiiS6AV/UTe/8k
xhusZGbm2uoQ85fh/v5x6BoL91HdqfU+EYDH8wB+zroi9dVUOgiSNHmJ9x/rASnZ3PCo8FAzmw0O
gU9fJ8IXs43uWouSEPTFB5JHOV60ImhizGMS0O0C9q1y2fdS+cn+X8rRP+/yH0X+fbhf8CPdTTsT
Y0Znz6a5+9o6HrnsAsS0UnAmHVankAImeNiLiHwWXvRmrI4g8DmP5TgHUEFHW4GlGz7WWO272Xcr
lF54VIKIOlVylh8LaiPY45akUoad594Xn5UnahazyNmzQD5qPQ8ICmXVu5/8hgicVgwWaW59LWIo
UyBhhtDQ/u2NrnNtoVBDtuuEok2g3AyNX9hsdlFE75bqMkhpkH61Cs/TsW+rFLtAJilcuNCrdnxE
p5ubHGoiF4VSC4BLTft87TuLlYzOuHeRnRAyWFlDAVXXv7TypYSjTkhuG6UgNged2sSmwjA2XJ7a
trPReJwImTKCDntTLMy6lIQgTMrxQywTCFNYINnS8ooZnx9uQmAgillR5r8KHUaVgJkS+pGOEXVL
gpZ6AGWY5kYJKmAkNPoLgh9gBxHNYEJKzIEFxcyBaNsKhzZuWtIrrDXTWHdQWMZzUxD/ogOLi5vJ
FFik838JLkltckn1QzvxzOixzVyAa4VaVxX0qrPArLmhcDAmRUYyYBqkej4bkAzFDu1+gcvLGVOb
QiIMksN2NAfqqECVE4OCcAvMkmNqYUCKFIwQvOJpBc0nXxDvewTEGOUti5phfsK7HAn7nB4pkeun
h8RYU5zexHPPQcu/pHz2Ozq2q17BnO9BXujylfMKUKDn4PU4wPm4RH3nP9IjLV/eCSL6Cn8tNhmP
fzzZpCHjb6S4byxE5fQgpR3o9x68aJX1XAZRXo9DK1VodANEFBp2PGtKjC5hoSxBE7pP8QTnoPMn
D35HQpyas08/xyITBNuc0XUcfae2Mr7gwLJyaKNEzdz3hzYu3+sYvyfn7t51OEuYc/vcmikNleGa
FD18MKL6tEzsKIMK3JLnH/cIdhUiVaU+xNy076cikaGDehCvaY/8YVzl01Q9Yc5a/fqyyMtUaIoO
uiBYZj1nUiJKzyRnur4h713+1rMDi9kN9x4rhIKjz1AYEhbdhCf7i/u/mydIgqf+9HWtxBPi4ig3
t5/5yO9iIzU41zHBayZrcHidBquUEf78E9Khsb4/Z3xfxJNgvghKCzeCOEFUPWFeRMRhdzw7ls/r
zx2wUu3XjKBpdkFhbLrt8HMU2q1WUgEwr1W4gee6cSj9hb+tNelUV9Rm96M0RtzWkaaDdjIOO9J7
z9EkzhR8oRwcxwam+eKuww7VVBOmuldmNWcNYo29vJtDMcsIw3wocXOIwq7OKjwMdWerQeCvPUze
4U8Lqu1I6ho9WLxEhfnoDyjW6AwD+xoWgOFuaBksFHNUNFiADJQLMDQjfq51llyICqJBKBq3Dz3P
uQVFBz01wLohHqJEe7J2xmu1R7ts/IIj32vNnhWMc8Bd5DlV6/Vt57kyjrNG2nu6BNQ4ycn8fI+S
DWz8Wu4viQEJMZAS4dXTFhMuybcqxL9QmR1J9+t88n41Fd6yxSDoLxDwd/NdFQwlWcl4dU0cPZgg
nGBRtw71xwc1vknb8jH6kM1zvOffn3Ivlz3/lwu0X6Pjxnqn3S4WXtdPL+NCwioyWFWGy2kGDQ24
1q3cOoUF4ldC2YRPOJmTjIRAz3OpmxCiu/MQTg1xs3Z3jMEOqkoRvSL7H4wRckkoJpPJE7wjkatw
IQBf5BkqPBEqLoVaSOk5ABNxUUyb8it7JgO/tYFGM86KmNzGH036zC7h1NOdD2KZXJrDtpl+4lqc
g9oFN4My90ja62gU2VzRe5g+ij5bCBDLczXvz+NOf3yg2rtVD739IMxLx7KLEpgeGSPCzXv1OJ5O
onyXt/y3j4MvgMHgGaqod41HI4YPSanP53vEOMebgxmSYdKr1ittcH38DOFGBIe++Wly2PDcuCgv
TO29F3BVb/BNQ5eNOCHIRsaj/xAgHOAIIIgQD0la7SfqLOn1ifY0K3m56OZTutpTUdukew89cBeO
KzZHQp6wS5gZshBqbF3D6QlXOEtqxNHa19TvaplzELkcAlBcQNT/j9nBGMxmhZQa6ioViUaAGwTm
1pOIn9QmYT5lkMEkvqvwgpAjjwPhuBCUoMDnjgAs10+ARbj9BCTzXQM4uFaSfweUJF5G5HjI7GDh
MQu3cWvrU2GLJhz2PnGalWrt/i0ZsSbMYYUennLNtOBoRkvL03lTWJ0wd1UglEA6q/MxnV/lbzKA
hq8ali0RfDyWID1wZlgA3dCVLdC3DiWx4CXbmtsPNeC34Vk3G0HkD3JOva63ypXBXZmYUDHIAv7N
VX7UOTZ7fU32/NPcoUCn0mVOod+I7/cNnV9ayZ0z6t5qMei3P5utD6FuMXtkxsenz/BFlUZTal3T
lctSXsIly0ftkQlrq98pNQvGJ3zkcxJwISkOHPTPPx+t/YIKcvf8rEjRdfKVqSYIm07vPQZMol1a
ozybr4ZHeZGQyuZ/WuxcrV9GBQwtsqc7zwcKpK43YlyMUoeHUgpXcH73OEyOExOzTxDCeAvqw9ex
ypIFTLGwl9Pedd29peuuhUOuX3nHuWlbuFeCtKZ7S8/yDUqBqx6oG808vhigaUD2Kd3P+DJn1lL8
vN7sBBsIk0Wb9SOoxgxNWp4lFVuqo7RHBnNawh0BkKdcJYQAOvNRIZvrR2XYefTs/+VEt5BtrmV7
wKEEfnK5MvViLGWCAi/Sn4qKdi/4ZEMD/gzBwp/a094kb07IfDa9i7c6xA6GEiUvwilYuBxLnEQu
rBXX8Z6iiFH2YT1/KMZNW/8QhJH7KB/MbwdpBJNiof6uiMg+3bhy30XMMFAMHBvjKmzxCNOTb5sJ
Ehpq+DkJmF/pzkmj+QGTsXmjE4IkBCLcNVtlTWw2UvlJdL9wUu4a4rCmKRBfdyUzpY+hJgBsr+zw
xQ9r41qcyQ4Pl5jOo/w8+RVP5O1RBHiyqsHgk7dbeTBHawqfDbItBFsBjkzn0TFooyNnRbamBecH
wrVEnW/40r9mmomYj4AAa2Tnm7wOSP5IiY7j0v2AdgcDzLSqzP1uV/5fuAggGlzqEiPbJUruCVu8
UqbGxgk8btMSRccGvnRQfI85SvQ8hnvGCzCMRjW97TYQWYqmsSbvVwuBrwlcvc8b4ZRIqqpumqN+
Q+6y0J+HJvQFXZEAWHWx7GwA+PBAAwAQumD7mtYj0iV+rZ+M41rOSDxIhY4WKxMn4YABIPJ2/syx
GgLGlwo7dixTMDQg173c9yKF9mZ6Oz2rxpWdIZEWWYmQlfpJbDBhtudPQOzLBRH4NqrwcBoqmXsg
Dg7Q5uyoz+dW3PKCHe/qQNfWip9ITGcKXXsFmuCXhDlplqSjcGXnGql/It3+55IOZalU11DNQmjZ
9UZ0JF10ENoJHSFCszugTg+TfgHAiWP2B5mmyhfJ4WC3ocHTuF+xINeXweezRD0+HlVyJDgFOsQ+
q2Wc2w9OFc24DWG9q2ekmIZoeDQ2jR6AKLvcOhRuEv/0kOh80vYpj7XGeoqM+bRmvJEGkRdP0ZA8
Tpk3SNPZ5Eb/opp9drq9NCSDrej6UJlSw87q74uMZHZzgQdgLxFQrEwriDgwhNYAjxcd+V3y78eW
xr0ibOQXqoQvUd1vRSrlEBEP2Gg2GBFnfWuNrVe42/Wkr9Cp+/e/Uybnh80kX4LSIbGt0HeoouoN
HuZ8WL+88RWzc4dCKiLFXVh7Tdtkcy5fPmemHdfwzLi5UBwZmdotyikJ9uxohBAuV0S7w4oqOj4j
FQMVHpfR55yM59fe8QZk0anb6O3Xy9OC7nPR2sY5XTWYXZvKnaNFE6Z7coS41xUxBkXxjo7aoaEV
9ZBB7WyMOdl1LbW6IjJPA2iN8RRm+nshLMdko9osr+vPM8EV+uFod+w9/skITgeorIoayqhDqoYW
Rpodjr7N+gLcFTbz0KlLNobijwjPTsKpuzQ2B3PqZvY8UO2Y4/Pz28eLFQFIBKSElckZ3uvmcNWy
i0Rl2eKI2ZwH3OClfzdv6a/F1Kclz3+njBl4OdeWhiG79crsNiBEY4l0D+Jf8KtBMIwyl8dp8Mpj
wzk44e0Kz8y9n5xptdq7r8SKuQKdmA0M/pMFBj1E9lj0TE+Z6v9omRKixtpWW4UcihrPvbxeRtjg
Kk1L2da6SRv1ajSAIwXq37b5IAvLxfVfSsLo1wlh99gItZV7HgA7+eEieQYLv9zzPJek9fgVqFzi
R51gQJNTaxqqqANbNNLknoDRKyywrCVPdWxcCKsCi4I0ivCbk8uZFFKRW/BhE4wjZ6yMhK+Qlnrt
Wo5xblCsYTeDwdDIJTE49uhmxohUjbb8PE8FvAz0LbVWr7do+5ygBOAxFJWYlJUBBLX23oYuj1ze
oasBO0sdvafrOssmyNbeFB/G9jJl+pNL0n/sGg4K8WMD7JdAesfsmqLsyjFGSdElAYxeHSMMLvyO
BZEUR2gFF4FlINAYAT8DFkeFIJAtl5jEsZUkww+8biiyEfjwoIoCe47MX/mi9TPcTOa6mdCB7WGK
SEYdeci3P89j1+V3OAxgMRhnZ50IsuZ6ZqnYX1iTn/WLNj5/bqalQM8GHszGvt/h0QMo2cPjNglw
BO7RNvb5RlZBsBssp95PKPRFgInILiJmSJgSo5rt/jiitAGvaxku0mBrHJuLb8WE6IvqD+iUurFh
iV+Ifo9qgkAOzF2n41OapS8So2EPsia4lBW7x3E0vXXJDrUdXs1GySqZjlJ4pmYA6gYCg3CiVHtx
IPz+WCG6JwAF5Hu2BIoG33i/ionRxKFBsmA0Hl7P99QiRZ+AlFk3q7omTN5VzYSsuZcApLpZbG+I
2W3BEGzF7J2BDGYVDfMm/kgPtrXotRZ8DJCNJXf8iYhsyDpF5TyGyAl+o/rKFOJJ4RIyy3SzL0qV
fty3+n4wC6TxyyVpZoJrKO1ekF9QJEKOe+0TAHQLMDbyWW1/tN9+wASV/4Ul1zHa0n634cUQGDx0
jNdOYwuHOQA215zQY/RofuF0YrJoAqtcXyWghGjiXB3fLB+KDC1VJhITV0uZhu+l3a9SygPgm1ub
AY9GCOtLC3aCaECfbNwQVfGN1JRKn9f7je5Ax+WDnpUdFWZp/Xu2AOtE0X1Wj8QYz+8rb6QKGoC+
p8evnRoOSbs+Vj+xAmavsRfT16JLJOgXTawQw1g025jfq/U/+Bvk7J0Z+FxBk6SfTd56EezD7g0z
p/6qzGZdnDKsNMX81WnCXi13n8WvY3FYMpXtd1R789eipnXGELOchhLJF5jIJwDRRubSZYjL80wI
+l2G3ip9ncB3fakZCP5Jjm8dm3YMd5pi9M5KPGiUhiHnMGUny34LVctw0m2Ottku58omvtsfucg7
6EDx6rvQDTYo1JtMWjXvKcl4OfN8d0ytUYuBZTq3tQggeop8QXu0ESpgEvX1Vy+PZrfuAH1LXYaM
om9TJPWNQI1UMUO9L1+vInm/emkUjerVFJnTgocR2tDkfruMQDFMnhgc5u9s4aMnlV9DgpkZZOH1
cX1yPNe5bf84khLfS33vrW609gOD9xBy9JwUGytJ0tOUz/jVgXk1NFW8IkGKTLmSqVirjUT25Cxt
+XW2E7SU3gICJlKKKuPENLt7thD1agtisBw5H9K5bwIzVRAwBirr1alwoO4IsMS9yNidr0mKIa3f
tsdZOVzAVSI7GVlMXFp9XaheC/4B2AXX+6Gk44OZ906z3UgpCBFvkEIASKW2u/r12PxweindT3P3
RTZ60Cg+jWbGG4D+7WZC+Rj8AjVFMRaDQDTIyOMO2OC+umY0+aUe9cZgXf6YQduT7B0H7iHK79bM
/J0I2q3bStAD2At/3MkV+MVSsMgC16nsLF8PbBGoVhFw7FHfkwZkCsDHvLtwGqAxNzRObemaI64b
TDZaLeP6q89bAe6N5C7f7AGo0cmeqQfbedriwLm591150rZbI5TJquvhSB7Xu8YSXniHGIjhiwzJ
KNmyzS9wfyT8IgyEYSzjoVUP0KR2JQo5XSFqu2+S0KE0jZuc5P+l7wDuI3H1kZM57SHd1Zlfx+qU
f25HAe9ABzMJ6e5mTkBowts6FIkC1qp9yln7rLSSGun+Ev1BeO+bSSxjw1R71Gc4hAsZA8xPYKe2
DuU5prA+iJpt9PrIpsN11Zy0Zy6xLJ71v3CO0iAaDjatjfs5yqvMX32wsCMzwh/si1O3dp469S2i
XqMEXOZW+SOkvERFpqtbDqmFT7wFMrVsLhzuvOoOYV7URYlfphXlPgrWHQzKqbvEpxJnFgxN2pmi
WJGZ3uvKVvunJYPFf8c5zH6w8w+B05zCgxRTwuCwNrES9H5Lb7gPnSmZc5EdLFCfw6kvqBwyITxO
CpsKo+o0mFOi1zyVObDRUkypjR2Y1hY7THPTV0lyins8r5ofvbxqjqpDyGIxXqQ0m4fjgoXIO+mv
R5cHlsBlJ0u+KwGYtfsLeSvuVD12m00skrrtSbcVIw0pP7VzYGqRGV+5xDDeMFUdAZpw3XjRtT25
NR6mUvEC/1Fyw6VKx4F+JCRN1MpaVkkKdPe1g4ta2Us6/oEIIHaHhAJAsJ+7Z36Nlj37hvYJ4aGN
wDBr1pPonHw8asYwQWmFb0LExX/j7MnaTAZAl2LsbCSA1R7iB7x7xDmBfWwp6GX1Q7hWPJrYW6pG
Mj/X3l6dvTfGvcrbrhAB/Bs8XaIwj88Em/QTkgDwwY7p6XwyaMUkJQpHJx25QCOOSp8muoLV7XWS
TFW3tQbrtmtcZygKFhDfsizCt+yzU5Lijk25tqCrTr61oq55T5y7mqsU4jjpkofTtqrSQqjhXw2/
r2ssrwT9xT4mNs4xEDWBmwl92h7V/4A3XkyjflvLF2GS6nqLH0VUnHAQAv7mRbCCZL3+YgDQ2OmA
BJCSLsWhS0glTzCrEtGUTbKS0J6IHOHMAgfPX+J2BKKUkKre1I+1ppzhme/oyrTBjbwTmgLlZmET
6c8KX2vKmKEwnYhiKGfJhZvjAVGge1nvdhUXPCfVSQtQNI70ryAUx6B8YDFNlsCk+lFALCg7U5/2
BI//KacD6DpY7eqmP0RBXMDaGFrrZCqLYafdVNv6dViReiVHYMiFwPx4jDNRq1Rn4hJ2bPiWPJpP
n6dQ0XaR9ugF0mrS2wrRTEm2j70KVyzBRc1UTfMIoe67BuifE8uzKckz8y2smjA4UQAIrP4TlZ4Y
0LwQ1hOZ+ndSmwZTPzLLid5KE5IybLN+WVKbwvWo7m3Ewi7It/gTdh5zdGVjfRHdFIOTcmibe7YE
PjhuTW1em5vlP6f0Ty4HilETdNXzPNGdJOdfs4MeydLnxn19hir9tsuekIY35XBfC9FEPjPTChgH
O4Th9nRJEsKuGUJ+eDxJ8fVa82np/K2x+Dxdn9CdKXDuP+JSsf+73leXuixzG6kFKqhqTBuWnmgB
aWdN873/c/lwGvZjcw5hbQlFgTckjA030sB0lXVGhyFDQpys0lxwYlU5LQI+f8lJPoVwB69gHUEN
WU+6YtkCjdzrtjfdNOibEELGBd7030+L8kx/8TY+P8WlUEyGPAynkA0bp1iVZeN90KFGzLQbNILj
CW31Li8oIWx9CMdTT62u7ysIedOuzkZmxlFtThxM4su3V9eZ8HBp872dQkDMZIPHo7muQ8GeJRoV
u6gqw2K/0PofAFFS2yRGqe0cQ6JfKx1vpNkyXU/yVZ1++6g8iDCyzmbwEkA3JuEo4/TnLVWJotsJ
kZG0ND2AKg9+uqOsYO3C+XgOHCbGCeHUgZqGBtPFtivaCgjDnPDJ63vMGOGib+RjwMNHyVVe2s8z
7LDQxN6UuEIcYBAuWIajupLdcLKzto7IZdrKhlTGKJBKKw2OFA2H5isItUJ66tDvuVavap73Qpvs
tCmIr0iVgKpKbOxpiAUIIR/mtCXdFaMhTCwytVv9qO+SBPsCsWGa9Vm0UYqWx3BZrxKbOrNet1Hs
DZJ7HD4DRKjF6wB+mB/bsYvnp/f7/6huJ6FmhKAUkb8Kz69W/jenkMkE7PKcIIQw4gxeZ+pS29XZ
wGpR49o3oLngFGVboR40njL8mshf8XkuiGpoaVMUSCMcsP1n0BAZxMzOIuxOEOZS+BvSdoogeKqW
E0N4d4VshvSmP62RoCV1e3RlBWcShCpDVvFM5g0lWBy5tyQkDBY0bzvyuGaYh/aIF537zRAAJyX2
3a9tCjVTB+4RsxVkomRqnUYwsPvmWEKmWRAq8rWf46YE0jRGPskAr526fyQmkONJeNH7xNqNFzr5
pULhfH1evCg2vB1SOUtB2nDndsH9Zx8pYUb8Ny02AwbhijSmPyPlYU98drKGV/TMXODKgTRA/3tl
isGhY7jJo537qiZgF9jn1xRs2e/DSn6YalnbhajqSIxOEMZ0Ji4d+oyvLLS+DianGsLs8b2brmXT
UheFhifGdfPBdmwS7pCTcu2f6sv7rWHgWFw/I4mpaU3DueoL9kfSazrTY6p3iGjVJ7Fg8KZ1Lnyr
LIFV9VKbS0TJzFsY71QVOWmrdBVzJr+D+01LH21kqR/pzOFHeFZ3wuGuvmQsF8xBDSSx9jlGGjY7
kdRORRWPJLdA7RXxXchLO7t0XFOhHEsIdTOHbOFLcV1pZ/0G11UYqz7guDDM+9ZNvj0kaenO2Zqy
GVsDA+8pJd3ydn41UV3vvrcMZ1akYnLsuxGXX9rkq5lMlIjCqIIGCIvPt7o20z4B46dyvDyfffPM
BwT5atQ8yOR8O5GXWfqvmNfWvP2cICAVnOeqrparpmiPdl2HdyJtieVywTF6wmkeXCyuYXKH9XYe
8GCKVtw5YDaElXeQSQE0abtKEeodgViReF26uHtfSvr8xthoSL9vEcNzaseu/xknlW7QG1Cnylsl
V2hsZPvBK5smofOdgkBp16Xn/+1nrB+LtYol+bcyo4qmFk2cQMZKw03SB5GjCvTIku7BeWqgh7f9
8UeuxbXCi5Q+tZSBfIkx6Mt46AI0jTZsjD2JfeLPW+FwFOWLkMSEsQnzFS4lIwRj3qMyV1fJkW5d
bprTufWTVqMebaSgupN5iREyn6li6Hmooq07HQtA0P4Hw5OKpCuBKcMCUgQ3jjMKxq8BDWEYd2eO
82gzLDoGb3kdxcK2aCxs1VUzkrOv78L/en1fA+8eXJ+XtQ8CJPMVcBYp3yC/CK1HUOR+WJGKK0cZ
7z1OnnrTVdLAbjoxvDdYOhGMNkjO/X6k/5SpzdvNSUX5ueg8WrgZwmKbgGAQIdrRxGUHwpStDJfr
kXZdn174mowh5fH6fiq8Ga5Iy+deZuNyx/Ij32Ww3ZY7NLmmpxDLRp7Zmq012yPDMKwQ6Wshrgr/
L3dNiDQ24AfsLbZtxkxb2n2VG8d1GccezRZHh6giLu34n0o8olwuY4iw9EyQOvixpZEEB0ryot84
berMavrRkCvm0vmUXAz8vi9SnOKizF77v1eWq5KPMXYjnVC35T56QYMGkwtmEEd6rI5mM3gRUtoH
nkOoDs+KKx1C229M+jR8CLP4A56u3P0QZGmlrIYygxc20GtjjYAvajTU2RH3DCVHeFaSGXt/XczN
+6xHQ7ateN/P3Hh///HLnlAenk33H4O5PrxjsIUV7yHN9gsUvQlyjEXeHwvIErUK1WrSsysQhzv6
khkuntJfb8Bu5iA6feotsvVuWk3KOxDI8HoRsW3J0a2LYEbVmOmHyuT183XmdHhSwjl4F79LeK7P
TWjI4TKREVY1gfabAN5VG9rtla6KZMN3SLz4ufgOUHyYFZEaDEkkLz9HZQg46fnULRcKp0xtF6xS
IGrgBktTJdr4X/GxDYWwCy2jKz7m2419x9tKAx/rH16SjveW/9pSg+GudluTbOnPmgijtl/5mKMI
57YS9GKrrxvtmVBjlxlmHn7iMvZ8uXwBmSqPmnh6QxhnJaCDy3IGpOEIQ9YRhHR5CyxgnjikYgHk
F5huZdqVf7yoBwEZ5CXUco763kYLe2G0xt680e55Rr2rVl4Wxr7e/lEMr+Kac6kBVyZ3rXOKlu8Q
SHz93xmC+QIuPmSGmLo/Y6H4TGcM8Tq8yRtr5TILCu1yE1yYg3K5F2tNjZrzbTBWBViMddnddO6v
mfFBl/OAffVs2YIkBQcCan5lX24dPoWQApGst3kAaW9imvzshGSva+2liMC499vuADOssjjSJhKU
C9yefDk8QhZRATzCiVveUTmwTNfec19eI29nkbC5tpHATiwwHD2C9JxMg9ICKmYtk50CZEOeQWwo
i//B82Vd90mk3rdOsyFPR5zC4gHeW4vLZzh4wgpa8C3+JSJX80SfYQWcrJJqhsHkWkNojFmpgJib
SAL4fcfD7wOUWZSgGqDKfh9iqsYFzfGykpbGzebp1eE3CJPno25Noxgje3dkkyWQbp0pLCXh9Ywa
tPDgJMexE14Vg+iw8qP0MZon+J/U2EOvRH14rVl068AOewK6LKKVyVXKt6evRfXyK4cqY2Wad6e8
jwNaynxE3nOnJR6qGjZrpow7+MLEa9jp5jazsOjreR8t/ABc0fP/PNqha3yfGW/I0Y1p+JW8E/Rm
VBUrOQSUFkZh7bcVqCOPdSo8IIGgqj6feyRxxOJy6Xy6c9VAbMjnlSZL4BHPj1A1l5GyN05wWpTr
ypnFyh1VnvUm26tQd9zoH/YRCFDT/N5g/AUmcyEM5LNqRtbUfZP/ZdN+wlxkZgxSD8p7Q2Kr16pc
5l14tuVMWecHdSKK3kVZkdq+1JfGNSGaTeWUMkD4XRD8JKa+pINXV77Edit6N1zOftWpoiyCRTbZ
sffri/PS62Snk76M3Bgn+krFOJ1aisXcCYrrEdH/3UUeKKfKF8RTjY9eM9PHRGwEPfRZIIGq0BxT
0vDk+rPKhq1aKKWHTlQ8FvC+BK9I3nhRa0JI5iFYo+5Lpj0DaLU3xIa7uAHa/SVPCaARuqGTm01k
3ntFqx4gl/qAQ5lAm1MgRROXT9CpKUIGfRzkVTR5yxVaNR7lkfNbjXFXu3UnbZ9msTFOh9JlwtjC
/y/K8hbRT6K8XaWvgjJxqF6TBnxnOpnMFFWiQj3cGKFJWTHi6h8HZkXpEPN1rhJibkcuR0VN5vWN
53ZNGoRQt9E3E0x6yzZHEWxIPbrQgkYSwWeABMPfNQbEEG3+DryU+DHFfTBjux9nKZoJSz22HCIV
ZfjS4Mghco80O3JQPpohEmLI2IOEX1b90er+kHt+jtV/UbT0sRYN+54Hezy6/M9bbA/l6Fos+UA2
UGEHMnMoL270l2i0riYPwlFBpW0rJ/xxBKzdzmGxFtYzJDGRYhnNic4oBOdDmqWQ//d+lhiXMklm
Zb2XeGOOZUUUBjs82v4E1qzs0fw/0jLhpbB2oIeWraRrwRDUga+u7Jlomg50wqK02XTpfzuu7+A1
bPFhStp1b9gk60f8ogyYH8ZpI+vC7j62izzVEyvbLjkhjS/w/S8H2eZB7bTY6Z9SeR5Bke0jmPL8
Z7Th5KMnI4c/pOT3OgqYYThHZOWHRyFbVwIVSQNkLeWMhToI7/hfp4GAJkW+iqqMoahUIEIDf11Y
Q6NbtBBznwvyuTt9SPnsL8dgaSdDBGCIPxeuTpdEmf23oV5uHtHvZK1T2FnKfrqLOSzkWu8JJsXR
kxP/zhAjcsdyASagRBXwpIbnrnptJd9Q59EGF34iz2bqyKegH5Qh27+oedgHKLIunzl17RMyZFfl
kTdDxR/itpzn3q4AlUqF+gniJ6BtxDIWWUm1GBtBfMfXqv6S3SwUeTA3mXwJRhq69En9a6MNm4V9
FPk+hXv1hqOaG0O7Wq6vqjGfzou3Vkic1MaAbkhDyRuI1EZ4lILnVLZCIW2/Elj70X55ixc7BY49
Ek/sIVWE3+xEUblhy5rOCxg9uUN8h3LwbTKDQElY/SonAtZQhzYypkfXWWdE/w0/64B3vPZJoltY
t3eGH905u3XyVSfwy6TZ1z762hdy/Iih0rn+N1nXsgGP1cesJ5akX1twdvoC5Mq6uLIq7L39SVa1
0ZXnQ5NxZQwr5+kWu5dq8hEOlP8jU6YLgn+yz5Nmm01HzUs+lUkXzp5nYKsssG1/1YXeEdcvmzNi
5u++p4bbO7E81PHqShKQ+qDiQMmJLy0c5XDWhSH9r+H7lhjOe+Tzb4Ly1C0DOnn8eq28tdZmTMvb
TvuK4Qk18Lj6snMjkQjcOGqelmemRBX/gHyLExhDizIGWX1U+/YMbOrSIpL0cWQzRtmkTAfSQXtW
y8Ny87w2aOqfF6H2ll7jHmNOumSdSpN/umVb5ML8Afu1H1CfQn1KXoRwqhHsyYzciRbbv3noxV1+
dfj/S/Yo9Iqq1nyo2mFpkVyNCHHHgwzbDFfyhEEZq1fsBwvxSxJyHYem0f2cZHDgiKoq7znaJzHL
v15QUNbcyuOHs2LvH5D/N4VfFKt/vyCzAxuEfGQIakv3hZgZ1YKXIfigwAUkysahVXFqblBjBd8V
ZpJW0U6pTCxC1saHXVcwAYOv1SrnYEYtC2dnDvbRuqAwljtzlj9O2H7nMgIyMCwz6uomgmp7+h7V
xAAmuLaI+SMWNZxIW60bIO73TYGk6ZDZi90U+GFzyS9jD4f4+iCphaqu2KDXhlG0MocFY1KxsS2T
kKGfz83XUPoqtDo/DZxI5yMTapfIltDUrOhwTKizEov17vcZZKQVKlDdxptRs3flEOSp988rcgmx
kqgKAsh3DDaWfiz6u6/ysOs9edk55SO0NspA0jO/hRaLXY5GRIJS30zQUrBjin4ECgOIw7w3paSk
4IzgRb49V2ia3nZ2/BfU+NtGQ7x5MIuzHdrnkbJx5KHYpV1tlXI4kzlZU2M2tUt47tdR1ImYDpzp
e/vB0WtrwFtInSZNDYKBMEABDnkis61kKs1A0KAwyGV7t5xCkW3QB2vvhcK8rg4gBQ5/GjqzLHfr
XhhbRoR6q17eZNAG4W73wLUnI6WTqPEtY5iD8+e+M5c0BZO1jSbErawU1Pnc8FeoY41oC8lJZleG
sTTcM5fGOcEGfOfEnBfjzTQL+HMusyUlG/7933UVhW6RSNL5B3CWq+4BJQNS8z9TP9cRVEJ29QS2
MZy7Sguem/mqxFob4usGaLpyauZAYPnEA6DZsxtGLtAL5EsRMYH+0lOEK2gxsn0vIWKrdDsxw8Rk
DRMXoapKyqildMIP1lmwpWlKWI2tYbW0MDm/BQugYeUtb37okzAjjQEa4XXZ7CVdP3RFpjDltVs+
XIO18z4PXvv64fV6KxA4OU+OUUoGQ2Lk7WsBiAao/rTe0p98riGq90e3+o8caO1NU1ygGjaLrp5n
wj8nz/6jpgmtUprctAjBQLncEZzpO2rmdIPJ+jeLj5RH8f/6v3Eafwfw2i43L9NL4BVeSF1MRLMm
WWA0PVkmBm5MJF5ruWanhZ3Ksopwu4/DYUmbD2sQhGKV5nTAS49V4Dw42/VIsylB3DzUbdTg4cER
kSdZx53DD4XhseBR1eyeNVCwpP6xXd9DugOn2ImLU99mUOakBvDxbwPWcdtwgIUFfFQlxbsPj+WR
vL/GvlabQ3N0Bs6WHTmRb+P49/Mh4CYwyjxJimay7rXnipzCl6Ckp9OFVrYN4br18x0B08ox4dpx
SkZuvjMuEvVnOEZOVRjD9t2ZK9G+gMp1J6PgNBrwAW+EGs/mq7buPMH1cSWNxy2vol+a8Cu8HaC0
AYy7VUP98Z1CTg3ymUCm8+nz8zbk7XSmjBVZwATSwH9j081Krc28eDjPXri/+bGhNC8ymKmXscWz
Qp6d0QRQaigwtofQUqZlBYaEYaDG0A5IYzkPGYOPmTk8MksypuY0iL0cZmR79Y5SbciMBhE+kQYZ
313Q+OHowJ+slIdx8+vz4gFihBKkUnM9WLFZJSIapO/rygpoVBlM0J2ubvlIkAiIPClDf891vN8D
+7qTS7g/4HUPc2q+/SaDEd/8D4h/8u5Hgf4WvM10Z2aSwpph8TwKP/Hh5aAWZ0+BkwwZgweG40qn
8t2e3J3jxeZUiDzMLxhwK1GwcBReOECcRizqfj+1IxlhUNEn7+UepuxHgxbWwyksnyE21bFu5p/Y
MPyBvbdAWc6CgTvVAbEDdGDFV0NPQyf/oLY+IU82ACklC04hJZGPEB+BLFvAseNbKUERi4adyGvh
zXcs9j0nHLz7pV/LBzhooQkKY++moNehTPjC2/RvE6w364rl+EqNh5AfcjQmIVMtqmvXB+W0O1Ve
+6MpklXOSRnyud4Y3nYzix2yG9V+cD4mB3Cy37qg0dLAJf9grU4wNBG9Ww7osB+rhvMD9kv7WEWI
xzYDU15t6Cq7uHFv7BoWDJPh9pXF3WzWHr97YWZ2kUwfCk8KtPGSZsVtSrDU+FwlEgTzrsi/biA5
Sq0HIv4T7vbNNZYtOsC7QlRTOK395/M8bk91pJFqjZjB6eWXnI3ucjSyERgKxpCXL7kECzSOVD9P
sU4z6kUB9h2tPQFHgFRxjeU1cbFSiqEWPLLjzqgyp5U2rCbgl4QY9ymETA6+evV5gBWalTINCQ01
SlaqZ58qoDGsq5UBtxleXBQzO8VWR6LiTeafaQRpDp1vUYYkTfwVwb1daKnL+VIAtymdPZDgRPla
hHmWZqq1KEMEsrGzodw2cvXXt0jR2C0cFQErKCu2NhWgNbvQHImxx4GitOeRRufQhmXyxTSkSrKs
S62ofVwEjLBIm1bZUPXrUnSPm9hwBhg14zj2uqdi7WZp/zIi5tAKXmJK4tf2DLiFF9yXY+SGQx1O
4WrzvvolsMT9UffNdRyRXwlfJOTruJ+X1DKT4l3QIfJk15HHZqekTNYStWeBbe5FTs24OHRN/8s9
i7aAxNeyr0MSuzKW5ccqqAIYygCrQlVzcAe2HovEKQOyDWmY7d2wplfJsBtbXZnBujVYeJE0snwd
FcrNGo7pw+qLhtozOZw493rR06e3g6Uvaiis0Y616KBQG1pZ/KL1J2z5vhmSarke0HJMpnJ28Frv
VaQL973/A+6JLbre7qdkhb+OrvFxxJFTTRnadyumDVIr6DHfUIiUiXu318pZA/Q9NuP8BR/UbJly
hUpse5P0VXCmrdvTbEeuz4Xfx8H9eTD6iGA0CN9dHAO8D2RbbaTI/YvFHRHcOqORnGpcojICrOGz
vSe0woKIxYU6GRv7SFn1d+oIgtvifZYaoFA73IdzlaHvnRl0upz3rTxZv3I2J+fz4d2oqEfVp6SC
u+nC74RUjKcd+ihen5BtRKFw9jr3LDiTHmYMWoxJLJt8qMOk46i0hrW32q/Cn6r1OsuWXiqhyIvb
urSqDSZR1afWewZwyDirU6OU3o8Q2VAZCTzPKrNgpNps9ItEH3uU6qiTbJmf3A8E1Pc4cacxCPs1
hb+ngCqwdtp0mdf4EG9Qum/IBudQf1Dcfv6YQ+0wuInY6YhM76m2it22jsINQiMtfk6weU3aoFAI
zJQcd65zp9zQ4eQZ/MjNjjNT+6knd4kSzr9fiRSLbCD3uXKvRQpLDNJuhPecn9mo0RnYBbYc9chK
t2cHC7KU75TbQh6gj0MtXEP8wgrIxawkVCqay5H9/EcWzOzL4R0NyoE1boC4jH83JuHakNTJU/hx
GTXs8MH/5giQx6xLJpn6lceOZ61VST4rqhv3j6MdAV1yYAsSWyy/EQbxErLPTr8V28V37EgAbiOf
clT/A5ul881776cA5ZH8zJUwgtuzz3YcZ0vdzHm6H/f/Av8OxOcf7NArfAMI6cTTPE72rpR766Ii
knVR+VBVK65m6PHhvWwpgyaP9Gcs2CSP6aDF4ghzD9Juou0dsg0jU7LRuBCcuSTrzJ/83p6b5NCz
4ygE4FsCVexW4asyjRGzvMptzbgXFfI2VTKP1vZO8df/uNgMedbK0/kEM6mHv18zs00MCKSYBEyc
7H3ctq4jAxawhbRa7GcxA6RQYxDW4U0W5IBfXm3LFMs3o8CAmbPG6Jbf06NsNIuRUL5sVcxfrvhG
otLyepneKQ4rkv1yUD6i23TM223dvisF2PJW4IJ2MAa4DCQp4xjJOPaz761UTu4YFsVM1hpRBO2k
8d1e1uCMax2bqRGur/ecH1Q1hrfCqCohKhHUCfepU8DhLN/Kc+U4ffWgdGt+0fzw9AV8H43T4z2D
ruoT+095zbb8ERFozdU2V34CY7cukFbK2hBbJHUM6QAhgKdPR54PDsYPhK6Kp0QetOv6k8l2lFHg
mbY/ZUdi97LToW8UulqB83Pzh3PcoFRnNph/TCCtczVtrFrUxojV2Co1oetXdN6TG2ZdsWvAJPZV
2BOuum9eD0cr28uy/nFDQ4+lmvJbek8yNpDT0Xatt4njYsbayZfbTyh8G2tUnYFEASg7mpH1PlD+
G7cJJy2cLM8Oe84H4Ue8odYuFOM0UEVXJPjes2+dHs09OONEBP9let8cDpeO2F+Nsr5WgD27sYI+
qaHZfXQzXAVjPtqA/k5flKLsmHHsru8pjT+F4yY3dpb6gg6hdFbm6DT2Lee2OlZvAaFHpmCwaJE9
K+tF2N7bDSO6NZ/5OOsBpnpOtG7/5ZA4yduVYbQ82XhK/6EhFDzugu8rtUApqeCiErIShP7S99sf
9kWDYk7KtPduZPDssiOqUTE5JjYhinSYo1MbHF49JIAIUJEsXqm1Rn7UyHu8Ex5YlKfJ06Kv3DUj
ClO040sIr93h9hJ9iYCn6/hsNzJgWb2oY8EtoapqMKGV59b9wgkHO1MMGHC7uORCIVMypB5pNN1r
qg7YIa1koIt6XtbiYlGuvYF88srLDacDyWBGWlmZ0hynw9I5EFqyocghkAAC0JlpJwue9vhxO57/
r2lK70ILvjMmIwpy6DI1kXO2YkDKbVeKr7MEMpFnIMJIpmhKlo6neOvsGScoIh4Bl0opYtLx9y4Y
XbXJs+9/EIS4zmESh45oheE/tnCyhZm9xqkQfOFhJJvYd4zChlwgi92nTy1niy6htPVrdPFv+iNX
4cPj3RgQxh5Pxikfidv2ImOlqUlGTmLqIXeoNbl3hPO8cb71y4ged09VgJ08AEJW4xI54FL8U6Oe
xk//1kb2Cy8LlI4qINm80Cuai/NRrDPYetxWRTQ4Kq6qQBOeuKvc8lkcnfbJhYfT6HKQ22pBHo2+
S6hYKNHvSevEyzDIZYFUE0b2LJzcHXhxK4RJY4AfsCYTxkug3t4NJ86DKDreMoUVSRepiv1sDiUe
GaC2Vtd2Daol6HaNUM5SCOMR11jcn8AqlCvMitJu1JJDyum1g+BTUNgJD968HKA6GWM13tXsFDDK
wAGGGF1Lh1wSgljbt3AL1LHOSrhRh+EJyfG8w0Ec1xxu9vhggYODyV3eDTuUTqAvjyHIQZ7/jWKe
73FUKHsqaX4pC+bcvXkDL5rU2gbx9EdL/QYJq8BpvzK59ukMt+W7Yf2MJaCI4Z+Lst5cWmZZApZC
e84hY3DfT5yQjAR7w/+a/uxsr7g3YlFEXO4GNeM5c687MwvP+Uzs69nbwSOLQVTOG+fEj6P+aTfU
k5oWF0zKuJj9Al9zIKG0+7zD3BtFayVNDdVazGX14XvXq4IKSnx2BE6y9grYbl8pASZPyf7TZdfk
3JjAJ14CrxIAwfH7yyRMyhxkl9Qi5x7P5whECv9vj25HIceTqbHFKylcLy5YZfdlwlpCOx7KSxq7
6LHm/aEMg+2RoCFDE5Gwmm+3oXwbQitkpXy6zMHSInxxjeg902Z5dFsRLuDrzuKEwM6KWypcUnrh
phT3jXDfDtAKoflNw/5KzoKqg9uMPAaDeV4s9pHEAkHnGBv0m51sWqIUrsH18vmC5t/I8LKmuQ8N
8+AhY3AXzxNtUESiBoVCmQiFdOjl+Frj36KCFOekdema3V8pl//EHNYSMCEr7EJ4p3HcJNkyUzRq
JHd/ncy5f8j9OabPIfEb9KER4z4a2OnkuVnjqtFCm5O6wCs5/VeqVDfaYkPp8YaXs+jn6IopvDJl
NehwW7DpgAhEBikudkiTZ5nQS3KS/i/isF+qZF03YeAIwwIXhUtJXBrbNJOFyqMjjg4FHUV+aEB6
iGddoIi9ur/eMj0kwk96z6h567KnwEIS9SaQXVFKBxkh064r1cO6LqI7mB2ty7E3oPg9HGnMm/q+
lRK3PHYsPioWqaPEQckgDNsRWGaysFKR3M7oxSUQ/CBa3Mafs7cUkkiSeVBr+ECUoe0Kcb+9xkAJ
SivrmlIzIOdsqsWKec5t69orVA+jBmgg9wHit0OJTS9SyUr8joeWk5pZnCesKfDPuWBg4d9YhuP0
VwZPRkfSl3OeW792nP5XDt21aTF+AhgrlEuNJf1BRgxLpFqJwO9WKMDsBKQ1Ri2+5TalLVBFiW+p
XMAchW2Rsw9knfxnKAonKOcmtvDMAqUBnlbGOJ/Mt1ejWHSLnZNF6Gr640721m0Nw1k5Saf8rVVF
DnTQBpwfOlaZKNnPE2l3Q5ILNbNtKLNioZmMZSCWpI35aRZP2BHQFJK5EPBFBtE9qvLTuMxb9Tgz
LH2DreqtjqYhylp7Fy4RiYjdP+OpJGsPmJJpfP0StgsQqDfshaeM0iAhdPVB51grt6S7/kzJa1z2
F08a4tiCG2Zz5M2csY/3IoH4ezW3PmZUQzyYPXWyYlIxwgfBO3lmKy5aCO4abPcbyWygch9HDbMF
gwLi+X8e0JIWW02wFROuKIveZNOYWcBOO3QFuT/rDixIesIbgtUPEy+RXmbVVZdlnqJEqxYlzXjk
X3pLtGuTCy6XjKWKiaOYNskFAsBO/vSxZNBn+yNldQ/wkr8iNeb9aCpApEjI8OMTOafaYhZcMHUu
HmaMoATvX6cjB4a7kuhoCea8fc7olu+IRTw2vQNuFwB39+NhBZSiDPED/e78bS0eg75gPpOY8Ni4
31tae/UNxTuxSQIHh9oonmSDSFlICqEk6SL/VcYnse5AnkTHgvprO3m1RRKCzkCBQf/xMUafaJRQ
8COd1ZYGcA06lhA6xYmfRZbwIJ49jXfvfmTllI7rylP1Q5Rq1IMkKkYp1mE3i0PNG2I+POm4UQ3z
hNlL6B78bzr/A/youcv4KRSAepfY3mw7bJoKFRrDVcJqmoirsnCFRPAglxnCCZJ4m0TJQ9VR8Ofx
1lX05+gcI5ZKR+zuUryvFVaQzM6XMkYjtIUYSBBZrP8C7nZgrgzNMs7jdWctjhFCNDSI4Dftp6Ii
y7x7aXTwfS+WoDyEd+0A2K39WOgJw5LRYwOM2okrRQVs7mI8fat8SEOn7UdfUVMnU24BMXMQzCcu
rncZmKFo4T5L1NP9k3JD3uD35vMOn7Q4nNFUWVU+WKHga4Ifb3uEAUDMcXaKCtYXO0iH/idzbMOB
WLyTr/60psheXkqVBvlILkknjbAtJIYmruMPpUF/iGzv0F+RLWYxW2r8e1NG2VMkSswkw53BTcqf
VXCdMNJot9ZruariseFvH4FQP84ye4lkUPQsnP1pYpQX1XxenyOBwEHAUdVoyb8hTpOx6LvLO8Zj
WREzweSvbhFoOzj18cbh/otoe2/7zmVnkNe3kHk9Y657pUDwwUfg71X3y/73F+zuCNl1JEO4oCtP
f4LMi0iZ2jukoW1sNH9jEVjMayV1foE9xa24RG7a2g/eerxL6V7lLhOekOJtdP0MU2hN7IQFwe6r
UwspAsYmd9BeOdXfJkJ45eqSoU/hh3fas8a3fzUj7OnBmOO9ACQUX7E/cTokG7J0QNaonPLDBDNv
gAPXT3ebzVsIGSlIRwn88EpOTtTkpBVx6h4OjaixvhRzarAZ9FJ30FPgc9LOX7LXF+zzLJoOWpSW
bn3LffoY4cqJlRzhkkLu/Gae+VZhyW5rnbd8yzEDLKyZ0JZkaVBKcdG9bdJeAExRRUhT9jnt/61O
3xWZLd+g2UElVGizRBJyziECwuV2/yi5OFVSZ/xYvd7BXxy8Gs8ffe2AQOKqMKzj44kj19AGlEEX
4ijWLqXE/ULkvTx++1pD/79SC693RGZ+3RmNY1d9aLjYdMuFX2FFNCsJuP4wLvVYHETEk29ASzz9
34VgoscUWtE7ASmFXLQ7Ma8NAo714HjjfSKdFzCwO0JPH6PSJQysaD3FuMv74RQDvPEK3wMiL7wX
1XfeEN04/UcZjv5yWUewzEp9AM3KBuEnRZCUKhtlibJRNg88gPAR8vyU7JpCAEMjAZnBTYu3MYu3
dc/MkWgDJrBtkFHq7+CMgn6BUOdM1rQdmbWFVcggcGwyztCsdkAq5zkpHJHe9qJZewP+9KeeHuc1
GGn7yucBUp4kLfq8+6jQv3UWlhXEgMg+575CSNQHK6CybyHsX60KaFesoTYJWggU5bcjQ56B0cJh
yWiF9agQDQcxO7ZVA2CoJ8vS9VEIIb2u/l9hOa31euBi/8MDcaiHLNAek6Hq8SSkh9jyPXPcRNAu
8NyZ7banrY/2yVnexmUSNEyqRG8wyZx8VMFh7cJ7DPdKuZTr2xRxYvYEMOURuMSZjGvXF6HLLHZI
GFq4QSOTtsZAva3sz2Td/O/xQy12GnJc17dK1SYsQrK46GePu8USjxfOWo6c+bXS7p4M4bRwFx8K
JNfL1mIGW0gnlNeJSTmeVfLTIEWPqCIKiKZ58nzE8BweQSpLAqN7jQMC584aJq8fd9Qa3fdZsaAR
H8upTYtJi0UBEpJlEtZWg6VtZU5PGP1ScUzeM7ksue3Sdk431K965dk2wJ8jRtk59ekudF9MoMHT
cLqO9IHTDAtcFKQuEoPIp1Vi5mcgx4mTVGbe2+YJ99yj0zY2H2o9oMGrE+dr1ul2mm9FakHd0jIj
pD/N5XS9Jgu95mbn0v57Wp3PyI0jQ1bfXNWI7bGHDzpnyhjVex609CKEvayjEhB6p+BWLgDrN/Rz
vnQnphLDS5EITii6uBED8nheWoxHpLDtZBi5Zs8bsqiNeOXO3Kqnr66IpL3rN8A2FXPqNJCBKVA4
igtsTZpXGpYIraGa2RtZHPYY6tZtNpnxwdtnsoV0Te9b4JEE+rGvWGYBpbEREB0yQ840OzQqrc8V
ONCItevfBLoVNz7BWzVZQiY2CWprFrLvPbS7h0cVpxBE6LwMXgP+kmqyFf1sYtykHCu6zHwZI/NG
zvmncmKvD2STcq5l4kAQ8Bd05g4S2oignxNyOuCdZ/rPejdFc3PRonAd4qmyBT265yBVgF7EC74B
69XaJaKgA936CWu/jJTnFYAOq8Z7kWx9f61H6Wb7S/NoW6ef7kpH7Fe7e3jZmTnEdJadZK8yK2TD
h79ehAwDJTtKmKivIKsw6SLf2iM6Lh7iP0wWpOXKckGJkaSsO9c0/s6kGXPvGx5IHKnfnjSsKWR+
Wxv4N7bOWslu6ykP8xrtHQZoi4EGtql6Rreb0abRHb1gCvH4njIj6IJhT7VRInsr7iMUkCKEw389
Vtiwm5V+YLcCnvXhu0eFzUBq4WhM6IRvZcLEGg31dP33nR+Hm0sBpn45BAutKlp2uSlLozYF69O8
2sc1dSvTvfXStRTXMPbZ5IB7YLDAUGgOhyTXIMHOws2ui1qhdHmwbfLaIMviX9DA18TCcUmamrql
snf1QF2b+2MJf9sJBVEtVQPqcwUFWQCHGUOwS+AcAwa+RQvXm/C/P2kkEqiK6Eym1S41TG3Yhe4a
2Bz5p6h/5SuqnX0LuQs6XG0fYV+bWWt3ClN4i3QL1Z1A1MtkdMbaM/SkwnXJ8NrzuJxJVxcylmFZ
nhaAq6OiKNM6UrzuFQPsTJ4YDpNC47XA7PXrPxxhNTcvaipe1KzKG5JYwce4HX1NUGFTpM6gefcR
Mm0Q0x2yMlXbProq7cSyICLxZL/UXFD2qiMsoZ8K7U+P2XHKqsa3GUS1ID55PzeEO1CjwT8dxpDu
Q4jevRMyaqbbEqMcL+bfaWscBgPBfIHDewV9iyXA8jmtGq7d77nD3XQOxWLzOQdMax4fqhLPcmAk
AqlP7uOiAwa91ChTCGVxGz01xENtSddg6RCeUgjGgGnXCMYBBRZLtkQrjU2DxsbYYPWQPH03ztGE
dg9AydD32tJlA1/upNlOA01+K2/zzicTpa+5fdBLsuEsDVMddSy5SjrDNKE9+xYLDINzxy+Wfth3
EduDdNEVIE4unDEnndxYMO0UhTthVzLve6DBx9Im7aZ9IDNE22e3d4VtJYFfAzLN4SKJ3kuxsZN6
1h5zSvKFkoS/jkqr65NCf96S9O32PiDfmXFsPnUU8MLKX2Mar8EDaXOFWiunWenY2VdTvSbTrO4X
isvwP2KwWECF9mkW3cS7AhBEWEHdmPKPd5ZW9rAWT41x82ytFo5sLdTqZFWRBvKwSsTLbwk3GGlV
kqgQrk5GS9LqfdV3oT11U3e/9FwcB5ZPgnC2edWt9oG38oBjCGzhcmb1P6BaJFjUMAqEs3npWrsN
obA4+bBsh7GtELXHdEBK/9unrXtIEIy7y60Oi5zpk9yDy9oBfM4jtskrZFDDtvehSrffsWw0vFR7
ju/r8bGznwJ5kxuDH55SRI0bwszuN20ZPkqo8Fe1y3020+ulCFsRFO/2lB5DOWOjtqoMyfohY3YZ
gFAtC8/2fsqYBW0oa4Dp0iy8AfJV2nAmGCIzNzOvq5ZslM5yeZJ6F12cMcvoDPS6oXcZZ7AFhJEs
L/bOKnE213lgVCoN+XgK1chrY7ThD/Ip4nW1iblTUilZDuRjdrUhoRoNvkplCvR62tI4pYqw2LQ+
JYsP7qX4VoZ6VWHK3BObRbtcGO3K937i1NXxD4p47TSxIUj2EEBGpfoKu3+UPJ3ehzJYlSn1AXUb
Ywi0S98FYq0NbHk8WDcLcuzZqDJ925Yd5bpSB+JfE17WXtEcnZBg3OH5Tv8nbsVjP0DCzM6Z7Gee
yTNzp3EnTpmwIKgOtsaAjbTsjsSajw8G5VJjX2ARVjlmYfOFXTF1pJXODcoW8X8kHfxEejIzIKV5
BZhGO57zZhNV6/IHiEcHgw7k4BvQKtTHOuZh2HTDefit9ogYTiXl3QF/AHVdSruGw6sH4WIUvT+C
sIKwxs5rQIdWVGh59QV4H/wEQrYFFdC/8rXG/UVVPO7yX6R95vsxf0OwCLZnVFJGNnGQ12LBxHxu
ibUu2oz22zj4vn00GDsgkcLrO48jX5Iv8kvs4w2dWd7qcoOOok5tPtK7G1Bo7iWAx1Y7ay4mSnOu
r1PRlU8wD5gSmnyR/uAf1b4pZI73wDWEj3TRK8+zXAF/84Tynbkt1ydZymiQY5beooJbKwClBJBs
ZpdQ0SbDZ3WY0xO+ZsGfZzgcX/PcZLzFRVq07orqJXsIBi6py7gEVJ/ApgCI0ykNnDB+SmptxKeA
9bg6wSpAm2BMS0jn8PTGiyObOpMMztx+RZoV/EcnsRHxj1vbe0vNsT3iGdhSZE6j1ahathFTAkJw
QuqMypPFnSJ1PzHH/YNJuKflN1SbQk2bFoudIceOeNlJ8Q7MjbhyrJMw+U2L7obcMtSRWuJB/t9f
qtkArHNQ4pUEtdbuEWIJMRv+7XtZtezrDB4C1d4t1bAulJ+IkLy1Cn6anJ/QFLQ6O7p0gEvX2dYm
ZJTF1B+3PUBXVgmJTpwek2Do1iBJu4LNW8fGf8wtS6hckObWZ1euz/rIVl/oNUab6PS4f6aKL2VJ
v6ux0k6HjRVd/m4gbSQveswAWMkMgX9LwxRDNeagZpq0F34dKDXHSWgBjBCeFcZ8KoTWdCUXCOFt
e740K91IcnH/XvmHjVjAQC7DWsNzKZ6rdlK/V8/m2ZsCYeRFIJGsXeffLqfG6UyEpZfUytUUunA8
B552/976SPZpdCOpXcrkRZmGd8NznN3bY1K+SArCs/2Scgu5B/0lVf4Vw4iccudrfpROnCKZ5EdT
WN+UhabUyMQm7vjabBtGM6usiWZTnX+AOnoyX5IOpffhv+fRMg9co+oOySJzD1QIeov9Jesz5rW/
/NSJHkCJcRpH05ofdp4K9bCyVS1rJJxqGh5Tf60sZ463oc1e04pjV7Q7lVcumJCdHXhiet8uv6nq
0nFX8JB0WxxoAoWi6wK5dnu1k6BIKm+PCTsZqzpB4M4FFBv6ZFkqiWcuwM2cJoe9MFoj/Y5FDcUy
DZiccNsX6eRXFVlQDIS8s+5lPO95UMqBvZl5cL9yo4je3j/+RIO+xh3MjYa157+V8Qno4ewwbgzv
hhM6YB/arbJp4aGBYRUU6dizdbUJH0Bb5FgQ0nYbMTTFRyoNKjnXG20kCvO5XpVgI7ksvlIodlsj
scYTE4THDqt9JWfGlZBLd6/Pdnh51bM1NewFgaqVGkG5xSwb/XBhaQ7RvcisICXC7U8gTgqDx7pb
uFsTtQX6oe0eCKeMP/MpbemcX1erLD03mtzAwbaVaBiVycqwQV//LvK5KF6pDJbzw+Zk1ilhcru2
BvF5n7meaS70ihKl4Q9nSr8jh54JouiR2hZGoQ75Xq4Y4/F/uwYoiLnpowDpEY3rESgktvOJDYGJ
vQSf0nBOZUPa9z48Y9MmKWJdWL3ypeQRphYJ10XfM5c1Akh/BpSdLRi+6xZv2ye+ZNBETz4lIsUM
QAzLywa96w3W9V8ADUzvZekLICPj2ZR44EFxUkPJtvyYVQkqsYekhNa46r5ONBPgRCrwuYMAcgTf
+R7q1ppmrBrsJ+6pccg4B1MzvAVJHiwjrrvd8rOcF1A7WR7afEoyF7RexmD+6qKtGG5QJVpEHdRT
aPZVSg71YtpdZAJ5tsVKYcl5wZaSs9L/N+d/6HMAwMxPCrfyQ+41DRQUoPFmwtQZwcz+6gBhelFq
bZStuTwPm8Me5WJRBl9RO8CyqHnRkI1gwf1ia7NhGtqpoCW0y5vGb4WniDw6SQjaY5Agwem/yYOm
iR3Ylqt4VuLGsLEtel2yb7FYZpYlCtz3U8nO2c6QZlaDBuxFzFjZM1z/VCJqSI5itsFwZtSRYAwV
HgGKqiruRjJskuKUSzlO+pGqk0DlsGxESFHPW7rZbAgwArD56ePaBG4JQRlehJskFDI+CmHvGOSv
8kIicULP66nWv2Lj8B6tK5GlO82ha1925pcXhakBjz5bLKiJjbjlTH2WiewEyJKbESvNoQY5Xq0R
s50QKb5OT4dpDXAi/02RoEl3wNPM+Qaqyk0G1KA3525gaGNakc0Sx3G5bIv0yJlcfqVeWEDdy9Jk
U31hk42EKUTDG9wkK61uX0VR1bJbbJn4AeD/i8wimF8eQkQ5hTqeYYMWBw3RMpKZSJSgrvemyBmB
A2feSkcQCwp3CQ5ZnDrfeKxpiTYKVeMMLuCFqSyH0L0H04CZ0mOCNOy79fbuDqtomtqdARo9UE0h
HSqkzcAvPnZJXGnECmRicUjqDXKZ0nxQGPM4+3WDXuEr/hc7mPHC7h+6QzLKedRY9FpiPQFKEExK
0oxBp3+e8UW/VFuRMiaazGHMWenC7u3Ao/0vQgdakiGlND8YVzSS9DR3q/exIwqBjqZIcTU5jhpT
BkaI7/BSi+VvIo7hnR1MLHTb5PuoLTYOdrOw0XFlJ2eGW+bxcWBbDsQfgzxKO2VMJT1heOVKOmb4
cbMc9IURPpLJLWD+MjYVosv5NMn/i93g3IwXXvgIFCNgHBBZHt7Qfneyzca0VPwO5lE5kK8bb4Kd
eUSykOZMwgxFRZTUVM6lJ4tOf7IHcLJNpE9s4Buz2cvF0ET7WfdKTY317OFQFqyItyatcKxWKv5F
xoIKQkmVz9UAj3V55AVqaI887yUfgT/BQXtnVD2CTlTToqC+2esvK6Xs58nsgIIYPB9++iEFjaMZ
dG0Teoll+dBRQAchAbr5mhFv706pfj0LoaQvkyKMu959u6z3shLe6irwM27mpgyap9r7T0JbABPW
vJ7dxdnEDd/YnetG3tVB+28DOCxHIPBwsVAK8k1se6TngfOGwLRfcz5S3itD+euCQ5LKIM3K3w+I
hn5yysiT1Q/X5Pt4TwBFpzHFYB4HdbtNdPKtehenESZPYSGTv1QlWSXhKK7faY+VimyMY64S/1My
wpDwQk/3jc0q3AAgSwOTEJkk287sEfyYsWIqpYzgMIFFF5lTKHUxePv+fGO8ikQVuI3p7JzV/K9V
8hNFW2VbQDTMt7ze8N8WureLsmExFNwElwz9urRR3N7PKao+LAAaJiSRDdx5KwIhrYdxNMavWd1s
7zsfmrNhn1EBbgYCxf7IkZfOEgs4Xt3AT+eJdwMSwTRQrJW1uPqZMXWT/yywvkYC842Ux8jzuE5q
DXKXOIPoTChXttJ4qoHwLscT5c6Yu5zO4npOGcYEU3fTTx18BsUVRtAi10DgAx+MnhRhfH9fRvHc
cT2Hj52xtFvtE05i7XP9PkgAIngEBEts+Z5toziILTTB/S9DHwy44eexDGc8n3RoJPti2oHe82NV
PKFbtFvifK3ZuSFKdsxdSJlS0rJrTFOFU1Zscq6pwwQEhRSoGjIOVRQGLDXSHx2QC7g/yYWatxw/
Js0qOruuZ6lSo/dUAKqR8p6TncXxIWAyyujC9Nz0xg2DmOTYarItRbjabjfZu1TJ1uyfA/jnXEA0
P80xgJiQQw5AsxpMrsG0/m7fXipxEVX6ivilbwdkLW3CiWdOpL3YoS0LOJzJpk11k37YRRiJvnmi
ZHIkrh1kJsTcPVVjkMMhvceozDqGH22UXkXsc8xGgGHprOdjyNtpUQMVHz7xO6RRTPLI9Tm0AJ8I
GJAO6tYHUFme4YcqzMY1b7ysrP6H+4enCzw5pztkPk9Ak+zzIrAYk28/buQXZpLZ77jYeKePLiW5
zdOSPHPtuNpYOKZVTa1OILFVXZmUrlNFskjPgljVK7xMJnVl2++WIS07IF5yAAIXdeJT/O9d8COE
sn8SBpUyCDpT2yl5mxtxsckkinT9rMH4eWUmXiAOpLKVHiY9qmjDYxpHwOLlKuQxvHDUHnaW9d7J
C/SXrBHY7PIyklFSbNsb0Vg4/LziFTcUhz4q3xYNJZ5SR+Mc+s8yqWSSftityAa1cZN3/Clu5muc
/UdcsAlg8SVrds38tCm+U3ILFoLejvzpDUx/KOQvH8dgSy66faRixKoqWvvr6dwhynPDGqlFoPxp
lIhtjCgonvsmySHWnZjpKJv3ogKTwWim1+Je6LMdl/MsJoVJrbd26ZKvB4sK6OsejEDdcXeHYxk2
f1Bh/fiXY6fs3gYp9q41UEKh/YaXxRcLYZW7vvDQa6zWLoo4EE57o7hMvuiH2Np+2lAmhmCNq8/T
GokNT1Q8dx4gYYdWufERMbPEGX+dCXmi5wrD73/dlkd9vzl9hu18dXkvsPnGfiJ10es+SRhzJiVu
vyC8BSG9oYzQmOhg6kLU5KQD0jox7em5lS5/sLsf+CszrTnpMCdYRllDN7PLhCZSgezCiq1tKtZD
Kwdqjbsr6T+pLeVQ3HIWfWbXydAkmq7Kgu8e5TOfBq37mik3ax4mV3q+7PxXWPF7UjgYxTo8OPhe
6dlGRkure19LRYO2RpU/XgpcaQssKFpddWp/9Y83kAmHcM3JyiBvtotomXRGs5NHsVORcQGpZq3F
ukTpKQTogQKurQY1P/fq5tW5TZ+Rif+MqjErAYULzkQXZlJsK0v8AgDY12vTNmMstdxvQUpxvgu9
dLkea0K+k/w0vGktB5LnMOCfg5Tdw/mxxZPlAOBJfL29IDzz87itoctS/QUx7NrsPDX08N1aiKXI
Chttviq5bXG3Q8pGc6bl0FgVPcea39fqQIE1dXL9UKOD7F1X67TYx7Xj9rDht9eFsm/xoRNJdEK2
qUzrNsg/PE/qbR37frvBZb+34MWmg7v60kQjUz2H+fk3mzKApQOBCu64KUOoBEP+SEBAuNnYHT9A
BtoKlSIBIUkc9vxIlyaOuxMITy358qkuHaV13nUBzoPMb5AFc6l3W1AtiF0EMXRejeHUOCMZLOeI
1sGJqpryVhQSaBMX3koroj9rmARKm7LECyM//kSARvLAfk3F40fZZp/AL81UUlehDskqai/Xv63C
DAZDxdTLTpYz8vj9AJanKWf4XulPS10srOO2vpAZRqr0OgJ9CovIgF+DYLPqiG4+FL0QA/88aBkT
sKqfIuEH/I8AbY3tJ17RXKT2gh3pvaVWl55iMpv65kzya/5RZ9w+ms7tsPUXWQwSHcrd+K3Dh8LM
klf3VcK85758fBBUgnyAuf469npv/5he7spzQRD1xYCO4oVjFcm+cks7eMnUbVigDVkds/BRMp02
ogjT8GgxVhw9XNAMtbbf3fYikJqP4LiRG3xMii68NxZa4RRQ8KsIjdO01yH7bH6+7BVFmkRC0v37
8aASak9T05qUkvD7dqxLhenZlzN5dsSVf19z1Czp/N2sqNc8pPIktiRLuWfFIkkK+YKgglBsiN+6
lYkXuNFXP7oRNN7XVocGrafuxDqiZN9EGfQpZGvimY3CTKmXMyG+2rT5YFUNKJ1eGgO18INH7rIn
kMk/35jcyPkgq8/sNExo4peYpovpr4iCkeMA+zd75UnGzTiJXweYtnRjJPWxtWsqecwBmj2V0TC2
fS2vgXCFGoEeMYmQ9TFUczf7/uWn2aCM1tEzDnw4Bx/rOkCzA7B2FI21m3QljLH3L+wakWaTrqyH
huIy52QAW3SgtYNfFBgSTgL9YTYt71rL6/r+FL+6b/5eWU/aVr/Nk9FBPdx3gpnYB3w7AZ0pZDd8
czl5Kj/M0Cxwsqp9eGXKdx4EiGEfT7Uu8fHFZgJsCYJr1BIB9EhzkoD+PO+t80BLkbmWUxL57UBA
MaV8XoCLfl3h8awdsCFqpM4R9hi+UIwESIEVShL1avajPdVh2LeIn6n4ZMWtYMUvDmNUadtxt0vD
a8bbmRnObQzHFfg+6Pnj1r8a4rQOAZLmmUFxR2AEzaGLK33PaAshcnczRDRDGfzJnGIEG0oTp7nG
v3GavJK7n11cZKxekogKaCB5u2EwMCMhp9CIIYAsKKrU2KKVj5iPdMRmWtOLigKSbXBmnnlOZQSm
PycWgZ/z9BGF6qE+c/xh7YppbOqJvJ0PcF9coKZjn9RaA06IBNZ/SyvtPehRiuwFMoFtsEAsTod6
wdNc3E7m4vbyCkWCtMyuB4L+kivAF9tSY0B4Oirwm3DbqA0OYzJBn6sTOPrrGM/byNNMdWGiza24
vVc7QOXrGIrQY4bou+iNDf6oNS/RKa3Y7ZBnvT3+fwKhtI2y7SX2g7X7HKb3XXdawlAfyNme9DsA
OvBvNMeWhn6zNNuz83LGxvvEs7Ns+x7nVGzhUzDXquH4sZsoCPb751RBWInGuqBW+1U3IS1qVia1
f7cx1xFmElZkHTsheSOFhv9sRa2jJAmOBC5BGvD+eD8HbGTycjzBNKz/aiDMOeleOkhDNjoFVnOv
C7PPMGZhAbPZrkR9kDI/Zx4MN0KQrF3cp+a6V6RUvbNJzlW86lMjVxXb8DIqV5W+NFIQ8FsYOYVG
C08xiSlC/acleTI0yGjAnC6zrGuklCZ0tbryv2rpSRJanVmVFoqohSI5ajbkNcRis+ZsVU7NHnvg
h+/PrRAnlGKtg8Fb37i17gW9aq9D5FcQGMEjUfH85jb7NzV9K8PhPpqbXXkrjuhq3VCr1GCtyh8S
PZO596Xcvtc0B5tzDIcPRcWPcOro/w0OsxppPDW9kUWK2N0zSvxcaGrUn54cJKUGzt3IxsbB8Xy2
N8ziuSny+HAMzmA9/nrkJSLgPV8Iqf1BQqb+iRdbdZNz1ouy5yB69MzpCLOq0OpCeZUYDKMQ9Ur4
t3Hy77m1Syr6wy2+t2OllN5ePRGW8f5gJwn8oeKMH/4tU/FHZFc6BFtp4PCrD/pBQdSpBoBYvlOS
lSTyI/bdNcaynrTqz8XRNk6MWrPkWIBrykjK4Nm0sXOSxsq/H4nuTe0SXhr3nyvTDYT2HpAA9t1E
LNhzYbe+MjyRhURkHFG238erglIevS4EClyNYlafsJbiUG7/wvLKAWJvcIDgLcb3yGvc/yBKSLfm
zkd1kF/LMicl6QMKGTE6MJV8u+8kcFQ1pib/WMjl8abxWINxl9YbTaZl9bdVBSoc3zKTkV5yVFLD
i7MvOiApjseqMM9hs8nIIIRYSRfIgX3ibgwq7bfQ1oO5y6cxhfmfSar6ywit2kMt+brQoe0Su4U3
iW3vxbvDv59QKKtqyB/ikKGp1e4wBKlY88+3DRrGf5V8lAeQ9/sP29sgIe9bAv1tkmwEJnqXot89
cXoja/tooHMKtQ1fBavobk68qTrEuzRqaQj5eOn6n6VCLUyNfcYBiW0e2Fky1aI5T8x6PKZQtT1o
ooPg//H1ocrRQtRKDYLY/svw2gm6zSGL+jMTxu0sZhRBRROXhcT09AueLNup4oXUSsxZnz9rg2vp
R7Hjq7EbL8m1WHsRUfw28SRpWA6zYBNe6P+VNOdmyQPQSbTC5QdjzIudL6CRD99htMZNzAp7r3yw
OFoeJ0pg47wytdsG3CT7mDA4te3NWV4QokJZai45L6Rx6eXWdL4nfR+0TyaMndZtZsiqMVOLYUFW
trMhjz5ciKQSu+Ug5xdAwCeo0rKgj9xod9YOZ7/7eBvC4MorxT3MBjLLAD5ZUUmsa5PW3YXzoUcN
Xp9HdTTtpzOFCP0ag/pGwpM7StpX6GoFshpxFXWHu/agmQVq5d8iymSTyBPedecgAw+UCvLmzWGN
91Pc1xvVOz6FY1TkocuzRKPz4rynG448WeQjOgaK9bVBjov1HHNQwQT08LzMP1ZpWN3RVmFAEq+A
ObNfZQX3WDBUGIIg8YQFRLgD8LRVefS94nLkO6tKFFRAucL/p1hM7OF2yU8cev3eubuKadgJQJl3
OfOPkK/ZNfeO0Ge5v222Q7HOOmLNw7kl8BejRMtB1h09GAMZcNwwpb63Sz598E/n+v3HedQkNQaC
qu7i0VJe1i7iZrhhIbr1iT0raBMZUhUfhoVeXyKSVwBEEwNITbx7Ru/iunMRLrSrnij265hTrMnk
NTmfnFTXMMBlRHKdtFtpMO4muDouDeyqWBDvAegSC2A7duMrt33l6NssF/Qm46RPMPT16ctrELF6
Np9bBdLDdQK0HdP08DzvNwi9a8LhOBkCZO7hwn+qgPGIXxc5wWKLwaeINvpyhqx3GqQc6e6ar1iU
1Bbfs26BsN0Djs55agMSUhcsbXgnRRlIbSDl8Fij29uYhMcAe4wLjrNOEgqjxF1EL9Zh7p24bNNL
HK435kR3THCjyIRIc8dqlKGMSSgu1YokFj7QZZyKBy/0NRhTU/JWfUpW2DUFBAXT5LCRrccbJVtg
UvCvW1h6s4Nzs9A+RQarnzb4jJkqSTqWvXIJD//czrTR0s3+rPl2SjkJSvi7OtL8rtRBy04ND3YF
ekXcLHwWswtsTo983vKhKl3/nMfq60kYJpPyxl8OfVIvGcryXe7FWlgWSrOdpgtVxfXfvIi0Lw2w
LavvN60B9Uh7Sw9FPYF9z8mxmGTVG4Agj1WrEQ2MPqAM1ilxFLX39T3VStG1hfULtDasBLDXZiMZ
z8AztkwOAXLE1UV6Y0UsfLLQaHCbtmS5wSrYE6SUOL3yarBonJtfGuDdScVakK8CGyeSGkfUc9wa
+GI186N/6/QHXksMLjlBMC5bgWmymsOhaqYefQTAtf1eIAiYtBOaJ550cf4q1qd2mDNHLo1FI11D
GdXqdBiyqWnq3yrjUntQlFi39acM6qWPkr+rxbw+mUuvfmRuCh5tQrlhmRvZzNPVyF1czGxDV8pF
t2aZy7oaK6088T1f5GD0pUdUXRMKAFIbKkMYyffT+UrRy0rz3Cgv6BuhOQxUzg2Qkl+Bbl/cfXXy
GPTmPR2Mo270b8fOqpD6766NlIU425d5XaRqShDk18Mj3du4MeWShrysIwdqaNGEE+LKoKoO4U1v
V5zLkSLYGhWQHXhlvIQ7sZIw1Iqb9gLAmbsDe6UgYU1DeC/q60cFYJomz8L6xxJidyhvMI6vlHsr
Ij8aiPBpuhWZaBeVkSFT6cIgyh4whQ3p6SkwnUXZnpRKWmnM+QJD+7TrkbdNPuEz1tYs9Oo9aFZa
hSd/6vitDPxkRbGhztHETvQKkahQz8+QJXb51ZYNAUznXyzMHyymQvnAEcMktjv9ZqMeldpk1utN
ul7RylbQmsQaZxSL6woZD8+hGthAp4CN3KigyEhwvkj4gPySBt/FzNWPJHf2XAQiI2fpLsVios2V
ycWSqOv/8csR3p5F/WtuN6PR29/JwxKQAbmiAsF5pB7sjtjU06BRVGfNlnxXlIZ5D0mYuwlvTjrN
4ZnQNT5jjhw/hiJkZC6nzEgBvFX7aYI900Zuz+J4WVszPaIiSHMPGCd4ct3P2MIs7WgGXN7O7cPX
BTYvvvsjySNWh+T3zeu1nBq3IQ9dpe7B51XYXH9f/oR0N6K94RQ8HITfVeYqS9UBjy3CiM91uCVh
XCFe9IkF2GVR9qc/4cpgCjC49kgaD6jp+YPdaU3rsyhulBFtZ26rClb3esatTTfj+g5cusMs08EY
3Iea82lPahpKr/9Ut2EY69ZGEw4XwtN9hHihqjO4yVy1tCCVTBMLlD5Tx1nPW8IFbdpb5JDmUuCF
ml1g1zchPqyxMUK9NOGUMRmMzi00WmmEV6BKjHnRXL75c372n+iIY7KA9vynfRXtEGAryL2b8YeT
XoZDcnv+tF+9oA00fe2I4ipMglwdq4lmbTtCzsoMrVxAKkrYW4pxP/FFxd4ycfZwP/nhImgFOCPJ
JtAWty9F3J93KBtrnXAxvrsJaiRVvEgH/aQi9lLfiutRl6EnlsUH2YRuVqmd+VWjC4tUNr4j+yl3
yRWhcR9b5Xl/C3DnQ4l34FwoDoup+ZUwSokpMetu3m1hF3rgPK/VfseW8pvTFLg7of4wECoH4XZr
KJZsXzy5xWI+uLBQm8yXDPmsm2nWlBkdxt+CXQ00lLAkPi6rV8j0acEdbLoaWf+GKEc48rMstTKw
1y4/9BeQm3Y29XU3H9mdEoqyeAexzNzi/cUHvipOk8rEYkWk0i4ZolPiyXq0veTU1Tqoa3rqMqZD
/sfoPVemBmvwGotf+NLjTCJBSSakxNGMgJAZy5CAWyvcvpZoV+TGW0k1rdAYGzdt1IkGXj6VLTdA
h4R6dr2VwVOSJiIqy6HxCvHWYLaCy3mvIvfP24CrQGOFTt/ebL1Icad2UdxBmciONofsE5FG3Dbw
nHq3Fiaf0JI2eg/3IA/AX8ylYcOjLA+zXQmxtc0cz3HeS3hNs7NXfQX4/92Fd5nrpXWffFVea49c
8Frpe0sXk+U11p1OEqbNME8nk537c9+a8LbU9J3rK6N2DyrjtSi/UN15yIM4gU8bPZO1SwfyquLI
3JcBMrqwhweMBwb4sRb122dRW8AyryameGPJp3Y37PDsg4ThEILvQJMFD3gRe/tUDGFOovWMBv6+
KfBHfsPxtukjEglB0UYoaKYbCX25IZVzAACiAzaZZoi6msElwT14ACToeialU5bP+wSHppxwOf/b
bAUwwpZTL6NuNJX34WgzQTc7fPAr4UIma1NK2n884ezqIV971rzb3N3t7w/pzqlMUXAZY83aokqq
9AMcSAWzYIm+mFjS9XOD5Ag6bNW9O2kHymlFyN90MDG70Jmwq68oyYi0u0438dbMlWDlODQry8ft
IJ51/8k4g7TfEqWcp8ZjpvdY3/e/PzjYVdXWUUkx1+ZvtU7QNp1Y2XnBeelOvLe23QUJSvT82o9n
P4c/pbzMxDasA1WA9J3XS83MXa4YI6LSx99TZjzQzU4HuIGetUcMWm9GtxZQPcV2kQ60CWTcW8M7
M7z1uy8w6mp49SvXQSZCf8eWFaqNaG/iq3e15nq4ZM3osgPVEHIDPGo6tDI+7SRS8ukauoPj3nfJ
fZQ14wL8ixmXAw2r2WGKfJPwKJI/u/XOVD+E5d17nzAERjhYvNioEOEGLxqVuu0F5YNq8cAgdSIZ
UMN2jMGqBx3pNHntIGkV3wvzrRZGOaqNs6IeH+fdKvIvhBb9bxmw3mg2hTUSdo4W48CoLhQ9wDX5
8jtARkyP8aQO/q2epCn4T3yOWElW0VsI6FpRmqI82+NRxapCa7UN57V6P/jGNb50AAOiNo8uJJrS
d2qKg/m1VtmRN4RIVFq9ckzI/2lAcd+oEvfuhFrVnSMdHE9ULXg+QjqCXvrWTwViDbxYWh7+Ytyt
UocPaZx/kCo9hh1UCcajWnOe0JObi9Y3PIAowG52Ld6gpmYOKHYbA9zvs4e6iIHkuh/9ne74ZSvB
tldvUc5uA8xscKCsdKjBynZwLe7AyrGVpPzV58sqEkKm0pNZzdMITRFmMvCvvtSenxKqVqmUeCvj
wYKY1bPtPs2ux0KbGYGVMv12C3bRhBiVYPRKEUX1D6bIjsMGdgqJnTeTW+c0NBtBremwJVoj/pwe
6GQ7n7DUXmoHp8cy5SKOrMCBNsBK84O9yH9V3e58O/sK6Yzha5OupEwxpTBtFu7L53A3eSS5zyjP
xca8gaByE5/HbFMdMwAbHK78T7hgbQKjRqOKoWS0qn9JrvPJYiUNJLCyhiHBYuyI059ePCMyDxJI
UbX/u5IXlfWOiGjjL1ExGStaWlbikaOKQcMiQglCvOxs9wbL44BrbXcqA44uv4GZLaKc7rCwofW8
nIh5A8tdtW6ZlV+Be4mthH6zxf1MHP8TFpyq0iPGjXRd10czkIdSgCDcWg9+LVuihSiXQZ5tuuYr
/knJEVp97+uMqJhd9ZZLjRiw9yXqaMroImwSvu0y/ugDi9SK7BwLls4Hfsp0i485WKy6rVb4zZQq
XxwzlRnYvZ7AD74IGHeNc2HOft3phj18uYEQROFKjJ5Bd69FmGjQfFtF7TmvVPC7BUhkVfou8On1
hxwbvfv/Wv4RK8QqUqBRYJaQ1qzXplDo1smj9ZgacordnZiUDGDqCf5sAOizeAIguc/jHDcZTMci
JpfKHz9fgnnUyt2J4zE4o9aniGItRgTNOwUQx1x50HhgeXxwkSf5HNJ0WxZ4nO+wtuZV9+oHansc
/+ASbVJNW0nuoabvB8wyxu513nsiQMlg5oFdpaB24lJ/QCt/tL/P+9hDGcJz9iUDUQ8vc/m6svSh
D81KoBl1ZnxTamTngrSa/QbR8zUJXeoXF5ixGLbhyE1m/lKm59coHzo98QKhfO+c9K34B0phajgm
RD4Xhq6TA9SgHDFChzyHtFzRhG+wmy6rMghM2Z/ahJ06y7OW7JofUpD3FJrhE8FvKFlg1H9udHds
jJVmQUOS2i3U0ulsxBR6KphcwXS4/3M6NZtK1qBDYMnJUK3DROV1MXz4HeUuuvzxfor23bQvXnHL
EhpafQ2PDG0lUigu3AMgnERTOo79aY3spGB9G37L15L9bnRujaeWpnxVCEYU1EadZuK7n54uGdOI
qX2j2ViXPJOlFTYnFNgemxjsoSE563xqWTEUwksO0oXSTPfuC/lM2pZ0ieK8/C53H2pZiSwK8jsu
KdaLkHHjevmhmiyeoAKMVeqrFyZ5FRYaSs6j08oXo7L048cjy47w52svfk+cEgLoM4D+hcZDplH3
uiLUCXC9XMe1NTeZkBSHbHrweHhIz0QfFwU31IYDJwo9y70/bvFJI48CDCI5krn44X3Sr3hcgpZq
AHoBOgwR+bp1TZUG0a4JYYEfOEoTJ/NgiKFqzU8404ex74KDgec36GO0vlRKem24BP1S6zOh+Amh
yc2PbLsmddB36xXryeraA+8b882Mf/Pg/+yOT6UU9O0DdtzIlM1k7hMlBgg7qsON8X+5FUGoiqzU
5NRDxr/1nphXJnm4Soy5oeLgmFo+q9E5ZoVyWvg7vSfPaQSIIafo7nRKfyiM9sOJbpP5sPR0Xd6U
yxHGf9XWm4LcK1wuSPDj3u7NpSHie3lXIOYM1U6XVDGxkDgInBvqQgX8q2UwkgLqDb+eN/Dj39sa
OqWOpGgY+wSZilnPQziBi8HtiQ8Q3eOwuDE0iOV/aE1VvHNUTsn2dR58Zd+cccm6CcAINpx/0QlZ
RGB0WT8t7tLKMDG/HNeAs+UYVlJqyl1p1NS1HBDymG3GQIvnhy2hnY6OCxoRMS4HbBHPXiIUsqYX
CavTiLUJUROYBEptuRyeDddHOuwA2GQ6XTI/VYX+Yy52g/VrSOurXznhcIubOhwH/nv8Tte5TTy/
ekRwUt97OEdvm8AkbC5L4HyKJSxdRE9uqfUSZiccQo5HhxgakmIrcgJuN9rSsfpgeaccWs0phaen
TNm3tbKGHg/aBzyYWmUlzYUt7vzChaNIq23bpURCX1AFwYCr2UxlicfwlRHa4+o6S8oTguN8Y7VD
AayXvI5xw+0R8b1t7XwfZrOC0Ixd+The3+eq1hxRrUIp5CDGJiWGvQueXck08pF6F7WtTIUSd/HH
FfH2WLLTE6oOn7Nsj2yUvK4kAyXIi4caeeI8eGI+/zYrtALJcRQBzHigxDlP476szaB3u2YHz95N
rZB0NsA0VF3nqR7ZzbZ10KPdO9/05hrPzjiJvXGy8q3hWNHMEnJh655Zq8tZ9JewBYgBB7Vy5A7j
IGMZnVCGigrY5BWso5i4TEY/EXYHG0kxKchBNyofblToPSimPacJJMahjjj6wr2TbOojXB5jIVJG
98rTLg0KRJLPUjNcWfFw2rJQNJiieBwfp5EPS39d6aURTVtJ94KDM1QqIXrAUHU+ngX+m7lLBwaF
VE0A7xoaF0r3q+fn7nrcOmQvf4qqXPpI2BKyG0nmNjmkmeCfGb5r9pTQMD65wV5zHInzllQdDHZj
P0K6zlNvG6u6xNVcZTwSGv5zEhJKq992S6IpESo3/DlcU2nm2TWo5uDsL7dG72aOUESBYi7tCEX6
20a0g3nig+HxNpcoPbpoL79y5/B5C88pkVblW1QfL7s9d85zT6b9ETXE8mcokRROhbgyYz/TKW1F
vnPt2bfXhjOxaomHAt1WmI+RWAgYecsdTlKd3/BO/3ar1Pdf9Dig3zCHtbdNyyQoFMxffLTZUzKP
J3p5JV+jQWLcx191mLieGD9Gllmqk7COiscKYjl9bfbQEhrhlvNwB+WpUVZCVqBKV2hQsIPYdH6k
l4dJMWkk0Fvnzh5sw43Tsw33TOn8qYD3dX9CB8UUNb4At/IFMKYhCohzuZ7nMzyDgHtXtkRPm2mP
GZ9uoxhAXMcQutvCJkRUWqt5eBc20U+KA6HrhW+aOpExHqtRAlOvXiCiMl2cunWUqnn/BdsjxDxc
phgIvdKSAyACmiuobUbR8LF69QpI/lprSXbRGVxXPxCwq7xT20lEKXGrzMisWM3zk8GwcBr4Ms7L
q0thvKQcdgyAKwxZmfUr08+1Ub+589wlyZ7j95Xm6325hMEvYmHmfFKCJPHeuGVXqme2KyUexSmI
gV3c/DJd31c3zAJVCTdEh4Juf/KKbw+QaygLSlDCDUS4s356LxpFu9NK9PdcMepmOCkA3Cfv9HSP
uNUDY9ycyUMAhEQ0YC+EAkzBU+xNiFVTffLRrDr6zEME6WYKl4oHv0V6PN6nEdLdn60iouhG2GQC
vMQJqeGfUSzp4F/QtUIyC6iIFngw0ZBxrmzk1KX+H4rk3dqCB4KoIes7iUBAEahKg989LueA4lPK
gnDun1KDr/cLZODK8WJMpsaHtBnxtvKjJa8EPEu303Qhu3RQQHjpeMSqHY8j333EbMaWF4fF/LCN
3OKo36Vrd0OxzQRRRuN4zJfNtrwIGOJIqewBwMvbszSr3gvEl2pddETMNFKlysh+qnNRVkEUKwrf
OyGvY7oZMQ5YXG7T2qpYNPYLvgSQO176BodiIYptLuZLZVC/kCcJn5xoX7U1EEeXTmZOgYNTnkjy
LxmmfAghuwt0671J6VtFH2eXp3Tfk/+SchD0tq9UoudIPa9m/3jae42WTrOs4Vo4Eqzj+2w72+xX
Lmb6epgpx7HQ42TYaocto4EvJMAl20Yij1HafY6aI2jGfx6Pic1f4ZmWS4woP/z+vPciBsrh/fJ7
Qhd8/5TMmXcfZPZahZoTk2fjsEzoUN2bE35qJWHi07JyhZCsIkhOxQOO50XeT9p0Nfkiq4uF9nSu
N4dSGA4tTwdE+9zPcPFlzJVFMg7GXdjsEtM1gXtMBKnthA3cbtVfQ1Xge+GkOHIwvV+sfFbXJw2L
yId3Osa0xyfeZs7hJGQIceyiBaa6/wDci57IkbYGU90vsoq2pq/Nefaatqj6e2fdxevq/SYejpuW
CvlbjeKrBpn+a4R1duc4723GhYmUMoE0Q6UCpY2uMvJDiSABa7QlpapMg1HTzgbWPD437aDSoFHl
/umOXQAG0UgoJxNKJJERhhjRrIgTswNCpTRiG9ahJvB62NPjzjdEthPmAcu89s8EHGBvJkUg1A4T
4ym7VyOWDwzu+hS9dRPsz7ivIBlnsuVh2EMtOlJxD0GkIzzEGrjIG2jTgXpMsFetTVdxy8oXFa8c
eLyIMGMg0/tv0Jhg0onkKN5GIhkFcQAnjB5t6Ya6DK3sL3ghfOwFGl7Cbjn1KFVgT20Fk/gnMh+5
C6kVeJSPNCbEPpl8laEOc7b+8rBaagYrEawwI6fsun2BjUXYNqXohVXHUJGcPw6dUdWAe96PzhoY
zQx92t9c0P63S08hQx2+p+uFB4m+VDsY12BNdYL4khd+ye4arh2QJdj3YLnBFsEr8URCGhCZwGzT
4GICxnTLxI94Bszru9xFwrXztf5wDVF8A53cAG7K47u0iDtzb7htLo7H5YT3p9y5RKgooDutXem6
g8WmiQdvksHIZYy3ZF+vOFWV537jM6SLgdgGykXvmK6hvscviZsfuYxljhW0J0n1qKsVVyfwxApO
sR9/AVmd3tModg9UQfYk32MMO2GpT3/zgO3pxQricMr5m+1IbnEEuTl939RoxG0vTtomHL2IkK/f
UgfIaHviRqawN+E9xzgQyEq8GsphGv0SS3uZtEGac47Nx7BubsBPF+x/KdnXieREYH24QxQVWrGq
jR50W+AlQV2jlPw+iyiKylrVCy6WlOJi04Vapy0/8151t8e7PNb7Zx2Kq+IZZnORgepO0dzaR2bl
WKrPrVJAX4wCSVHW4L387h5ihlwUKA/c1Phdhg1GXYozRWTP2QbI1bz4e6fgKegETR4bpBGIEXs+
WzLHfyPo1fKL04lrvAp2m7wCrxuLffs9rdIyEPMk84iB+GTgVGCCIb4Ysjlzzgt11g2c7nZyA4Ai
Da6eTdxRTr2oRMjTHFy7D9/SJNAhqoS4e1TV+FRV1m1MKDJk37ritcuvu+Sdoxo2iIhzwKM0E98R
xxBvYrXV504wQwTj5fzSnt6uyh3EbiV3ZUUp8aHYiu43mdcXMnBDyuZVfKxbAklImTFNWOzF7RrS
Kqq88zeBJZj9Sm53+LDKXHW/6807QPDLK9MfuWjHu35B5o2dRV7E2mrSImOdifX0laT/bxB6cOke
AI9wvwXRRDY552qIy4XkcnFZ9qaMeKAwGM5Vbn6pecypyMmdYn631nVoffq4HMO3+2rt8+vRa7SV
wjvGvhvHRPhh7QGLzGgtZ81rkYYZ47ouZ5sVMI4Byso4m+3+2JgwRCVAGxtoZ9Ct8yDFpkXqwyTy
Necpvm03jbatcgII5A60t4XuihtydJZ62cDdgNYmBCNEmHKS+HZn2fpYECK/5Mhb0XdTH6PHTasa
Invm24FMnHBZEjBcm+gikJotcnlskRp+jafIrb6D5NVaqvqJXXXNKHiRh9mkw0xs67am7VbeBfzS
mnlu0zjSUIOxbqjndOFQfzXlZVWg7p3z+6KlHeQEvBy6sqS4MA5iU3cOIm247oE+0JvUGwyFfOPl
s41ik9MCKcYW3fi5S5FR5Tlh+CResoTtH6lnWzaIY4dPGH1bjj+p/ZSjnh08p7Y2kLHiceQgMCzC
kGGD9aAa6OC+xZVwbdwTX1nSrHrsJvzSDa4xEksTpJ/pY/qbM2bk8vxvq2PWLycM7E4G0n+V1jMg
b1Zf08e0GbTCHcnxZkCjr4jGHqTq3Jfbr2AK2cVIRsecHA54HR6dQdlD2WWu05kob/LD5MDbswhN
ra0WssNZmPuofzG59fN0+SyKr9IEaLXI8pm4wb0zyydh/TDthH/LaFH+MkWhpkQ6XBpYqG3L4n6R
ASO8NFe/f2RjZqVyacFagdjNGUrWDxcqQki91dOswlZVgHJP+ex8+Whnl9Jn1giB+DcUTEEeSuFs
gwGxeQan/LAzmhXlXH3HPkdqbsS6r4bvKJthqm/Q7Va/m+/Bg+O8Valn1NL6uPfmbyLYit4xZHtv
vMgs3TUbyKFm85kp0WhhihpDymlGQcGeY6BEoIRKCukFa4fMxaYSjxVhEe8cEijWf/xnzNfTGblR
EDDNh9CqikH6nI/CWv9qbMqDdl1FtyUXawJHLDoavLfbZZYUDrdzPhdyE5Y81dOsxu4tcerSdZzC
OL/NY4B03yIDe7h4TkqV/9jNKVSl8388GLTNSrooBuh/7135szBJOHF0HjQL37eLBveqB+uTvD/A
jxbpZQfUAq1tdCFnOgptOBzg0qX7FHXT6jeUxF/5Q3YbGyeOG8+OEXxgmOQja4EjeGgtT+8qOcPS
jHpMHhU7nkz/svNVCR1lfB/y7lBROP1i0r/iUum9R0z7zpM0jhr1/RvtewzRPhH0+UbKIMJvJpGr
fN8FaqFaOlmyNpN8ZFfNwoRaFfpp3AxJqK4+XyEX/uznrbF6ADwO0Mgivu9ObWBVQGazh7/BI1Qt
RMoQqWplu7vEsj7Z/jSfXjnaxgzJG9Za5F0H+NOupeMuTIIL3aoR204TVNOiEcqLS6nFUBU9hxKu
6IJV7vmmWnsPtW0LoGZK7D8T/oqRUlsf8q8UjACK0RlE5taFxPD/+2ORAGsu1HeXngLwgf6lEHCO
da3OTscCBx8fuo22rAzGDylHr/b+3t+/bL/0Ln4dfw6zcWyumCf0rc/+5K/SAe2sQZHbKffVvOv6
O80+CfV7RhVfrh4hy3+0o63Q7jmg2dEAPXd7g/6L0wCWDeW7cxI0EaoRP1s6JpVd44MAUNA5OwWn
Zjgz+H587Qp/3qX6hi07QlDK8o/Wfap5F4+QifxJi/EG4FHVPlfBRHhoYTldkOaLgIDzU0yooG3t
aBODsQgwYgGcqriCi6HB/lPFLcS57mV3ZfOV2F44Gnm4x/onWee6xP0BdUjZ1e1946M3SAS9R3Vn
iI6vjiDDiF16olLi0c5g0Iv8jH+RALXMgKHGgJwe1gU0E6VrGCcyISkozZPspCMDJBSHiEwA9H3h
BO6gS2n2Om1RuD9ePO/0w5NCsnJBC7tAhzXa41nllTQtm+qQM0R5QfAKgkYTmZO2T2+V9RoKiWn/
qExFI74SIvmYLrRCax1d19UAHF5DozLkrSykj9Ns3XwtiTodIL5QLIlhzWOo9TVEeXEM43Q5SUH1
Qv85x1aPQle1sLU6N3b2Eh+DVN9xL3O5v70l+K9X8eRkNgtut1XDQe9yrWKe7hX70pYlFg9iIEVD
lERoOW4KcTVaEN5/HxxPQWBWr9jkgC5/uvqjN1HLz7iwo102iy011rPZv3UvjZvbZMXPnaiS4yFR
bOBNIpo6XzGMz7EuPTAcdEGbiaaGmJDVQmua28JdWe9Z6svA2A99n0OrARMhXsfb5If5PQ+3btWa
c3U8W8kop97wu8WL6k1qSQqYCaMmbjebqXTSLwE2vSkWQdeMNF9+lKYacoDrz8fu1xxp2pApBz9T
sNXELgp1sZWLbKxAkrQfwmdBvHzHLnEpaoBrrzTnJr/LoUlcscX7GgD85TT+ECST6pqceUwBP15G
2kuZCQ+O11m/8lhlKNAmUHz5CNAEww8XDavZo6hdS1cPBTaajTAVQbonluG5Cz2mb/s6F231N9nY
k7gRsxNfrXQXhn6rDcllPuDSYnPWYST3wu0cFGMrklzFfZ2qfWOq/eCDwdXb5RX3F83C3H1KSxOm
wV7r6aD5r1eR8fNAmCLBb3MIvwT0ob8nH69rkItnyxeNhcfTu0HvNa88XlFE4rzcb3Sjs9ZVMU63
SQdbiPZvqEcmVHBjgDT4Sw4jNpYjRtK0xcG43mRO0FzbgN5vPrxYK4YUK3UtkTdsCN/jMXy+5BZC
BxScR8fd6XQJ/cOKejFc1J+dtg344FYEog3ZjZ+iAz/Tc7oZwryCsMnogDad4PkUPpuGgeIaFuvB
fEIIQBGUNhvEpMu76GENLV1WmISOkv7M2hl2ij35r2WYMoHFpsJ/pBIhQqNQv4r/DSeYM0AyhmTH
5ujnI8psI03hBYSQE+Ny2Pd6hiPL1pN5ZfWz8cpYRatZWvLPSRM/xLMs5Q2M+K7OIpoeqE6G45IG
rpvhGTYDtSHxbdaEKlbHWIkvlV73EenPu6hvbImtxLCHrcYeupGU9o2CUTQ4cSqEMIg97qbvVGmM
d1MnjY63QzbjzrruEm8veHKWVc0rSt4P1QUKUzuvUnsuQuRHBi0hYuU43Oe9Hmozf4JCpAgumfLG
DwOoHP332291iDTVSUay+UYUdvuZnnK8xc9+RcBuBirlC2o/b2naNb2R2cidSdmhDxJ4rEdLGS5T
Qffo5WExztGmKm0qr4nXwgVbbMl3MkbkCagKihP7hedXo8/m43h/QeQBJe9lWWfB3ZTLt3sTy6xE
IX7hw7QeanP+fT7HwW2sUXUfzhI0ILMl+1P0OZc7xogPeNGMi4OlULcOcr/8w88vyMagqY6sALGx
QgcGoFW2VFV3itwEENkxo2CbPfUqWUUPk3c0lq73iWmqkumbDm0NrQx6ReqRCyran4xOmfvzAOS6
zyP2bKqZh7p6pLZHXvcFg37MlswSJJmKgMAz0IpTzE62yx5YmTT4EVJ1Bu8I3o22Eufa1DG14bXT
ehQy80iv8NVXykvEMvdikedV0PFacCitDpbMG32bKIXfDlRSAloLhh7owhd3Dvcb1yqi9h5ZAXbA
FpBVutvzkMTUZxlZFrO5HTW01FFLt94b3riOkLQ0+E82ihmi0GwqFFb5Yj+qX6HoN8LZnjrIrEp0
yCJANIWPv09hLQX1kgwAEUCRJ5WNx4v8qJtxyu+DdTWE5XRi8ZcEyNxqTDfRlIwBc5YXQAjogddn
PtQ1Haq/K0bjAS6jDMvBKicXDJBgp/GaCz8Pd1PsRYNKO+mm5I1uT9pQNCVxc0gEhXuiD3bzZ+30
OtN3aSnVezuAXnLvJOvhugLZDSDuZ6DXmycrH7hK5jCaLJksXlYkfJrZDixhlJfZQcl9O1ggTiY8
Vc+1BHjAoLhO8/WEF2NVWzAbPtRjGLY5obrpgZ8VDBHUyBA+8K6lq/KXq0zv2u0MQAtlJZesv5No
jigmDlKl5jQbW9Qe3B0X4ePT5sGiqYxBq+GaMtNf39XS7ZVbLALkOMQ63MY1CQYxBmVxqSSEUJJ3
jIIKDvrJCvgAHqvHBR10AB0cXpj/5ovY6kKALruH/w/Z8QcSJhU968cc5ZUzzHVq8zqmGWWE5BPM
mDK0k2xHcdDB57ElqudmeitzenAHpJVyoggq4Tdckad5DeEJTHN/mrK2Q7ge+ZuG4SYr7Ngf1YCZ
1ZycwxQilQlqCLhDlx7lrUTUcv93lQmMEzYeUf61r99ib4Fwo/wg6mj560PFqK+uP2MEHoXFnOVH
jWTIXBkwRIwI/E+eEen+uppHJ2JK3tNGapaoFHkHXJwbJiUBoGR1ncnB2mdJ49sqkKtpE7bupSFU
5oKTR+oD7xnJoO3pLe2N+/iOBF60r0LoM/u7oQ1wBGpxx86T+ipGWIYdwcUMu+z9r+jzMcfWILoT
H7MagFpJtn8DHzWawIEUwuB2XJoPwJpF1XvVKFUTbN3o61kQxXgbzO1UzDkND37LtA0ljxafbrcY
dyYiB2aR0/2t8gY6tU/u+wsWY0dEH62LeGJ4ODmHcSbfTgUKEqAdXBy1bUvcLc2qPYgkm3hWn5kE
Dk+jNOz4ijySiWSAoCl/uNzwj3FzWpO0F3ZJ0dGg4Uxf2ITcGTlzpe9KNnp/TkRYjZML5r/jYZkt
PEBna7rIdJ3Wv/PABP6QGwopYLn4NeP14GE7BwCG3KpKp4mHtFQ2CgX4wcOLMEFyUTDU5Q5FgdO6
5/VecEyQ4jySHfJk7c5XN7g47FSLpNNbYjFSlADZZcIQsb06hbFMtSMCwHnRw4WcR722llEt1gGh
GzeRaOPUoU5clJVXI94MQBraT9UrKTSRWdJwYriAfW6A9N5+fm1TxHbSpn/o/lPVxCTSKejKwG4k
VqwMbU28sqmnsoYw3A8MLW0+VXN5CWq2fauW7i19GxCrlASu9wsXm9bXf6b3CKxwsn/KTTESJte3
BmGdjdlf8fhkqMPbYw8s4WUG3avrw3Szt5hWO+oqCqQ8rbI5qpOgiQKq2HTQGvU4O59VC3Hyf2uG
EHqy3L27oeC6CG+SoGYisjFqG5ZLpmgHLvUTdxrGIar3KXOh4xQvkbGa1uOBOIjmARKbdcGPxnLg
WcQa3zuvV9IB0PI8j3oSYwpAKDY17/G0mvJVrUZigPFK2aMfKgFkyLpfWIu2P/J3uVQkQlyXshbB
BLI6PQwzPW3817EEc+9RdXftCHerP6gTKJtG30aXjdqxwOsDiKIeMJw2UO7Ht+1f5938kQH+TU0K
I+g9wZhAg3vXcPnAf5mfzBC8FWBR5VmZ41jgSrM6Zx+hIdp/D1z/BXedXFVEElEnTjvAt5sh0O4o
q7HYcyej5eyNA+UDRhgzBoEA6teVTBTNoGpzbvYAOPugBEpZrHEiOa0PoALPgWi04k36yq5cabRP
RNJJOy1WKHktGb6uzm66dLkuzIbevgZyWV9usi9UGOqduwwbF8xxiCsR8/bSlmAmlI+oXRdQ6iEi
2LG7MT9rdGZp+JtC3fYPPebkUKwIPuN4bDVB8r+UZ3L7F6y5a9+cto6upCoBAh/72Oq21QkVxaHC
WUoDctKBn4mf8EYy8Ypn3v/h0Im5cycU17UokwurGqCKzLZXqCywx1GOi3AsSWA9YU9TIgAyEoU9
Ey7u9qf88v23zeanJo2CbURB4tshhmjPjfdLfclczhKPhvVlxpmGUKlHCm96EWVlnaSjMgrwuywT
YHHOMLxn0ytwzV3GJomnzHYtYGQzelLVXJFeK649NMpmukuAndiNyMaVQesIvUOuNEnoCeN6bf5x
jWyppwsQIwP394F4Gc06UXNAX1bt5MX0n7DejLoUJ567HFZoIPYGkxrGZyDt83vwzgvo83y+4D6/
+DkbM2YVm5SFne9+QrpAerwI8en5NwEuW5KCakmPKgt/k5/pu3INUDgGl4Bms7qxLc2UhJOoyOFk
tqxX0A9Y4l0eyfr3iJaKvJrdD8UITYDZFOGfJe//wbvJrw7mDlIMd9O8ETc40RI9mg+NVAqoaU6/
i7v/bGHlaqSBU8Jp/aLJdZzvnGxTzeXkdjDSi9OX4pP7HHILw4de4A460VuqBEQuGy6o1Rjc/VuG
BP6fKEdHNMKUfEuknqxayiSquLzjrx6aS4jAgovalq1g+G4ZpeZB3aiqtUHVmDXOFNWh4PS9a4BX
IBORuwBGL3O9/HNhzYn8dcNkfBXnkFfpTHB154UqCtXz/4x62zmkDkm6iyQCpZlaMzYS74Gs6q2S
TlD4AvOU74NUleoxfAFw5oTS4Qeq6k+Go03FGcKPdOIYLTfkFpDvhEsI2ybwd5TMxhSskU5cmRhh
5ZpFr4U/L3in3Zn2Si/XChuWQVsVVOYV52TvDLJXJZBs9oAuC6S4Mfz8ymqJDHXL9BeUQoDAsrMm
RWcj/37h2n8AFj27p/e7+4TqZlt37+dCEJ2n6kPGEiys2500xdNc8bWTRuQC1boMTP4Xjo5tnWCc
1y5keY0s3rmm7sWC4O7qknBVx31spQrPu5W/crVHutYUEssXCsCLfgI9EM7u/q4IIV2j/LAo16o8
iK2BVhds1V7ijApjIx/HYCNJeGBl3qZt16qs6qhRJRlWaB6TxL/KpAguFCpj0ZH9W/qWlVuJ8Ljo
8BvUmsa5XtDp5fRQhFfRE2WVtRvHh1GJo6kMR0XowCeqmWZWDJSWEztBEaI0eTNY2b7y58WJo7ot
5+LWGGepoJ3k2tdGQRAWMaCYbQUXC18dOMkI8123qHfzcc7VaixBjDQcdgsKQjNsy7xbVN0Vh9DY
5Liv5/HY1l3MCFFAFhxtYO+gQeLnQSXb9BBYo4P7TdhzG2Ocgu8jwne5e+qJPJMK45bSH1Xi3aJK
KgrSN/ggMRQYkBqc+ckeWaG9B+pMVZFwKfE0S6idhqkljrBN4Lajalwzjlbsv/mfI7LV0lZxlQ87
y2au8npDkZZVzU9tdLm8CqWyI67JuPXfdnYBO5VUm8FN1+oTEQFJJ2TSgq5DviMK8/B+WI1dKdXw
iXgvYPU9fnMZln2v9ycLZ9dyl6cFBCGp6KkhK4NpRxiYvFfgp/wHqv8PHpset/hFCtJ3GXllXrmk
fbz/7eiKDo2cFaxxDNceMI6eyqqyrvLT0QI7jmpHmbD9oOsW0W0rY6sXzDrZ59sDyw+sxj7QVn18
n0MabaSIcL0iXzE0bUZ2rr1WksvPJCjH2p1ydBEOLabmwiY1kCEwhgIF+NZzgbVEe7BOTmTP7SY1
MSSk+b4SVDakb7nTLY9KZDOub1HRPH+JGb/xJNm8Gbxj17c2vsZZl0YgIeKDpxRlRMDTs5J9oOWT
bWYk6qC8pOPmwF6r/uZ93pMgMsSQzzNz/eH6D4vWp/LMi7B8ceXclHlonvaBKSyZ8NCJ5RdLScbX
v/ZvqvUNIg68DNRXYTxiwCbzKJqYgfSn9HOYhL2wTpJd6/v8Wd/aX9c7uFPCVMh/ORIaeybfjz9n
7Hq/+VAqonFb7G8SE+s0JSGWUMecy2sj5r+2VVu2QDtKx95pUf2wUA2vZWN1FC9AiFCAwnT/TRJ3
9aOuGOeXRvhForhVEtH0xerxowt7qwuPJh1Z5FfogSKf/YhSVRcB923R1qHKmRRvksZKZ35vgj1X
DI+QrYDpkix2sFKbIqZV0u4I7rS4PCOyxdsAz9g4cVsjwk2Eq3qxcKc6d9dpSBy9VZ9kxHrRNXxW
FRYJBEKG0voGlaNe2AwxcKVBEJYCCZktUNwcGilaZFOi9Y7LQn7wMaw7h6CZgAw9eL8UVFMGoKzZ
fV3svfhmoqBHcziN0nMkOK2cRhtWH1gamUZ5cFoN6wgMUUc0bpMTi12UVqW7c5U5Ml2HZ7HkcInZ
O4poWE6BE+U9C7JPtFh2bc2kyCb0wTlOfmHJrtl0SK7K1SAOIaOQINbAFPnWAsVaWMtIX8zx17yy
82EBJl38UVHr8705pA6/NEqKmCPmg/Y3UxJ/g0Aos/WI6lImCPmSuEhfuPA17NG2cdBl8D2PxSMq
1LSMMj4DbQz/dGVns87LjMb90Q0JoakTzwRQi/nqRde4mYoB9Ug+tZAZWuaANcKehbEq0iU/eSM6
q1vGFSn8qUrlgedYpm25ZpKa/n/mPt1YKn0B59D9O1sHAXR8p/50Jjqrr+qfRfKgMhQXKeGrTxzs
sp9rTKQ2cjU9G3+4hsQG++MIwo010+3FZc8pYRM36ztmawF3XTHPDYCL5wrUFiw+r6usut9RujoS
pYzlUcLmTuZ9drORnW+WZjS3du0Xd4rUdDaqY0Jyer03clcqUt+DfxwAdEZwxSo2wg7U0yrl4Pcq
jnGMUdjeP1hq36fLK4s/kXZRUa4Rb+cE38AQtvYnxEDcB7Kcieb6YM31j0AYgzIEd2r4FpnKD5d+
ouOtApajsRJZiWc4/LDbDk1J0OYUzAxCbc9X87wEXRh8Vm6NLNsn4bLVkEcIeqYGpcj6XtkrhTM6
Bqoqt28oYuHeA37NMaULkKhG0deQcsqTOHVUadrvVLLbfGenzaKrkO0toIOu4KgU6YcIt8J0+aiO
RiaxT6fhPsuMM0UMUTQX9rBaKs+QmVJlaGGwFFXbNleOJNCXfoCGZYZzwBq25+607Xudm3IFCIP7
q/VNT8jt4K+YEs233EVEE0w0ClTE56l4tsR0i+scqF49Jz3KWLNEcLhl527Uz9fio/yU7JfBwmOb
BAGlsWrgMk8NxnXXIq5UsfER9/TCokGn/HnKRe8549lHb4hifk5TyNBFby25hMCtAvEexd/pOec+
wTYj5FEbYZ93uDRg6aVUTGX5agwEtmVvkvORXlazkrSz9p5+ux1tY+BGUbRnCZ6lKC/q82hC0W+X
bZnnwqCsyHfr1GIH7zFr00zRHDQAKRAvdO7MT58uo6nfL0K9VBZYdXsoGjib4u/k0+/AdJ97CLHw
hquMnrkqoZjbPRg/QAEL7F7vFz0obz1BVMFukMqsSr+//4cyGoA8zebihWNa7Z/3IKkcFwKQkj/x
gmx63jdKvlZEs4gYURwQBCFZLbTWavQ/BWuSyfBgdFnwqlT1xjaS92kLKyOY3pm4EbnEUJAapyHg
XeF+dP5Buu8feG5kHqkI89LpI85hQ72WaW4X+orvclrh7C/dlvlj0EvULrYSqxY7GkuIP8ijinHp
rA/fMYybdjLqWyJgk5Be2g6qFe2SdXqCcigsM8WzkAGY6wUi7PXIlWnlgL3rDayKaBOnT390eQoP
Vtj+/s+quczWTx2FZH6nurEkN39nEPPkjBSOo4fvlHjgM32cqAA0A53hJ3dDL/HVjnGnJT4u0wEH
qng+vINXADPyT9k5hAWnUN1fSZvzY7X1OACr/sB63wleW9Z/7djky+nUvIfArYyY1JsXugOZDfHe
FZbQMI7qdG1hpfbvslRm1ecy+bNixCSFsfD0q6FzJcseFGMZbA1x3+ywuWZFA5iMfALcprHXpZAS
HJQXYczteucMZp8D/erdMWSJeetdkD94HYzdE3gNFMzKXmenKFRCciDEDyRglvPhXM/vicKR5jWX
9apKrk/wCH+SxY6X1AJI/ObKAS4IUG0QVsaZumsijnIMxFI1zecwEaKE4phOhs0FF1lSpv1Wem34
Bfj43AVtp1E8tdFKpZh8MHXn7Wdvsj3B4u6+ZUjYsp3tXMgu5LxCMaUDeVv4GqPNDxml62anrmIY
oulS0/7HSFUniAMzc+/lqjyg9aixxd2M72/YIdBV55BOevGRJtpiMEHu8hmoYb7wM0KvTkKmbcSO
FRnpRKdZAEX+VLZFS1HvriRwfEAjLRqJkK9JqEb3cSadSuBYb5haxcIQp5iI+462FB4IEazNAhTf
6B8JZYtvKiUwiR3Wa98cK6GtQocAb2EagKZVRqKkRKu0BqG1UOU2J0MX0JWFK53tg2G0fR2DCKB+
3outIQP740E4ypKOBE3UJvIW8EH5DtkMrOGOqqGfRv1oV1wAPWBIMLqDHQTIvJTpYSEeL6ikGs7Z
AgMHJ6qlxfKFHAMWip6cYE8/gEDP9EKwL2pLfziVJYwUuxGaPGSNxH+25zofDJq+rxVu9lcDNRXV
FSgP/qkR4cMTAf40UjDUS4emiH5iQWeQn027Wf78CPazWhLj4wDMMfplLuRk1tZQyft36YIazNkL
glk4FJiXPvq3RBCRhPyAy832p9YIvuuBibLBaFyrvuU+E4HuQbAvkXH3TOldZSNPO1i0ZPOBWaP5
4qHSx/Un+o7LRkjA8gPHd7LnuGyQypoqhK0f/heNpD9tF3HQ6hdErJ5+QXYAn3iHI+0LVamlOe2q
YYqiqAw0VVV9rPbNMutpAEeoX+FwcFhlGbMRTo2Ll8p4THo4bS1fCbp/Chd8OOtvvllTI8zMP/4R
S8zQXim7cOh20Etufiu0uekQcsCCp5QxJNXlV2o2ApF2USP5zjt2azjtUL8bkSkFNzikz10mlQz9
bYYrpmJ9JB9kyCsa/VG2rgRMpc9nVmVMO6t+LKKHjh+rCWh138y3e3h56nsy8GfIGLO9DG0BOLIA
xpumPeLTlc1rKn0x1T9kVA/Ijw3w4mUYNqfALx9L27lStAxlQeISReE+jQ0VTs/1m7SeQzJGU5O/
Fxj2+LtrAaZEfFtnj9z4b7FEhDH0mBzJmy0X0b4328/uEFavv+WUPfD3HbI+riMr8Yguasr+TLXQ
PW2j5bVWwkx4TUq02P/sEmrI/STuXqFrmTosgrPVOMrHdZxsa48UyXEbzkYEJtUqZovDdXn9iJeS
GihZ6NweLNXGZRpw2zF6dmdUsN6T1S6Pa899gIM8Vl7LhsIAL2r/akufKL+ykYBMV3WcYY8uAR2U
GWLDXt+djayLHDH3dmWQJ11CgkEMNM67aPluoG/M7jxWnUu47n+fn1Q+9Fd7dtKew/f19M4txjLg
ycKhs2NEsyVn3Pw6lDsv2CxkON/CQ5k3mfQn6lUqLDqNA4/RZs9667lSJv3UpIJ1QtUYKxYhSSbl
jR3kl04uL7zt/qqOXbfhg+y5/QkGCU/nuDqnp3HWJ/AQo9rPuEQdJ7kFERZFpcvUzrfgiku7Vtv0
3wUni3ae/nOH6UU1k+n80nPPTlZlz13Y/X4DxGBWsMLKP52jXqLnoTEYCprNfiGzy+ORXEhYYPhL
WiqIAhViKzqIb2hDQifi7lmwRlCrwUKciDqQC7b6YV5GBADO9m8udv1Sg+5pgYM56pRg6L587TYe
SiKV9wZDiMAwXZ4OKl1YCTl6gaiIOmOiWFgVpkKaYWkS/vl9GXHTpLVhh4A6cpGhfnBRDDfwqf4O
MpD4nohzJ/6Y7g0GVnkIwBdLeuIJgwTf6xCFulBLQ9KOfnup4OGppLs+8hBT5pJcNtIFDIEiU21x
1bbQGe0d5cL9FS4nXG5OzHEYWicl+iB007zPyqI/SurmRjJrU83Im0pEqjl5S6TA6h+M/Wqk1rJR
B2xsni1ITTW9SYS5M/sondskpU8+fhql5V+umbBCFJiaTCiURvlg+oz3+S5sb/ZiGrOu1YYzpKNB
CZeFLijuvUbpN2R2umv+ZAqkIYd/eucXwF+hwob+0qLLIMGmGFkHwpX9BUXUUb29u4+5Y7pNMokC
lhfLwv343TURSx8X/19Kc+gF206GLxGIcqlw7Wn6HK42zKN98mRZTMiZh4ISIWEUum6FYLIFOvEG
W/PAwqVHidqDBQuTMWFw2nWqGFNHzrxgyRbNLYjJIQiHxxlZG1xGgfmr1zyt3p9mItp/zvzXuxiC
1qNqJGzYwa4JlyymT23zIe/JcBo4ESmYHsAR4Y4ZC1aPmoR7D0OYsDKunviNrMI8tL5E6W+3yAfX
KlCAZCHxIStx6yIakbjE4qTxLuJdQS3iC1EPpIkh+ZQwLcbOiBuPrUc5NoYlFpvuZrmhBaulTAFD
Kzn/6IlXKtF73n+G/1t7YaLXWvC0qQjruNbZRoq5fyh0IyGnTzxuiZj43pJCWNoro0xjLLqCG2lR
9BWOVzb6XVVlw3JJQ+ob615UizsfIyqlCJQiXC9viKjHGcpsSWvGCzEVoYB+J0JTjbbxvQEG6jwZ
VIO9Yc505g1qn/Nn2o9e3J1lTgJgmq7p5VvfooonP7KTNQSGeVOVE7wxeXMxwn3BCXRHVTmU0MnP
ZuchhMlpG3NUIIQC8o35YKXo3wHuIn3xYCOnMKqXh/UBkKItJ46lOaK91x7Fnms4RepFOxopQEOE
JLAVVevPHs3oz5ltpCMsIvtQI7vE1nf2mPWL8sdG2sAy99ihSt3dTpvUIZAgbwih91qmnqsRUDxV
I0y9fWTIWjZ2SCCuUsdDD1SoPl4s6eTGxncIGQLQHdBYCJ8yh2C8e2cuUaTbAVPmlW3UTqLwzMtZ
MtlR3KS4++tn/AUlOhDQ+0WRqYzn7aUp/tyXv4zXo2B9UN657wvl0DGpaZOmRKF1JmeR2NR5+ztV
XTSsyw9HfM/SG/qEEawIfT0wK4eI1YflPmrT4aKcUH2Z0Oax1i6tLyUQ0Fu653znSADF0p5B6x5m
GkG9KmBJv14kGbCbk0fioa+6+0EZ/ulTSIcI7GFlWGD9ifMNXzv8wOBTsrlZGQZblkDNYi5fKau4
BP/L2xsW3hMc36+SJ8UdoiDuPH/bntUO0ex+q05lgo/lgUTXhgG7vNM6nCW89DTGGNZM6Yt/eIoi
KgRnuzyB4S/foCaQfeXFBaLIKBWZcQTGtoxZuKJwkmaVlUf0CbXAOafByOnlv0jNJAskEokfZb4v
6igFXVFZpB/cEZsa2kNzz90qjKH+4prk4eEJckpMuBU6eMaR1Dg658/JuLf2g3Q5OE/iO7HEJPYn
Oaf0nXqTR/81qjnHDFdkWzrVK5XHhNAhWLoPFWsEqkneWIMyhm7791sXqoA+lKhEeszRcabYxVZX
o7qVupM9J6VtA+0chQLq1BqliJn+lE7yk0akXTrf+s+KhxAcipAQEnDQgSLBtQWKzb6wT55ZyzhN
O5m2yJefk9lb6lq/6WHh2oTu65pkI5qMLwPc30+UOeysuMjjcTyVqqm/lgsq1UhoyhA1SKgsIoUr
J6q+sBiVAolIcl7a/xD81cayYgZkdAG2MMzsWoVnqK7HLQ7nix+g0ILw1d/UeUPmGBQqNnry2nF3
7GiIS3u5mtXoY1leeGU8VI7Lp+XLZXj4Zn8q/dFDrFBlwAQnGK7UCGVYzf9qeWSBZDx3JrAt9m7H
9k0U0G8ObSSP6bDOXd7rGFopvmQAMlGntXFtLbd3XBe+QJPwyvrngb6MRUFHFX5O0MG7XjcZMEuL
2ljIBcwkBRGYZ3c6fyGFmNl9zYkEdNgfZNLvcEQnN2mJ1G9fT9+50MEIpBMq/8J6+6MfrlsTixaH
lPGe49r4zjsuqDD96BRPkNV6gPmDq2b36cnC0Ndkjx3B/R36iAnRCvXekF+NetxkSzGE5LmtV5Au
NuEw/T9Mht/VfXvL6hzW1ZzPX8JL2/7GL7YnNhY6GyhkhUzg21YZCwP+Mp+vD+PDcBcJ6WVEi4iX
cuWU3ApSHctiQAJPNAs9eDmQG64G2wcxx/hwoqwm8lnsEnXtESgFaToRc/4ahRxowMxrVUJOtSZX
8tzxP34UV5aRR6OHiTIKRv8+nnHkWo6SeNtGhC8QCvsVyZSIGs7dMYdKUYnTWR+tn2WPYfcI39go
IHega+O2fn1sROrAQ1OYc4Djz9SJKAsATTH0wRWHY5ejuJbFefe7W/3/82pGSdCyFxSkNjQaXgHP
ZHeyRp3Pxj2wWaPU6fk5JAEgWXufE2N3hgxlF5fSSXaSFlqyX8XMDih3Ze5l7CynD00Ma1Fxbzid
vJL2FaAVIdATRi/wBvjb7eT/IEIBJUl5+AhVYArBaZHIDMczsZej8lZBPN5DxpZN3IqLJPTcBg0j
J7PBhpiPWr/Df2sMQjthgaXfuMDf1LWnjHoRRJ+HsUjAxpyR6+wahen7cpBbKTm30woaLqpHhoko
quWs/sBg4Hpa/9bTPufsDRw27zr7f3OOIIAdcyAgH8x191Ux9+1qhu3StPyqlXiDDgN08m5edDz2
REZA03beZDYAtGAecx9M4yx9zZWQ7zU6qchLt/pkgBp3rQryFBPfQ5Y1elBQt1IvlQLyT4XLf0+5
tRzxoEMkvr9pgqHgSu9+dTYyQ3zDbS9ASCAfTbPtAzN//z7XabhS243YNpSC2n43JV9A+Nik0YPB
GNYXw78kCnIBuqDscdGYhhHbB4mTRYvtWjErLzzGGYSlNcCxnS+OcygNUga1Q4x108htejfb8AoT
7ADaxI8NH83QA8HaxO9lFSHhViFDSzHr+FD5Uo+jTlyQRrCo4o7/H49IhK+D+jdaZaIFE2NutVcT
yJjvxFIQIET6+6rjqhhviuW2LPpIaVCipzEl8aaIvbKZZ+UUKH5QUIM4gF2bxpxeWxOdpWGjCoPQ
atZCmb9a0ayGk/M44PdFG5giRn2rA5zcovSGHGAAt5kaJu1D6IDDlq7yz5i1b+q7djLO/7cHIV7r
My44GkllyKwUme/asD8pXyKDj2uFTY9ruCDaKz/qjU1NEZfAsJsMP7kJfHALmZPQvm1eTLTWWiMR
vHKUQwhvvmTNPYatysrx2njRYc/fFXg5btiB1Te2LJHr93OoQRtWtJSlbtqoNxO//ux4Y7xhp35L
waZPasntoHEHlxLqqZug5pooCOY1F5cqltL947F0llr4PqnDyaTeuwW0KnLm6U9J1UVPT/WanwVK
/UpyapjPbDtkYHdBCeFSrgRZMWd7CGkwf4Odon2/flxGdLn9d2q+edkb2exQd6aTok3Omhx8/QND
QcLxjHEq+dGbI/ffCJhet/5CUzrjW3sIvvR9y8pR5pSzvW/suxoPQLw1SC1ae98YeZSCWqurvbPR
3p5PP4gjmzv4mxnvPO8RG6YzonhJduAleO7HVJTG8odXqG1GkW/4BGYFjWlbOuHIEmBaZRHiBGAc
ovGcICGibbrc3FNKPf0nnp4UgRFTqKcN8IHs+65L8MbyQQxKWlRziQuLb6eOjC+zqhZ7W8yVcDR3
UN0YvkEpzDrz5gUpspXh+pUlW7L0XUF8Trr/8jlo7Q+zZYC1W/YhqN5nD6oxZd2m6Vb7jbzdoWek
sdNodzECR5mRN2kTDksZC6Tf0BVjsVdZ0qiIl2qsxm0yjUPrHAsLEkH1v8BKWsA745L5PNjcSJJA
Asv/piYMPCQlOp/epAdAMdTOy0454xknTFho+AwfpAoLNq6R4oFlGJ3r1Ypv4Lde2KtOknmYFhte
+Fz71NKGbwu95xQw4KybF1ylN6v7ECFPxBmyF3BUoZC73OMolSyql5M6QI5De7aVGDLcdqDlirUi
n0CugRAl+gdxcy9eOVZRKuYCcJSNrA7+dAV4MOCJ49VMu7dawQyHXuGob04FHEXRSp81iw4LNE37
fVrXv8GEZkpw6CZYfPrzAtV1qo6evy/qqpaiZA7SNnrO30kgCI9wrCd31B+aLRX9VeyxN+b8WoTD
MhmgzjxyNF1namDE3bUhOVg7cMEDBNic672kGOv2mYp/j1pzmofTWYP+wS7rmO2Ipv+TEN1l6yuw
nmOyR9UwIdlMFbTfMNKsxz3y2/gCwP+lrwmM4/q2r51d/8u9uAHhqa8q6N49SNpRdbtUYrB2UCfN
7hHDgKnwGrcWhn8BXj84uz3iXvu55pVDI079AXBfGISZchYCpCJHw7V2NywpRLRc81T2eMQfIgni
pUBmgxKE26VOJydvMSDc3rLfmQTQ0ZZRcxqjrjLQM8jqZ9MVoUg3YwFXY9KaZaDLgeGCFxzN30dt
ZLpo+144oeX0K4MOHTR9eHroikCECkFqWyRrqKB9JTVVd/NF0eNRJJBvEh7GxSiaCaEesIgVW2C8
PtC6vW/VRDKuNW9mtwSaXy2fuFkzD88lC8aQ4YNo107DQUvvvasp48FbJlvmT55QFOiZRRVySJnQ
vJkdyeeIyMNMA2mYoa9YsH00n0v1EVq7pn1KKUfUCZP5/hOy4Zq+jtz57PBfIQfZUKBqx6dVyBBP
g4h/pzpGeNRA/5McV6wr7D7tDfpBiKPZRtHlq4oO7Nzepr6BsgQ2u950D3Rv3YseByfFXp7xYAou
uAVQDWQlrjzrN/JAuZJM9cnaL3njPRHWQIpHG2DQUcMbxD5kA/Bejg6FgBgKY9uGozKxX5owS2zX
EEYR2J5H+mRnGWk3GVx50s2qqIIWJOKujA1yUNe6XSB4VoAsPC9EM7PAOEBcCT39uCl52XKxEz3y
3N+dCCHZfHCE2kFgcY1ooKU2uSNynU78feDGezvP8epXAqzzNVRck9j8OX/kjCZdqvYb/0PG/xC4
xnYtaYax8TSj5NrJROtxlRNf/O+RpbpkE7iX0kGPW+7dTZc9jhlhnI27XWpvn9AVK/fMsMUvVnyy
5r6YlWiDiK8zM2+uZ27a28OLZRtFKZl1dAnjKqKGMOt5x2ZrCIgE+PIH8QvwMpHdBMloSG8LIQih
/i4HIZm94VGoABqh0SVJY9jq2bDzr7M2M2JZDTnPVpEL1Xj2X+YgnxkGCHuxAOi7I/q4/jJW+mn1
FnOsYRoabcA1H2RvwZF0DCbTRk8CAtnYuhhFy3ILpbNMhCSuHIqN7kiCKmb2d3cMHuZ2ptdgpFC9
4diQRuP64evwxFOVtCfiO1i8hk8XmtQogKfLpZmywdl8FlPRJEZlYqhfgLPqZ7Ssy4AQKMEFHsFa
VqkRxdCW3a027We67RdGBn6vp6aUYZNrTQxKPnc7MFqk9X9steUAXDiTyI4A6CTgbESvjd1mI4vG
UXn2EDOTsH+oCfScowEsT5WpXZ9nCrsKpdUJWh6+qiEC264HIGwjs2tP+R1kmAwCyV7Tk2LwJgz8
w394X4SwMISM8nJiby2gc3MtFBTcsp1aEwwFib1l1poyhLQpj5ckDESZI/Rx+uWjdv7PrXD+D/wx
kBhOaiiabn6yc++ZDv5/gaFDWYjgnZWszlJdsm8lIaqkaOFhRyrZzkD5fDEgcnbyIQEjibCxFCut
j0DDTiuqvQPFVXC85X5qFmwrA33oFr9djJPziXQFV6c5d6d/GjJJYvErefNFdTlVOrS0jjEWDldu
fKOXVV5lGp2c09xcg42ojts4v4/KXNCRLW/6ulgZMloYpxKfm9ATIMuIRf9xdeDnp2c6t2AMFafe
cBqNGi3La6l3uOZJlCxWGxcjkGRNEuqljQns5n4j/6qso3qqO/pZ5NLUxielMX9QVmXIDmAp1EdO
T9/11t4XJidhua4X3JYtA9Oe6lhFFCb7QCtdqODvXMToLB4+zNcD8jEDWwT7N0/Feem79T5qCWiR
wGRm2C1kXsp5N8oXHwVdyyEGdK3+8odm90sLYPFQqSQ7xD2NvWAW8EueKCWf95tfAhGrFN0oO8aZ
jlN9CDy/ercGmrwJEmXmGbC3NKcXVAoghFJxn6NqsshB+IiyebSPtcd/sg/TOiZcintwhLXuOC7K
kDWPg2549FrwfiMsl1fSXy2+8Fm6je8gmNvIXJPxSLaxY8ec8O4TjmpXwCobpfGzEZozAsYDV/zE
Y7QZ6PZBB6dKNJtTZkagb35axawLsvzXx2AQvO1OH704MJMLJ7m53qhuE1o/u9IwtTjyPTOszKvi
yKTl2vZ7/XONwL+5izFM7GksRyrKV6hcfub50wO7CkKMeup4Y9vSHzbAE+uPjx+GWkOYVR+6afD9
lEMR6qAVw5RQDEHqjRzvOQbRjuoMfe26grBkUIgVv7NnPHxoeGl/hLUC7CEQAx8ktZHf2/rVOnhd
To2srovmRkyE2VcKCY2BdNwOFc27xvhYzTIhKboKO2YI0hIiVz55A4PpwE94tIXrhyRb+YCGriZb
jjefKsu1XMJ13oFCB6hjBXiun7RYP03Ny7RnUE6HtIVX9wGM2apSiCiEHT5D5XfoG/k+UrHgipvX
eIZHyeNGP3eNc/z2U84V4RB6RQ76QW/B6/Z9C/lcizqIMQ7XnIoirGHsaCLcPlhnPNYeHGsLDDUP
rjcsC6skEv/BDoEoNtR0qJg1HkgzTmqTRHd+aQuLwjDr63ubMR02XBjcPKou5rksmi7imC11fR7W
1ym39ObYJFDo0t9GncIPYtXvGiYyeHnNnS4/srYGOrC5PTRhOkUGbC+qon766L2WbGgOlisZuyDe
tpQ6Z1Xx8ayXFHj1Onl5fx/h0LEU864yLNCva0T/7403lO1xMjCW/gwFNnQoL2O6kl6a6eAoB85K
mB6ocU9cW2rbidwDTHP2zYxmFNIIh4p4FiB8Jf9I5dxkwkqtEiIKkgXd10XjrEoImBnCmRtPDRJL
P8TQcZB9G0eKEXV+sMVd3vwhwbBav2uG6yyUOBZT3lhXvHfbLQapzK0jItw+v6qLmIFxHTOEMzBn
HqeTD/QrCKDxGDtdUeVjxaMxJN3/PPxzfcA/V9gJ3lUIczLYbOV+ITDsyyxdUsTmzIpTWaCjsx5A
eg8/bBk+LlUtAgL5lxB79kqFlHUoKXnfNYmtxMnUxdLAnLoOdmp1puwQBTXTknbWlCKojbp/qB53
vMG8zOXhmA7hHqU+hsiEEu8tgy0AG4ea2z7pToF4p688s4FfQqjfwttZj/ak/0J9yPmL3eoNS0bs
YZyjNw/GBDxYKhMUe6f3Ymsphw68xzQCGcZlAklkbJ4jBGPMG2i+19R2DXaa0QEOCLo/XPcQQqux
DtCWCvX5p6+61EK9fTm+qjwq9OMV9pwNuFGH9Yh0RNDiGuTt2f0BeATLJeu56NkgkKlmJhrMOg0f
redwp2Ji1WwQCvhApyAesDzTwqUJk/XE0BN0ciNSCTG+ns12+SMkKA1bpvW+gYh8s+sA7ihGbjps
2ytgMGYhAxsPYxfW2YjOX0sS+is/6H6T1babEVNl7PSlBbyi39AR6oERbOl6Kjlvef50bp1Vb/k0
CRGIuKeIS5sEoEW5EBosH9aai0MW3xyci/TY3EPRMPCCHzdcltALyHEDhkZLzrhRtEV8jIkQ5pbZ
fRv8eBoF83j7l1L1S4UBMb1qhClxM9cPi8tHfdXxTiCnBzzgZx1ailEfyp7ONaHMUdvgKS1lqDMo
TECJoe9m30bAAxJoqjX63Bk+t8K4/lQAmpBbBMkBJzl14ixWiDsa+vbjEQM4KqzwVjEge/dHpVOx
AbpJ7fAwOY80klv4pO0CJtkoHjqFeLI1dNaPdJ6WRBEcn1Z26OkXozMjtsU8KI2Oq0Ph4zJj9S9u
Fwa9pDwnhKj/O7cTRT1wx44umqw+9nk7Wl7bLJEsvXSod5I9zwUz39wjK4dCipNgIIEghd9/YrBJ
1zLuewTlXNEyG3knQ7SHAryi4R3SmGUKR1W/+MiY0BhisUf6X4MW7sYW6WaIP4d+cnKFSsqBaXKW
9Czx54yhRdpoQSpBQCpoejjP3Sqgg4KGuZknP2s4+QTgbU7V+PFQQvnRBQDehB5vo0ML/7kdIeTA
YrG8N/RSxIkA88wvtmaIKwYTVZJhiXm0AKIl+uuTTQ9digSB1PAKA9DQ3Ja9dCsLnnXazsChRVDM
5A36e4oHaHHudBywIbjwhIW1jApvaHGcw6ZossJHll/SRJOsVK392siACo7XdR4lZRKUmBqMpArL
1epQIIa+PG9hqz8FUldgCdNagOOknIdeYNrKx4puFV0aUyvxCV3FfhBhwyeCaZVWax10tj3iaw62
V9wN512Sc90oVX+q37dcORsM3Dj28xQjkBPzw/rsKl/ZFQg43o5NX7pZyBIpQlX+sbjIvWlcPG54
+I/qH1eZMlLh6of6XIDVwDOuruybmLSJbGSAGUIsvvB0iKW4vLwzruIkNrgU+kqAoyRBCM839YRq
p6ozNjzmeQMYvKKgrfYbybyUwTb6jb3Jk61W/Jyh0l/iRKVf++datNfkPU5O7f0Z56TvDUbOa9g8
525lwxKbtKIrxNmwKLinLdrmymKSSi0n3uRCQobRm0TlLKjiGbf/V/yr2DJb1X94xTiMFx1ATL5H
pvu2pUkfssGcgDOM7BdpErNkuX4e7dJWzqe6LflO9DgX3TqTZmbFw2VE4EJkR7c2lwcDFjV2BnyJ
xqH9q/6Samg1qvJpXWhu/XjOaHc6WpnKIPaSk64Sgu+fqGGmKiV9JMLNvTykANY6xQ1nF/CC80pk
F3aOiE/oCgSOJ7c3gfuTUQ2Thw/xpz7ZlzpG+rhZSs7OFXHfVLk9wt9M+9cuxuudiyTU+7aZw7V/
yrKq47FpQ0WlsFmFNCu/acafket8IdySOC76701vKIOsaoTLmDRABWPu5jHmykSk1Dms/eIM2vOa
HTA2ZHOYAD3pDhuUCCwe0R3PzUIRCMRx9Wojvjig+diXg6/1wSA7N+DSkGnxPmn1oyFfbk9HmT4T
oQvRu2Elsz5fDQMj5sD8KRIbebeWPYQznuoX3scA1aY9twCY54K0rjVjAgC0AB9zwKkqWmenFzG7
5nIpVSdJnxa02CsyHMU3PGI9mBYnEc7gnLxv2Y+QEbyPWhcynTGibKxSVJKX1eMbDS6ChE6nALxs
0+eWHl12m9FgWCvIal8vqaDsyERb83mJlwTnfuKRZrVfCg4ziEtf5nyZb83KrkvqbgiEr/x7b1bm
noHrzc9nX/vP56U/Xiui8fMZFsh0rckg0iFcK178WFbrYZiGPLJnYigVYjk0Qm9P5uDZCJOgAmWZ
e/KBwGmISDtKbgL6FikQ8CGpSiH3XOVC2Rx5E0CE4+drYWqlQwbSnAMJyk8ITWvbEfOPDATIscyx
UMWI/AO92HTD4GKXMkNXD1wnGcYFOKiWduIw/v6nTl6eehMDkxiSyfwcvYfOhgYSi2R0cvTmVTVt
wepo61DIf3UoUdLf8XFOPiiKHH0eRRF0JxmBe0ozFaMJsnICYei9g8mKM+pg11ILoJCUM2o3ZduA
ReCLIt2J+gNKKbZELvRURHLk/+wyHGRwMXBLnJTEJqZn/vHPqMr+ccRaMkAHFBK872iWyTJ6plMb
DXppF3ppFR8n7EsOID5Mkyv5N9AsJnPfPQ0TIWPo9ncq1MKqAsLMTfJHSVeGFDSdBK7oZlDxIWm7
7O7Q/booR7rFEfd9Pr5nHz/oXREB1gEKZmqViU7aI8Nhh3OV9/ede3hS37e/H4d8pbCqINw/bmjd
C2q+4FYjaNLpLj+qtK1d0lIZp4nvvjwGp8VLvKq7iuDgbv5m6FzLi09qCpYyQy1OKZ480E3zKoZL
Vf0wnlaIQLj40uIgozp776/372DOX6+knxd6XAk3x1kosHeFXHtBivjvEMYUX6J+Ql6r9UNEWhY6
Jdwjy7+4IylH1DbRLrrM9xbPZg8eQBeOWOkdmknn0QlkByXpFtaSaovgat2BP2r6kBd/2+qrpnFF
9rljpi/A+tRotomF+OkM5goY2AKvXjj/SNKgKnBjS40R85B0OEmTE+YjzjzUUMBy+ckwy1qdniTf
GQNKCuCqHbyzoVg2y0H3KRdR3Adt2SigkOw3WyY8UpWsGynnWb3jqVB5OGedpredLxlr/InoCDOO
Ev5w+ccQe7DntI+iO07m24p1qxPhGv0ZlO3AsOYMk+QUfVgmY297HDVeNQDhBfp/PWsxsW3ignPE
sI+ZTf4/SWxqp6lmkT9ioGx/rBsidoXVwRPPxKEoE/cgqb28gxnckMQOMLgjL5OgGZtLNUWX8Q7C
mKHOJRQ0uErcWXfKcrIOG4occAmcZvlTNETt3gKvcCt3LwQQyxgwGN7JBhkdJmAo2G9oAMkbYkjW
8opMPe5kLvkqa7Zj6Z27oElG2d7d4J8UGytapYc0v3nm4WmejtaAv07x3juRZoxxbvdFiAxVMm7H
h4+UdgSM8T7p8+hUH6tjDbi47AJDQvBus+N0CbV3/ZciDDtNca8D7x+PgqMdTWc+QSrvh4xx+itM
AxFQ9Tz2OWepgmPEJjGBfHLYEfp057KDiB1yMYo1zwCPysY0PMKufXqNUjtHLKVM1KPvbCiUuwJ5
CecJyZ6ti+bsjD9LFcFh0nLz5BF3UVtuKHR0sivHkD6GK1sICUP4MraEZJCbGQlG/0QjkkrgnFiI
NIEIqQWbDmWQ12qkacUMiZxMBdpuonMe+8iUpz4whyRePBK7wvJettX1K80UsPUKr1+8No9TPP1W
F+DoNaqmNh3cx2EgErtnbwqX/U6VqZNRPKWZiEWxc2y1K1E1NNohEoFSDrXB6yudaGqzh5dXO9TK
jrXMAfhXrAiUf8WH0LuBG60JMZw4OwSur1VBuf3gNwy1KLyakNWMrdgZ9xTG9GrHk1kdvJ864LNu
FdGz97B0IyBVgvqwnfPKgXhGLOU6nhgCIHFDZihzZkWWoL1TSkHqT/hU3lgeQq1iQE/wKnK1m+d1
htIjZiNKB80vkf571XkfUret2z76SQKs4QfJTfuiA+UzJETwZmsZkE0Ri1lgWiTAWWWcOndp/OBu
s1SUgib2yDRAX6Cw1CDtyhcJWXgfzCHGs/N6qa1cAjkj0bjqkVfpFERYjXT+gBI9b5DayOmMGe1L
2IrAbQeHuLexW3A6XWN5drpAcp3joFegJ5EMbRJxGkgcN/BuLtfK4cHzJFBK0xPGKA303DHxxlHS
t1jZizyM/TswdNAb33Lb34NaSI/+C38TYqvg7mYAYNWDQ2oU5VsrzjuTKSx/iwllWOjJ35apf2fx
mD5zjQXm6H2vC/sSh1zcTIujx3FOTG/dl3MQMr3PZJKroBbmPRN/zOFvg44mqqYaO+IZ18yxFcNO
X/reU17VaLNelJDYVDP6/gNwqruGgWToPj6t0rXQ0jBtnbiCgeI+MMwGbwFXY6C62N1zs8RLhdSU
X6P4DUV7pObaEQkgPn+2twaFb90hepbKH1/RkrB7rPhU4XXt0IZTMDXQmrA3tUnU1Szll9HzdwcQ
MwcaBYN17GftctkCmug3jfbIi1VRpoPvCeuDWE4yDfsmmpb5HaXUHt6u4qGFfdCO6BBLETZTYGgu
O8IWGR9YZb8wn3SMOp1en5kJHukKry39MLrG4J8QDuKTpa0lmRGL71Iwsfc4pfT+ydwsA88O1242
qcN042YkH58fFSkC/NY422npvNoFASk0xH1URf+JMbyWI7OmZAE1VxYw0AggKPD+cSI+o56dYmQW
tlThrdNTQ4ovLqmWKmVOkBK62PhZOXODaSIgIrpUkrxvJHlZJyfDgF+hkrFzRQ+sL7jStiKVWHLW
rBeGOysPejRVdtjRVlSZL7pNB1RfUiubyNyStGMdRrT/MoN+Jq4ra5HGgb8msyB3NhY8cCJDKCIu
pmcITkNGL+tnUOfUwXhjLQkUPTx5S06xcs3GX/Xqwko2JbPdZSQt2S7Hey/goTUze0nbEoWmN61y
+ZqKSIvJddzAXPXlmfPhkK12AFWsyRFzH+etL8r86UXfNXab8+mwfuT87zAbCWZnDMZtwi/sKIha
RsCKKFunqII97a65j4t1AD25fCYeMOGfJe3FWD03fGee0t9otNbX3GSG9SPET622PpA/AKdWCDNV
T6gTAwpNSjBxZTQuAQgPhTUuwynFgCSfrv6H8/jsg4+YMQyPHEijF19XpsUA948PWxPsmxNlScRV
S7GFYEkD32JMDjjZMSff5Kn+7EjhvsCRz3SoV7sxo62eRPfoU52vqY1FLON0kTME7qL2t6kI/lK7
3bUcXthFpChi4L5/OvoMbdK1L+3C2z43mflS51a+4yA3ZWLuL1whpoOzamMZU6czavo1xDgsVXep
v+h/9qAXnJSvMPI16y7CySUEwENv87pIBCzCS6onUO7ecK7rdssLG9jba6aucGHYEjVOi2AjUDH/
rKyoW0eWlsEVTshx5VTCVcyxHlQkVcsGaT4CYehStgXGKK2jG1RXvSZ2jPlITxAu9tL84IMnLMhE
iqE5x+ARJDp4slM4JV/gsD3EV5DVCHR/k/HrnAkx3tWJ3qpZb5b1Ot4/O53juMfnu+tXqawoDY/f
u0LJxcT+voo/UfrieIjDRPcdkap5toiSZ2v6mDs02GErRBYP4uXkVyMDXtzykwWUvlgNhqwkIDTc
500iHdz3r6oE/3f84Na2ZYNNku0Ods3LaedtpIcvqFynPED/HMYeIaZ+zDydK0F3BTl0x8mhmrVc
qyhb+GBzY2stiJccYcwOYzG9qrESpqbY4HFre6H5Uc7nf02tnjwAsw3zCpCA+6swt/h5zqxm4IDL
M+bnMPVPrwbNWjldCyYgHHsCs/11WyPm32wTXqazrObILgLCT2GEyquWj8CtUqfzzZDBk9pXp9IO
uGvD6wUgPkZeIZje6G/SD0aNeNbOI4iZHtn3Wr0zmlgPWwCkdVyDLPF+VWlTp77IK94Bu64KRnrK
xZdnJYG7sRo7yBSdTmsd3Nu0JuPXo+W6Vijf8pfCThZtkIYXvxlFoj/U0sYp+3DlXC/DCffRFtHy
HMFVvdycWeQQG2u5pryrT6f1xTMs8HruJu9IaHegh740WS2QNBDxyxilYh4Se3Dl4lOsykuC5wBy
CZDwWssJx+ehYnI+xDjfegmA5uZ+9RU8iEVbZP5u8KN4BzQBj3+xZpSvdAGWbkmStkoWD/8jKXYV
IQhypGGxmZx/A/OZm/nO/vWjtLDAc6OdQ+sPHfIXu5uTqcZk+G/eB4ST8M6nJhX3utASKJm2JbN6
dTx6yFiD11MYh1G2wQTKfB1MTTVEtum6uWY/2L9cckN6ovEANHjSSSCd054x9a9cvSejm/nGpbka
dfUDZ8bNgtKxhfCTqGncmABZUE8bU4E9FJMV1rfVE/BDjnevK4hQVfZETvl+7dcn/P9n6YfH5mWi
/vA04CkGTOFT1QFh+hlW93xOBDBbDD0gs5tEc0S+0SDRc2YTcatf9Mli3ZcLgABq+o4sF2kpq6DU
rQ1HNUNZUWU9m3Eg2wy1RG8lv9tyLo5Ky+VDi1UgvMICj3AM15ntSf4kqIjCIxuP57cuyq//9OlJ
p32aY0a0YH8uFpzTgKCDQb/18xMrYJdUTmtjFZBed7EnUswtEU/dO2rHfpeFbV0EDpMHuTB4d46y
N5ado+WtnJdL1KAoUZbJIVBWkqhK8/Krc8/rCitumyue5PCylapXV8IRUdM0f0vebnwJbow+TfPi
WlQ/X8TGfNbBSZGa1acHzZ5NRA2bxlcidFgIJZ50x38h92m7WuztGZxz7sr4KCUWxgmqUrUXx/vg
XDcBN00TQdDYuPGIw6Awxy0nXmIkmAeZ4T2c7v0JuUo9zZ9nCIYWTiPsYgB4wFU0WSbpmskS5lhL
N61XYYpYhx8Yyu52GVOkphLcy4J+NE3Anz+WZOXQGXdTlPr1FTF7ftK/rS/2aL4xo0liV/ldUSi+
iXpDo9T/c8viY3oMkZ8zd0Kco1EKS4tDbVPcD/Q2ZVAUz6tt2rxv1pRWo6m3wgRnh0wBkLONUrEZ
rNfZzRsCBXtX0eTfrlSWDU5i7vt3Ivvwb39ABYY5LJIv9q29bzsn2jyMGDIG1dI5Nl8z0mz255lb
M9ge2tFC1u8pIqj5tM0GCLBzMTWVo/kN3C/pRkDkmf/eXaXy8+ccL7D1h9Iz7F6PMZo2S0L4rXoO
RMOfBkA9/M3k1eZvOieMIBnkyoZO0W36gwmLLbWRt9wwl8rAKjjN2vPrrxNv5NDJoY3FYBppswuK
+9/u02x8ATH0MrvbA40D+goUKA5+bQv8+kLPRIHR5t4fCEHMCNFawuRa/gTMr9Ogl1K+a4s+1K4u
+RnN9TrDgtiypYJbPaN8gCvT7TLIZw4V7MrLpTKp6dcC8jziQNtAEkpK5T7YI8yZbLXVd+tltepw
DuOeeflnt5LpJb5dzR2372827b4lsLJEirVsront02O5ZwjLDxMwDjTCFPH3dmNvx8q5LCDhPH8O
ZRitGIpiJcqty0mRndRKdmWb0Jws7oTFlsMheONfBhIBTAa/sgMOAdLXNn2zeiJYs1qPP7tJ+6Yi
/zM0bbo3TfAyHSgjIBiba6dsfQdQDWEfm1eqaLMPr7aAVYci9ygbcLhMskLiDgmlVNbWpQXKROOg
E7ENQwaCk91ZDJhEQEqW8HQO8EiunoSx8leuhDEcdq/6HUR+2mLwMPdHa1g1lUWp7xdhLaSWULSg
lkNtq74JLhbrmPhpSc4fhXpK1B6354gF7AaISnVRF9MOnzvyNph4OZE/jlgktb04UnTT7ylAPFhF
zVnh1kqeND5IrIyZ1JuAyYMU0m8zVm/1ogH7/Kd86bScMGsKHFLgy0Uk05/mHbrFoNEP6T3rdGyn
Z3TyuXLTZ3j2fPlZljulV3kRngGqEdfb/anEqmt+8UlqxG5O+XI3N3jaQZvlK4p0TWHNBhCN5PT2
BQ1M5z4bkttZgfcN4eMQy5lOkefNLDL5G4WSkU3dykwIQM8GSo0qeoNwWQRmYCAa0jpzF4OEKEg/
VMSImE4XJ3firX0wpkzQ8L8cQV3aFL6e5IpMkKD/t+cxSMOCbD7f0kdHd39NWPAfFLgpTnN/QOzT
fPzpdrLA7N6vdsSf99MpjSBOztKsbdYukj0DhXji8+vK02Yema4W2eLS5KRkxM0y11irJX5FRkFR
b9kuS0Cp/WDdO5LmtdCrqvQGfBLij1N1+nBHR0wjmzKDOllOMYKvZX/z+vQA+SVwnIii/THCDgyU
h+os/I8X0svvxZxbMhlX9NWG5T2ZzA6aE4pX2TBfGNwCcmEg2Hde3PeKaSeukzRhqGUrfV/1P4ZS
yvbB8HXhyT+kRInQU0KH+ekyB7bFFg4ULYtbFp9gT4a7T+q7l2oehVuBj4NpPdqnrdhORtyjTcon
v6c+jOlAyGfpjqRn9xzls4dZIZSfq/b4LQy7hBQ2Dc2WVs6VwwRS+cXbmwA8aY8NHVJvS5XZbrly
fSFngIhAYtncTDA6kIuOqq5H8h6GVL/MF5yTN1XaGR/aAs1mdtncK2AZcZPH7arMSOm/mD5bMOaJ
+evbAjQEExHoqlULrugN95CpN5EDhp5CsTrKDOkjFBxjbISxgj3aLfvueAqzXsZcqRTPFPNeTbkE
PvFBh2AJ1rTVh/5UjXhviKSvz3RifzjZItp6Lg3icdFMCYQjgF9fXI25QH5srkPOJ6L1f5jW2uwU
rR2wiui4cW7evb4YRqIkfPXqMdddk0VictT1EK8jLp/tBsNm0AEMT2UFS0/vQ9mJaFNzJtfYESRH
wwRhYjzTwpBUNy7j+LWlevRg26oHM2D9eLBtXq3bYsqvlEnhYkChWihPJtsvp5QPIJfgEPSPjask
9RN5Eayz0KEYWHg1wvnigEyEahJivqNLD0O3PsqSELvLuZPuKAl4ZY5vSxlrmVURVZJ++kBkQjwa
TJsXVxGbRWq6LESKF9k3ad35+y+moXzgUXc0EdE8ATqfztg4i88S/AT0G5coiHjgGTsTqF8wvK/M
TgR21M/EoPL4QB5rXLrigcMxSwSZYAh0P6Bt73bOz29Jio4LLYsOkrOTk8aI3oz2tDu7Jag9Rr4x
37ahuoIzt51xk4RRBVbNSUhTd91BlNKfDPWW+eHmOoFyzNuSrde4rhuRlMIZ392LOIvYlXq97Fy1
+ahxd+AiZgZKQTTagppDdoJ+aTgTPRJSx/UIXi1NA5SPIw6ZPnsum1XThh/63hVXSu7WrmSP7MKd
ftmiKjjYQ2YDOz1g9a8wrCc5C2DvvIMemd4vZqVF6vjihyxCs08ClO7h+xy4R/hW/jW/dl+hCFQN
Sh2zW1CdsTvgeVSVjRX1rJHomqRojfom8j89l5kVIg/5O+Yha8Nyg4Tg5bHxADIcHL4z3w/9Lr81
u22GZ2n9CThIt97AkCMOWoEZjioLg5QFey22Iajj3Q0YFj03Q8gJ1HKgcvb+404v9qa79QLqpqdV
L8B+5YyA/uSD81pOpWyf4MX3KHanyZRGyuTdzd99WuDI7TjO0hhYtj023kkYX6IvSVJMjZzw4AV7
F4KgXMJHGJi2iMk8vTvU5hU32l4Yj+LeHY2Mk0ovtLEGUb3h9FyAh6uRh4vrNr+gJWBniXfDqQDe
3aXqxaNF2oaqBRyduXv+VJU6PPqXvLIvY/wXQ0gNdWnYp28814F8cuCsbWoflBmuz8G18AUGL4s9
BBOKiMPJbHF+RFeVYJbT4HcaHViR8ZVUj4DUP+kfl4KYJL0q5MYQrSyLy0tHIKnRSMpW7kJbr9xy
GllmaEUqAlkst3+178X8be4jyqSozHPm09Gsu8R1nu6T7daeNtMSnTGWnnVj2uMPF/STcXatwziF
FGkwGO8aa4+BQpwagvKJA/n3aM0TE5DvlE3E9x8No+fAZrq3OK5g88rVnBye7nww0RUmISGpxk70
t9th8JxUfsB21gU3elyP1KyMW3gu87tH/pAEjsqedSNPu4gC2z/QqU45aDuaUfPYjUunw5ouHOTC
Et5+GinI5WkK+8mfFNJFBpiTbTbNBYYpCFsimmvVf1jyvVEZbCcwvNfnsiAaO/aH7opMQoHCWYYe
cC40ip10UqW37Kw+54LnAxHZiFZN3OgtYPA+TGR3+d0szK14YI4CZaccadO94UaRzoUCeP2JUFJ5
9SkdxR4jZTsglD1Ls5kcfa5rkb+UybM9r59mJYafhpGZJ0GQTOmHmwHSr5MMqyQ3GdT0udku1rvk
1dlzp/yK7Be91VbOxONOhK6NLp2T9hIhqjtEAHMLGO/kgnEn2ICL51C2S0KnCKUqW5IVfFu+Aq0P
/HIL34srOHcwQIZ81zyADXIIBzPz9CdUTDl/KTd/ByewH1MiP2trG4bqQQ4EmQchYyGs1A4shOul
1XR10/tkpEXMWf2PKRCBfndL/kGbeMLHrvRH7in9WWtfDRMLEcEWlOWUBMiVvt6HqLthIwNTFdM6
0EjB/raQm44AFpoGKnX5DqZTTMqX7tqaAmySxjxzhNaeHBSCvSvhtaYDb5/3burG2dl8ZilH+NB5
meDWbe6g6NgG5kBK16pLZGlxfDdnpm2isoH9TqXIjudDtNVQsspAgZh3A1hgasTzzxcRajSdWWMT
3MggwK3/jeJsUFaoJVQXfraDmq8tCmfi1bQdj8sJafa0QlhGnEYKIvPeDKGK6rwCt6hbdjKiACJK
CbAFtqQtUWaj23voBw/fzkq3nu1C9RcHe1FHUrDmcZqLb7t259bWg9V94SQ1ID/Hsnwv64ihdNbj
qHWsKUuYMpcZEPhJt8jIOYfX83MrKr5UiNgb3u5ZV8k8fEw0Am+MsDX+K1KogaetBwkmCZDunKmx
n7Dk+fcPtH+FhZKQTpz1lQCOJAv+pI7kT8Vw2LqIbD8jdZF589i7aUh8UQSY1BPGm+9LJLcIgi1c
H3VQAAjopldmN3o/sO/mlvcVPQ10ibd+VZyCjfsF9pNU+f8709PcIYpNRAuBxC4tsmcWAchoFRdg
6sHugGclIiE/Gptt3xs5JVciaXT3YQNRcgOx0WtGjKl7AhDBW1yHtdceoosrjPtYfuSt9kcS7Pbo
jfFFe/BwUeWiPxO8GjTEQ66ep8KWBy/QCIxNLboAfYopxpegQAfBRVsm4qJMtSmfZCMEi1wL5iHX
MnNjPR+9HKE6g6ccKSvB7knnu5YIN0Zz5ju30DMTQhPTW3fF9gJkh+0wfG5mC1MYSVjzAuICtN8A
C3DUJmcp0rxJu+fcM+sxTNzobQnftQyjc2wlwiOXicc2FWYFlB4as5z7WdCsiWQAinGuIxVYcOai
nLh9fCabveFgkJAqAJS2IFmxg0QJmBm4Hw/V+55kC456do0PueFvkkQwptX6KbGLKLi2JWhYDSN+
aqlceA3xfop9N8O+P3Xc1rFKePdisl5l5XHQ0r/IHE5m2rHVRi5M0KEnRHE4K0gWcqkNFamip0ID
ohGGsNOFwXs0cs4ZgEGMsU3EngCbVYHOh7MfgstyRzrnuq1vHT/ZnGetu/6JlJn9pdFYyqnMTVO7
HrCWnwcyXVSIV6guGHiKngVl8IOgucPQUwlqiqw0fMirmelIGyO0nQgWGCGerXC7EjMd9Iq9mf0y
W8bL89QDE5AWj+wzwpd4LC2wayT33P5/EDBTRggCMlMJvrJFiJObfZ1VgMWQCdgp5WkxZuzpIN9Z
qAe5FjAZK2dzXfhHCaospzVzCZkn6oIgGiTOtecW6PFHEpYQ/t5fdWUsJwDm0+xNdzyGqNToS35h
1DdRy9YCUybitmIRkLS2jcjh3UbE9s1ESp9yJLPkbFUXFyPdNkgQBGhXMq5LA+vYC8ywb1Gata9g
1Esdf2pETQtAq8J1Ube8Ea0gAo/0F4P+XHYitssxa5wZBNjYt83w+hNrBNGqWiDEEDDElM5P9RNM
Nqs4PLDI7SigvdDFrcfUUo7n0rKifPNREg9dWM6ALnWznWzZq0IWScHm62bds01YIrC5hhMosuf+
StWPrnaXSrkWDBxnyQXxgK8sAr8cB/euv8DOm++S7+DCAYK7tMm+CgM/WICwfbjZVMccJAispSZM
nnJD9tYqw4fpLahRKeQmJ1zUad3l+onWlg6E1JxyNaFGqbNv1jeJXfpiq3fzo+/H3ws9PF/stt4K
td8eY1x0cukLIM1lDqrLrGnwE0sIbVTdNEVo2X6uGoEGR9xvp7FoHpWAo9r3pGKuytPGwFVuIv9a
e2EMI97s7PnqS4ubhU/LipvU6Tmv+ylzp9STP1iBSb93FEKJ3xMW45X1+3+HrC3cGpYuiklq/xb/
Nf9CzFh+B5s0pRSunVNrcwIsOxmV6bah+532LycEV6+nNkjHoyvST5i4Iyr2bDMUPPmZT/m+Bs5K
2dh8lPhx3X/jVlW6TzgEx/mwdAyvQ95L0hu9kqj2MEFYn83k0aDubcMRQXRJnAK3hwb3fc2+7L0Y
GB3yV5tOkTmCaKvm0mgD9b+t7ZsLm4AfP9L2kEcyWp97HKHrFpbvTS4UzfEHAjWggSl0/5japsWs
3rn4PpQ5SANeDgBTZqaXdbVjsVMq8XtaSztI2Tlpc6UFyeQyLmiIi/MAxXBoYY4ZLWef7bFfpKIT
d/8yhrC22xrRaG4smMc81z/khkgkWlxmWZFNmdafOROnWoZd0aXiWWzrLEq1OJxTAKRKsrAQ4ZdZ
GzdeJgqOlYHGlOE3XOfR8D3ky3HvH/tBNbQakqDUCvO5RJLG+JAdjInsZ5Z7BDiNwnhPsHzqbk5B
nks+h5pBxiVviDGxAW5WVtH2hnHKUspTS61LyloxzLxLJgOfdU6YdpKwkyDUq7psgHP4cRjIkES2
WTsQLcufJZJQ8IdlInqTmiHzcIDw1LhHzcq1sA6bDwFquIjh3HlCDy6kAmbRWJAOzOutdOalnFpZ
qd3PJMsNn7AVN6DN4xRoOGg0AnaY6JxnNA4/Gs/rHIM+bXhDivzOmjXPSxiR1iS/BxQx2Kp0W2LH
qRQybytqN6W9CHp8BQEsZRggFasH4blKMa88X4VWZchjMHh12KBDYRouLBP+92McnwqqWM7Hap3s
EyxHYqlav+CISA6hWrmCWU5s+Xi3s1ZUxmBVKVuNQMoIqe8SV1+dmtkb+Sm7LDZV6zz+jzez/idT
JqApAuIB1Rm308o3cmKjfOaLXLURYum2GDoEAJoWJgeNt8bQyqAVDXZ5WYfxCQg09ZndKLCOtxRo
HqY6Cib4xfJ+wNNUgHSlymF1mch8RismgLKyidHZGypICjx1+9/R1R/pPUc3XI9A2a/d56gq8W1o
+aqCVejI8TN8oIcW9WJmti29cXO/Jp6msDCEeHhKzgAl++3/sufUaK+ANcSseajKcn2i/67vFdF0
xrC1hJnEy7r8QynRM4boln4ziKR7p4kRxNokLetaeATSB/g6HfEvLptDq+5igXqzydQasxZ15TjK
fGniXKRcxl84NU7w0JHoYcETJffzI2QC5u1JAegs3VjtUZWYQXSnGr0p9w0y6I0eOlY5TvD2N0RB
+9/gwmrceWbTCaOORzkzFEzid72nIZXCokFE1J7OXlZio3uemw8KjOOn/gf+02RQ/Sio09+BL1mm
hwhfoFL5rJGRZuQ+b1l4jaXhACp4ZKZzC7j9Zs1a6x87EP4fwBYGYu4q/urOoPGjz+7jRlMEIXbM
E4HB6ewzhApmzo9L71t+XTpKhKs4IT69Usy45ZfjSykdsnHrZaVWgLSAenbwtCJec0V4DNZTUgrU
UH6B37bBp/b5/lR+yirUpq8gq3rDhXnzsJzhl7ImWf9mFb3HfD3yquHgZI8RzmPDyw0cd5QIgar0
LxiCqf5TSpuXR4wzZTz4/CPyW0f0lgul3LaYwYKgIMt0bOhCyxLfbu3r+Aunghyp6VKQHomIYkH8
Gnp0tphSDaEz22ou5qvzJ/o2Z3Fu3Dar/vmfmhpNQvOTw715WTjUOr0Vvze0Ows57cMJ2GXOi/ni
ztRXgaLo6vRLz/I680pHGNrqQUGwf2faSYJrI+Is7DyhHGqfYKn+1DEl+GOAZ4y/10HKLrQ6GUG3
xrYmTBTw5FTQ7tGoWzyanDM8Hc7O+O0dKCNeWanp9/WHl/cxVdrSIOG0wZ8ohE31coTsWefTG6rx
tqs/XwHSoRjw8M2XPIu0fOBGgl/uKxavvNaTyH7KGpnhbgq2smvOWKP+JEc3gEWGxaUNYaXFL88N
ojsmkgrS8Bnph6VssD5znJZxgItwwHqzjLBQ6HslE2bB0bNoXWX12qAyT/pGvMs6mk6a7WFsUtx9
Jr1lJXX8Cw3cIlfHIjQBctt9PFjU+caJz1uNN2iAc7WwokBb73P7cQGgEE6BZh5ltJtAPUWfChtZ
z9co5c8USRzlKh0649klmKxOykFF762iYuvafKWpKNdWQ/UBDtYl4GtIv7v/xVmUZrcNxV6+DHGH
fUC+75O+MSkkwJD1M6jGGdM18gxqKFR7YaQRVA6cK+kBLc7lXAJcu0CehR55b7tgdxPbpZMGt06F
H/aypsSAFonn2MRbn9kNueQgw3dVo35FtPH1xJbc5JB1Ldig/a4d+yXj6kHliHSLlhtl+I5SyIV6
9NNXHOC3B1CoVbZ2xkgykRA42qX3dSwVdVUotrgDZNb/p3vCsKaQ+h1Gqx0DhflvlRhjIoAa5gea
YfBy8J84xNAfSnVbpAQKE/9k5BPDQrXx65e8InKUj2b3rAS8o0rZ64cq1eVyi7aOI7s5yjTPd9k5
sbsxmJqShf0RSlJcFyr7HL4fz7B3fPXip7mBmGwbDqAXcfZTNBtwZtfOw5Lxlvz207bGBfis74zq
sQnGoONkY6w7IygvENV71UyJxSLQ2Dgm5GE8uhFM11gW+zYbUfe5LauSPQsOcfxahIJySLJ4k2zP
Br87WnizJ8yGbgJlgxn33ikVc9r8lSyRa90rYjExr4BhAlsxtw29vVDXdcKjai0IXJ2D+EF9AWNY
Cq9aKTySrwTkkv+D8cUrdm6wFLoS6Pi61WmeChMY5DEOYO3pCkkBMwEMTDIodlL2W6piTFYtsCIx
j/eI/s7tJeJvPNqkiMXk598Oe8Py3akihVm7Smc7VJM8uCvx6jBKX6YqHrka7rm2bJsmqlsMp502
a0Z1CWyCP8/PAv7ynABEHDeP390gWU3OOvCWsK1pRWVxpBod3VXh4kE2Z/HPpzx5EGJJOIv2rf4D
hJwwuCLQpzl0Csipzkg4Fh+RNBT0UzJJMmKcDEe5rpWAxY/n6Otmu6vTY/JJ3zmtS3oDTXzqrRnj
VtoZZx6ZBauLdpRS+dFHf2YeDyy2AAj+0pPQkviKI0zgdAJxExXYWno/egivgBQm0qCtwMDlICpy
u3iEwnE9/Ad7/1s0NTOeSz0fc6wp+Gq9fb0Y0B4W2bind2BuBNQJHL8cspj32IAfWImUODLftXw0
GhMF+iog3YAdSQrFWT4B2n+0gH3dcVNKDpfEFbLLXMAqSm8ud/sLJZz2+3PJlhAgFvGDZuJ5YzBZ
QfeGzdefAYYIbNUtqqwLxU3pPxt3Db0LOKQfj1nVeX7H1afii+bM7PeERBErXEnJnOHFtX//GT70
TNLcpHJbKXQGxdVXbzon/S7FyHsDxiaXvil2veZiIoTtVir2ib3pzjX2X4/Df9zP9Zcq+brt+aFw
ma8TZkg/e7CQj/rVY8Mj3uolmU81u4LGS3hsluY8/lilXPShypkcb9RUVmAfVc86e/2rwEFCR57X
RB/kwHzy2QTSdAIEz2tBBMCcyGpz2Q7ceCPA/RFE7sfJdxMJYEL9nneggmEFq9tsIRPeQJvhPKcj
2GOrg24KMywZqRMD50z9MPIT8wKA9HCy3FSPNzLTKLVLOKOTIuY9PX0eOEVTgQG6YlSQGtH3wRA9
0xEVtE6Zu0Runao2q0wrArJszXbcePo7ULfG1ksoa32/grSENZfFQZR+NV52V+kj0QAKYlFql/tf
480X26uYC3tXenAjc3JZ+g0kz9GaVDspFqQRhZgHLrH1dJbo2Tq1yZfFIMWaFNOfnJy0Qs1QRkUg
tjcI1xYXAoCgJrhBbTmZ0cPh82JwQ52v060CuHeiV4ngI6vM6WT3nVpdaujw6skYtT5HcrE12mvC
Ft9HEn+dLrIQCEcrP2Qp/7DdwnPrwBgAt4CmvFaR5r4Ucbtw0PN43Wgs7fL6vRgCrwXZscjcdwhl
dMx5tKGS6EWMMrZzRpmkR6u8ku5BriDXcCCpgNOOkm8WBzsPnlGS31LiAwp8qCqZa/YbHVmhf6lR
GaWFjqm8hreRMDQj90p9SS+gtzi65+y9rgdsBvzPlfF4AyFwAsR7QKBDTzGplMoANbLaI4LBQUzf
tISIYvUUDYgEdBmF/GoC7zydyH8y+ye1AB2yTdNFEZbIRP7QnUNwZbeA8ZwWELXReEpDhvj8SHJo
VwHIIQ7id8wKzF6RN8//lf+KUbdKvS5yw+nRY9MGuljm83FytmfD1D2bk85qyeJQrRLwQu7E2qWT
GmStaOWQqT7FOpz0EomUAIRkSvrB64FplyDAjy/hM+gdoX5D7iJv/lvfhwlhusEYYMBcc1B6+x49
mSpUCbDrW/T5IoUVnJMbghhAs8GhuDBzje3VOnXB6r2MWlw/buWzhNBoWA91PSfxMqYtgLpyu6oo
CUYxRUhQTNd1fOLEl1kn1Bn3C1RDRM2y/YgtrOuAnxxAOU+8FIqmUl8hoPGDq34es8qKCeDfnX6k
FW5cjrmAAVXN6AgFwD5Nsfr9mv3vz616r9v5YjdprucG5iFzL/xDD1oa6ZUKslWpdhuaVWXMrA0F
NEAsqhOKfZ+v2BewK8KOOntMKGDfrKkTxvAJ6kyVFmZXPGfjHt0n3xDZAngObBWSktTnIwwpVWsr
K/fIUFz2lOginUmj04XVlKKSFwIi1RngvTNjPqUna6ERPmzZVYCq4luYuBS4VazuenjCEmOIMzqr
PGEjWdqItieAIH9TW+Qez6/93GNIq/wEAgiwWNgRnI1OlnXt4U14XLN+mey/P/+0tWSTJ4G25OZb
BT13DuF07mtyDAaENBiImbv3oPsZ+CQlP08rKZv6Fst6GcimmY+zuTlgzVrX3YPMjnMXjp4FMJS9
c4XI97xeykCXiDSYfC5+O3pyWvocp/M2ZxRxniawH4DLWogL/VYaHlv8bPKS3ftloF6j/rup/JKc
UdY38jRB0ET9IEhq0ItUYP9K1yGm8A7dhRLSOWcb1uv4FD4a1vB4JxdLm3NpXqdL2BByxHDDQt8u
sbrqnHJn3V/U15ETg4ufJzag1S4VStOuS1D2Ey913jqgiTzXejN+KQFgQyn8ftUhYBQmrCJP0zct
Dqh3Ga6UD6HWik2lIKrwmDhepRYOL6GQSbOXrOaq5/lSxbYDmxhK6jxjsiC1h3FB7vHtHizvLdoV
qKI97P8BnFzgnLJaXiBee/Cwp9GI5ymbbZNqzQwrOILqpu9pmyRL/HRcHp3gm3ELnx8knHW9CWwF
PrdaGZer7iVqpgjy/TM+TrCNJfEmzUGRx3zgzPx5rPGjkwghXGuDjPYKrwKlkC2GYIqxpTt03eB9
bV6JS37/nOHhJUmPLB0oCFBmM7ZqXpt1Tc8NS64UAGHcQebSzS6Ympm3pOGksdWpU7katPNanKue
zT6NFSkadigg3TusZ/XYXM0O7B5c2x1aLQHUQps0Kg8vihxbcnXeztnsO8AA8Vr1cxYMmjO/3bWq
gdx+P9CcR5XgbuxL7LScjzFWBcb0Y+8BDLyps43nPCGSR+OtWZ0QR/b05F6W+zsgjBgb8PZLw84J
mOhnSIjyQDuylz0ZAiQFJKqeOv8Yo/HKFbqqBz6gU5aBjwu0CJ9h0nnUiJzDPdAk0yfrDucPhsEI
C7bYBoX6hTvrzAS849pHiHlMP1tbIHjNXUyBFXA82VzYmV0awxN+YZGNxecnY/bqSFkXdBtqcTYi
XRYvepmeEvngMG8inaboWjV0yA7chnWIRjl4xT6mjJOne3tmcEOoq3wQhQPf/945s26xaqOvEkcp
Zemg7cV2oGDYJZZ0Bk4vB8dsUTi8bWgrdDL2arKvQNOd6BddemCPrcbtKB2wby3eC3+3/H+UOI97
W2+B1zMUpVOGOMY1SGq8oNpSD1ckJ/4QZp+/6OEr0nB2/JuOOkm+qhU3OKHrcnEupI3/ux6aVaki
OQ67Iwg4GTAJ0XhRYUbKbnc/qCnx55P54f++5weXc6BwmDI5n7I6lSb9eu6Ta6FXoL61s+me+hPe
d3+DVL+DOcAo5E9MrBzi+P9AQvjzHNb45W5fXmmb64nJyszIvnhcCwmTXE6sguYdKAGDeLGp9bA7
NZQyjVjt4wk6OBK92+RbB01FPDGJSDZQJcr9OXsnH4/w+VgEonCHy0lHKHia5gdWETNfa35Ygmip
cu1Lu26ExgJEqvwvrzEsaxM64s92nP31fu41HgBsInaKeBAcmx95WPe9zFuTNzDfKRHi/bkvyi9F
5UlO8wh8lBJNQqQp51+oWlisY7hMYU9vdWLXJ5KPIPfrnK9zeRaqOoss9UfttBGcPUdom+sKGa9x
rElgsxE1qdiBMasI+ooCriUe0KiCaUVJNVmMSaYc0SXSUuGW1iXiSYjlr4GridLNGGXpS5SXokKI
i8lu6u1Ay87D7jvX83r4lWs06FxP5XEOeXVA7f+cY5SGmmK4G5jh3aBeuHpx3VsnW6qj8100cqHI
1HcCmOZURjHRaylCnOUb1r7VfYxMTOlt5Ryd1ulDrPWQQAenV0Lf0tNMeidJrvW3JivJuqyd+SuA
l+4WEbt5JKirMW5G3vR+z+NIaLaQVM43t7OCm3UiE8pDRPUid4SuQL9TlUsQl2Tx46aUTcE9sznL
VAZn0+P/04gGxvbf/i250+TGMkcCtmH40C4vQ0YEw9oDmUuRp4te5BMsoy9ssV/hlsGtffNdJkdM
lZvFZD87Eqh2MfYXRuh0Ys8mxR1NFM8UoQ6Ae9BYicBnrl3GfVlYQGU0yZek5oh0OIO8Veu7yZNT
yMX1CkCxPffgw0jP8toKIibqTszuxrYbzjwFIgcW5Te5r2PbqPFkCh303T3QBfXw5FAGJikBcKsS
DWPmhEoJDEBNw/Ysd4ItEIBogeNKq4C7LR5t6tw60LnX6KyhPJcxhP6U6Aagw5b5fPkeEX1seUob
GJdx6bDQlBahYYiJZ/GRS6kg1CxhHB+Bw8F6ZqRRZ7aDhB0wWdljHshx67zoXVFNRXs/nZ7GYh29
9RwxOweIfCQxiLw0byTIAPEXtEv/AEgqjQps+UuF0IoHlI01m2ITpXTTX+i4dx2jIq6GPjtRMI5W
DCVGN6yVHJpged5B1YkuIAswi5QYxogf+6yMvw47jWxbIrvoptNi7IhVl/+7EOcQrrM4Lrsd6Yg2
aYYqAHJF8QiT7Y56m2eLQ8ivRUypy+zJtqGEvSXT3FU4ryW+kLVpWJxoxkpkTXSZbrTaT/rrJ/CQ
xt5HLq0QikjLdy3jRQzfqmXQdXOVLfp/528L4M3ahy4zYyLlycqZNgzt25RhEsWRwP5asOsRSio0
Le+1KtPDSThXUvlcKT9zIdaj9mTR0MqTCopUaaUnifS/a/f986SFQ/586SAa7FMVDZIAQ0pRAJBm
ZO8DqZdiyh9cQErJgBmKki9PHUmgRjoeFqGOftTujhkjBnxzb15k4PJ8QyUUcA2oWwzppRoYm3Nz
43YvrOXIlk3dd9SEBqeLG/buEk/fKR9zPzLosnKr2ezmjP/Oco0ZzzSGk4n2rO62S2k1QHbfiPta
9yktQ+54oGCJf7DoRlYHdUefoqw/xCI+YjrLdiOVzWK8kbQQ+J24k2PqBkhb31rrzya0LDqH/NMt
R/YtDtSO6qEHg/W92Rza1fnlFBqy2rdV0tXmapbuXZPYAXF3dLIlZMwpBaOvxfs0f1ZXZAleksTY
5LlwuZnPZznsGA9HuDKU0KWZzHA+cjabuwpu1XRq1SEs5xOiCleL9K95pdsyl+T/dSlFvTQ+0J3K
y4sf3l843cHoam4PJpTO8DHx7nYhf7PttlB9H5hS4cB+AxCQe47u4tEqrUPYklszC03Dh5lgqkI/
kQ+uFqbJqpzEPM+LH/LjTggbtQWtAkbMq4SVy6ccrQ+d0zcwScorRQuE+4WUoPqZl/7/QQdi/XRY
4Df2SP+ncKrMOyppWrh9snviL6H0Oqjmf+fIb/vvwmRqR7TuAiPNzKeVGeYvXauLCcXjltd1GAc9
X5GQp9BxRKz0HgFxyNJxC7NFCsGKc4uazrzb/iv1jt8nszgTHk4GXC3mK8ejPf5VBWYm50VI/xz4
pRGFoHhgWL/4veiVnpba9KvqGo8+GIwfgDG2Nltg0EEJj9etMmHxm5mkVP7lrddL1AzbRpU9Sbsh
0qQU2EMGYkV2L028MM3h99RzDgTyOXETD7hmAbnZaFLRmudQTWKTn1tXE674B/MV864rSnl2qtL1
nt3o30X5QQ35Q64p8NqXVr2OhX40sfOXwTq8ymCdsjNF3+ooxM3rrq4TN3lqp9cqEtH7TOs2Vr9I
EriVEy5sIxB6M+pdhZAUr6O265RkJnOrNnXmMC58pC8PRG2S8WnCNtlB45hqAJAxwrppp/QiiZ/t
23L+dDB/sP9S2iZKF1n8YV9v3ASkdRZGpng1x3I+DonHltwffWjuzZHTwJ0BP5eVS0m/gi+Kr0QT
00ZvYe9E+vbqtXJ8bzFbasGDUPyvHGfgwXyvCARXsX02vhk16rlhRH8hxA47ZcSb2bY6zVffy5GQ
jteZcAub151Ay/60xyE1Bx0bTYO57jPAcPh+HXbhp4vHXf2H9GjXfRAwkfMwJkw8GcgKusNloFH9
68O4uC3RkT6iZX/FL9rizbmO7Qu8YeZm0Fq6FbDS1q3U8PDnQY7omeX85eTXd/VBYO0YjrHP1zwJ
gI3547P5SQbI66EUdvI6uYqtNre+bVXxbXd0vTp3mHjTkXrVS3XrEEZd/xcFvxEy4wxGNTv7S2dh
Hr2GBvTbG//M4e0ldN8PA+KtJQ2v4tqPu0ylgWu0dLFDjwfl4kKbtuUwxg0jKeVuxHJ4nv8Xti2w
Lbu8MCqps8XYN9+8RxUxrusz1cB0l+iLo+1fJehshMnQBR41zTRIPEU7CJYNyVQrAWl0a05Fh63r
RwXG5YyHXQBupi6oFSrAq3VMzCDclwLAYuUDjFuKFdwQW3Mtyx+wa8nQdisxhozA9g/SNobD2Hfp
xgclhuX4dJ1k2Wo5BHVXBQgeWTikS4ZntKigsRgKQA2Ck7XFHu9a1vcDO9Ii6spUx+ar+YtmfZ2k
FJSNDLXir6a2wUegy1yyyYJgW8HEuqnyo9TInRSrxk6hvF+D3vZ+plvVwmR8GpHNCxvaVvEIITT6
1REWfUko8RlwS+GIIgCEHxyMtq7ENGhaqbFqvbN0eKbtwn+AIaytUQ000+ncrk6AWWqc0ERXFrxl
1MvgR3LFsJBn6qmb1bXq/Q9HMN6UIpT2CZ65vnii3Og949XH0YCXYcE27jIUJsOjYRnpee5rvfLs
jO6TGBegb7Efb4oloEzLLnIWUQTtGBiTPkYdbJo7OM+hRRFKB+c0Z6E3brv3Vsc6g6inb5pGbyt+
eBJxyAHrjatCY+WYG2yn89hGPGQIKOS249c1uexbJqbjwWzoBvrTnCIOzMMwZLcIqlbNkYEKMyyH
SUQ5+JulFW+ugKvyoXfkqSnoUyWthH4cMtqduJ88wmyMtLzEpAzXkYESkfdXmoJmXwghSvP/ypMM
S+iBD8A5Rt7vCQNrsHC9+68tKGEp4yn6pWc8/JFY5099s4wQOq4pxNitOWO2CWaVWzX3OA8yKx9q
KEJ0XBeUI/YFb8VYRdsuT+pq+QDtr/uax9LtMCTYnwn/bltuNFyIFz2JjQ3M59YUgAPl61wVCTKz
Q8z3tjmoKXyaPfuLSBQC3eC/i5yvu261/KSEtPaeJATVdrARmuNbEV73nA2EIKAJF3Wz8Hdt3BMf
ymjhY9G1j1kY9x3NcboLKpPatLzEzUuBHfHC5AY6AxJZGXBGM+SaEWmcgeG2qZK+5cm4WDoKatE2
+wQGKKqKpwZD5RRqRu6syWL8sRGjM5WVX27MuCYJs1e3kR6PuGLhjHvz8Ceia7chTOvH/4qsqMKU
OBfTic1H2KjyDYlhBnIUoWleIBPJlORYFZUu6luZiCvUsOgXWCrmuJp7P3Vpb+ulwmIjGfkQlyWx
bmCW3QxXVIIC8dfJ7aa1DK/MtIl+kOZ299rcdX+DB18NrLdC7Fbwz+dBbftPSlwdIR8SGXAGGN0F
NcN5JnYYXzAA1/+19mTgW5IYaWld5Sdt72JgV4GuhyZPXYDBKsxB4c2PPMWiEAVEhbGV+23hSOTp
/YlmaMUOl0l/yruGXyEm0UVPAV0r+KGVh17dP61dEBorPKHXJXmv6ILNySKiawnvtY2W2w24sNx1
rPOLq6ZOdAOn2z16bXjzU2eHZmWYetTBya0XyINAw89l/J9t1WuLLkiiqOfKQAIVzX7syseAP6OZ
dMRcEND1NvflcxKIMYRDv/H0Y1CrV5JPlkobD5hVKSFgK3Oh351q+qxCIdXny5ATu4K7nbwJlPX6
D9kcq/gLjTr+d6VBAvy998WN4iyO48mpz01mYrZGtM73qQT63VNW2ViKwN05Tea84r2/yZVN8BBq
GGAAzUOaMhk8lOSd6qx+D4O8xk4dXUMJnnZpclYnDLDfe/2aLBrAl/8juxCbsWlFSlZZik8+VXGT
yHV0d8GrXKcxwKGWmS+HKHPoxvpDGGS8W6tl+6cso3vaHdDoPkh6Lf6TzZ1180NPOs6YF4QsMmy/
Zj1hUA3e2j8y0UkujiTIrHXIHxjUKoDsijEICmV+awLlg/z5Qo+mZBUCPRnOBwlViGRKu/4wGHyt
nbG3XxK6mO5UMYe579mvRuKva9qh96GAeUJE8C6ANq5ruibzTrXBiXGF3O9VcxcFswNsvqMJNS5u
ERpbdJWg+KQauB08yiU/jxWD2jcz3RAHzRDNbPpkAHURzX9ljnPHFWmJieDM7mLI6N2MPAVgu0mb
nmDS0e6YWjxnqwo8WUDCpY7SYbImtr0zSdMgFufFi6QC/WdkLt0CCkRryVRk5WL6AKT5nTWRDjW2
NhcvBenq+GgSlbEHiJwX+e8pBcPJIO/FV6xBVF+qSCnMgyCawEvYEW3D492PLu44gA4aWh0xcmd5
mORXYKmNgBzrMptaWpD/PLQ8eOQ23oq5/ncac9bJaOUqN6g+TdsXwyr5dDN51d0mJNsOj6auvVLz
+dJR9X+hGYg2bWdpthLXUZ+yDe0TX7m6nQpwNl+9EBGnZeFgZiuOCpb2
`protect end_protected
