`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S+NPt87NQpxvGaf7XnzMdP/fozLeYxnmGHUKXjdEjEGgTytddUHon/69Ruf3u2MpijL8bYh3YMYT
BA51J62O2g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eWhq3M+oG4VhbsxAoFhy2N5ckPuOqfzYjFoOdIvnmFjZB0XUaUK9OjRWeAWJ+64PFaQYopky0Fq5
SkBYJ6qTTu19vcRrPzkFhidefwIdFd3RbpMr2hTYt72GeQEFiOqvjNTqKCDsYNOsePTj71Ipj5wd
dL4PQcpPvGjWJDGFpag=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BKY5exne6X+eJLRV3fLUX3qUSafuGMa0WOMANSIXiCFfs+cajksxAlVfV88tCmYYHaWrhJlEPvQR
xkT8LQoAnw+tZL4Ln8RKebWTRuAOjySqiXbo8wKwJn3Xv39necQ8/vETp7moOCtgUe3/HeVPPce4
baRQNPLxEaKezVhSVCk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a0XmVcGfv5DYijcftaZb1VKT3qaG0lBBjuA11+j48/VERbpZ0nci3Ixv6vTTp2coLRgRkdIm88X7
sH+2l+X74rn0QMI/s1D33046hbEIOJxTLbL/oRGFYB9Xatbwev8bjLFHBgV0G3dZlZKOwckD83JE
wSFvi/Z0yJ195Mm8+UWSAsv33yOqFHNkAdlkHj7wtoZe6hAGcT4huN7BgmT60GSLVo24qBZKcJSe
W4d2AVEllk5wTRpWTaC7c9QgQ1W+dk3140cdFRGBUXtynaV2aRH91pHkcVG9sQ3XqjBKvDbu4v6q
FeyykQLxCbA7TH/GFMdp5XhjCoj9KE6GpRplQw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I77KOiMugv8wDv3Qpz9ol3oVg4VmT2J8j1hDucKPSch2XyHXgKzaFSUzI0stUpCF6mhMBJJKaB7C
0VJyPqkc+IZ10Uy+CwjZ3gik2aCJtFHgbPZEhP0+XKjQBLwHhckgiAsQKEFBg64vuzWzJTKcrd8M
y1dHROrhJIJ2ZETFcQq82/pJKlRJfZtZ/6hf4Pm8j1HXf8PipItmRfk8oT6gINQTxdgPn+GPPHQA
vOqMJgeeNWmb798ytYKPyWjNHH8AO5w9pVD8MtvX00hVtMN1XB0GzxE3WTEp05lkA2cus+O/sK1U
qXLYWyaUDH2MrudJxWFhrfcMZOEzmYNkFxlVsQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dp3qi42ziRXBSD7E3fpHh0ylwL65MH8Anyn1ckdFcJOcolKl5/mO6xYc65Lj8dDpKGL8C+hgatRF
3UCoiWfsnfEn7zVRIzWcy/HoIWT7NAa6mf38jRFNz6x8/lkJVjX7fShumTdbhOLLUB0egoIZ5xoz
V2CyjRk0r+OjiBqnq1+6G/4SPn62GZ20BQbmcf1ZCHSQYF0FenJHIvqOYzEfkkm+R/zQj5ZOgPVL
5lRFhgk7DGi4HUUIOebvz8WvCEyuJfEPx2GnES+CuAgPWhZjz4AuriOd8BhXLQvgSsv8yDsUnpsK
h97SJlEQzELELZWb+djosAWEpy2DHJ8EvJoatA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
W586lrbjJwPkA/cUT6LkPYkoU37uTL5l0rnTISyfmy8YP2CQ+irdPfNKZUnJgeNz4zvUerii2KTV
HfEo1/Xxvb5QjFyH4Bb+dVNCNtSfdQhJnfKHFN+fuRUrNm4VxmPCWY2ZbZ9as0Jsucu/PUk1a8tK
3usZF69e5bErqilTlhYG9aZ/2KAfpE3W1oU99vwageVTAphGgFLSnf/Xdpy/OHY0IxF/EUdRBKZP
9t32eYnwZxy+UrpgccF1rEq1Qa74SHqgA9JcmjE1n+EH4UOjP8NRB+8Vqj7TpZvI0uJ7YM8VZ3Cg
rJVpJtAFFNBXIWGcLPYzmUJuk6boDFjp1kkodJNKSGqbq1m0RQXECL6UtzG8a9Bi9QTMoe9oOqGV
3q0oNCIdl3xKxjrf26s53XW5H6NP7vUE/g5zQn07oao2/25W7l84Lyy9m4r6qTGo2mm1vjSrelaS
pTUSN/3pIEp7lJPnmq3Hp+183xgafhA6QqWIn0i/hQXNxcd02vpA2Z96sm9N4RupukX+JXVSD9Pr
p83SKWwixHFermRj6wtaqJlFzU6NL7cQ8EX4JPup12oTWx4Q15dNOejYToUyOL/4D/ziuphZyNRX
yZva1ucmO1JXkvr0kcJBw8PeT8X5dCvOZDJfOc336GS9ZJ/wOCBrmGSvx0u8G2IKVtOfltbf+PgN
gJ6OCeIZv9jQGb/pMKgTT+IRO0PYdAxR2SK0+J/DapQ6tH//fC9sfOMG4BU1EaKzQ3TTZ0Vin3FE
9gxpzl3LmOb/CIUMZ5nD9DQJoyOh1ykWJ/rBvkiv4nMF8Zq22sKP1IE0UYIT408s5gTv5VyyU03s
K9wCOuTLN0uaVL3hL5EHXJHhWuKeN0l8C1C/4mK5+6Ad+ROklYdtLCqLehl18NNFs/STE1ApK4+t
F/4w4siBHxmn63EO3cQdPXbRQSW7uSWeNErc9bjZAgQeOw4v6k3wiPuegUwaVMnmFxKX1j6aU+/A
oPrOiANZM2xyo4Fy9MtEM4vkUk6/RZVdtHQ04euHnGm/tTZQ0FyFZr35vweaxUwoCNkWWxV4XHKW
fzBZdL1ehcRuvEmhunf56CkfzK2IVTbS4AqYkOpLDqs6JVjE4mUwde9iQL/8OeGfRQvBoTVQYB6y
iJHu9SSsIHp9Q1IXboyKRrYrvU7aIa2QysEpL25yZliDWRllungWlvouxIMthW7M7BgiK89xRcHA
KaMnCT49D9PHhgOtkSO6xro1rxfKZebDa+U7TpCGHEy2E2uNeDiLmZ7m8Vh9SxlPGhFPFa+IAIgU
VHs/Bt1YT8tH1JuFJ1Ocjk5ehfj5imZtAns1Lorooy8GmW6ezrv0GKwPX54uHKsp2RPA8YaWhUNN
4LRDmfsiI/KnGhjsCiKIpmxfePRPsJNZaIvLdgfwkHp6ezkoWXjR33oWncM6vn76UxHN/MfQaGqd
tPNP7umFuFEe9EvKNanXPZfQD3wvfemUZgV30IFx7oz8S1SHPkNisSV11FlL/MFlaSW+slklJEVq
4iZOr8Vfrf9IJtSBkmnMNTEyk4WA7qNKS6x3wsRmhEt1dKctyfLTX5Llj2yAmlYykbBGwmHWfMv+
US7Yv7rG1taU+C1m8VjcxPDi5CB5tvXL7t3uZHYAEamdqbIRKELeTScvw1Lt0iirfikTffgp/d6k
wgIM34n/YQ0J8sPCOCXdwqE6qsKliMwrNdKvzZTDgpaS5ET70DuHAlV1s8O0kcX6aEXetAmqxHmY
h/SDcr3PiPFk4rwcpo1H9fTGfDqiDY8rNrydZSm6IIQVLS/JQ1TfL/+KBh9wx/gcvyiJkmnXgS1C
G50iacn8ZIeBgCkEn+BLl5HDiSsHG0ggRE6eIateA8Vz1OoBljer3/H9IQGD8WM8+NjFUKE4/Umn
sJIpFXMoo78ADcFOitcV/k7ExoVFetnkqpsFXHEfxncoaIwufMWytEucYsWQstVA2p+wYe5P4Vza
3LIhVfJaF2LsiDFmQuTXVr+RWkNQjkQqgpM2a5Ig1Sgx+O2SpkEZURgQxf6IsQMHrkOJgNl7hdSu
T02fNSZV7csO/V04T8a5wSFw30ij1d6hPTOHGAL783PsgWbVc1X+5mU8JqlH2RlBocHd2KPnU0kj
RBH5yNFbT896W3qGFFIp6S290lVWdhXGV0S9kWBC9bfdUsxqBfOh0otAKd7CyIl2k/o6Ju2O7BoL
rul1vhq4WvNMjxB9IKeiC8/CJ233m3buZYAsD3QiLbj6xGdLIlf0xsFuqhpv5Pq2RzK7nyAsEhgR
Yqisy5p5Jx0Z6Z6/ONbzJB1zIVdYITBvAJrx9aGOmdu4Jw4mWlegxQqFaxgotfgEiQOP5ehspBJ6
KBbCXy3i6utS59lj3uuce1GWCKJGijkUUxhX3IbUPN+Vd8arBNnAJsS7i4YaHmawCGD2PWBLgGSG
Ja6+fy9TWENkQuFTwkbNdnY+7Avd6YJ/myg67eK2h+w0ABn8s53rSbW5UWUb0Lv0W/Ui2BephCXA
w44xPL/MxwVOT66KA4OyCz8taUt0qr9HsmSKL/16GngywYDLuYx2Zh06eDkUuC+hO3b7/Y9Mzz1Z
kv7J2D3uf/jPd0qIYqA2heEbsT0nFelBYi+6GxZTKoTK7iEi2sjRolwfXW8O0Wt8XaVGZnUFloR8
km+A69GYK7sgkOH4jmk73unOMKV9x0QJbwZyiwcKgPtXl9tUcqIjemrj6Gg4WRx7fSSxtFGSBvfk
9trnm+n+MQO7GM5gEWqucW5Qv9snp9peYINNcZW9AoayZVST1niagqobbv3178eYZ+HsTFFOBmaU
UMdZhShqX9mVO6tJv1OLuqtnwENZ5ia3ydrOV7fz+DoUFTIXYfrq5VusR4CD+VJ++3y4e7uAEiaA
h9S9ejKSAif2AnwR+sMlOkWLfbbXroxGDHfMe17OAkB7WYOrv9iqxt29/JVh8cdfKLZMKIx8Fr2r
+CKciGu1eZytb2nSTp9pSrKOjEVR9EzG3kdEfZNHwL0zdRWz4YLz2NfjO1rrP0sm164Gpt9kV5dl
Qx0VVFooC8+rYHntISrrT5AHdpnWBCN2GhqruooW5DWdjaX87EaDlbHfXmWpL6lmr47offDFqng3
hgauISq9DOUoIqU86rgj0B6J7nE/fuTTcD6kzkFK67gC8847Dka57FpOkNfHDRMVH1ketf/9mHvR
aBV7Bc8eWDE9jGZ0tInHSqLr/MrFEAyKsaHsk9qSO9FOodxl2kBw4q4r3skuMD56Z1g9r+hBRFac
MXXI/K0oV66EFwQjpq96pB42jlKA7yl6EI72jORJbbpz3Iw16PQnFDvRH4WTdtmOJwWYXrmBgwzs
4DkfD/3oIL37oqMJNtbF18ilCdpDOCwBaCSa5Bp++aVN/i8Uben+zkJf4TJRojvLZgW7PRlWNun0
NGERaq/8D1C47M9MdAmwEPZcsgLvOftLZZ8+ruCSq1ijLj0LeqKEq+cufNd+88lmKWDN/OK2VmZk
aMGyzFoEsIiJSp6T5h2CYEGtd1cWR80qi50YSifVHpiWD4YC/s1mEnLz6MzOUgMHGkjd1K1U37JO
fAqXLK0l0EGZmZ3Xx8h/DJpZbVXyk2CdaKOjP8vye8gZ+Q5jJfx/fFgw63PJEqZuCCf1HqYqCgB8
2lJM5/llQ9yZvaxjgmviRHtG+9IVoe2XVY/6mJUv3dcXdDUCgdwAuq1r1DnOX/Rj0v0lzSbZcX/1
XYSSocn6jt2owvyDJnnM/rfR/j1Gg9m7OCYDkvk9XuYwWa2yWAmkhr1LRxHmrkrZj3aFk8hRhEG3
3X0Otmt1bQ4DVpJoM9mkE+lsVDYLgqLE9Vv9YTjdmqSwsI06UNV5iMCsjKY7k+ltfnJen1rMCZjY
sCqyNuLxKCN+svAWW6ZUDVhX/kY59XJcJJiikdQqQk6w9gNmOXbCwpHEL/8nvjvjD34gc7EpfBmo
S6O46THooWJ9MP6hzzLW0YVwVc16N/iTz/xlnc0KLWD0nuLK2zB+fkHU4q1eNw0NuK5D/tyn1MjR
szyerwh5q0z4dE7BP3sR8sQzzJPFdO+XQ/V3lbNZIfzV1lzH0p+nFyssqex/0qwa8t9E7dAf2G7b
LKN+O/LAIyON0ZufYtr1LrXgGC/tBx7ReU+nURoRKoTALuQsIMTHMcUq0aGy0IWhvX4MRb5+jog9
yttSYwQciqt/d85CA/J99gWdlFMxiSjGnideeI2unK/36BX6c+rd5QljmyKdKm7mW6Mn5uoibf9G
zhn2LRgkdFsFHuxgVBOjJnrdg0b5vHzfwsp4y2LhGIDdBpXrNTXGWssmKtObapjAhWCrZ3hldqtx
ghmCv4M5LlklNPUU0PaFgyPTGKiH9m8bEfHuMiDX5zPmugeqgraQh3Go5SxRZ7iIYL41kCU7vTwx
p5PwoRQu1AcAN7EjooA4b9mb+IZt4IamkFC6scWDthshLOIXfe2mNJFH0zZvog8ybg5QBV3TRwd2
F6+4AEiNte7D/rIM09ia7QgWpg6iJHMVI/VG2I0HSKZ1RKZkzw4ERxyMNuiKrPFBGQTzWNUciO7T
KmV36OP/ih6LstPix7vi+qxm69DP71Skrse4OpS0oRpRQtf+DyjZI2LQySHpzZBwAEMRsEgmcF0Z
Eetvn6wPFP5roOXrXi8OxUkWc+IZTcMfK4jbw24ck2jCd0Ua4NSTMsv6r/LPMIJw8d1c5wN4tHnF
uojDD6hLjbkasfnSCjOJ62moN5B+EBXLjsbqvl9Y27htcb39+JVtnP2JLmzBMwc63IXPNeojE48l
P2xD75Jqg1eUb0jMy6icIcew/1kujWMf2gaMeBB2tLJuw8H6lazScvVJDJTinJbKG68ruxrRoNdH
U5f1bINSbG7bt+QOCb/CYGC6YW30cDVzBjym1E10GfD7PEKMo40H4zMTC0DfTgahOsNrZXEqlAQh
3nq3XB+BAt5X19W9Jq4YcUcQQvuztIueZugOcOPEKbrVwkNUk/INJg0IkOOCXfYkRW+xcUdvqoA/
+ot5aYc/Gk3nBTmwGC81BdblUoetZU8PsqyPaJUlnyykCezUx4vRg1f4TJ16EG2cXzEW56idYpWh
4mk8RcwV2ld7qwxVj7BgDGuXcen0n3VjsAGu9jaml5c6zcJQO7mOM8vXZkrUsvIpRvcFbUCWGqPw
rv/qnRS6siBdP8wEuuqIBjFTZwQ8s9lZEyLlwd1qnWjgcWpGuJ7DA53jOX0m5RpaxQWwgPPsPgWy
aQsI+hmvusCPfcIj3pdp4aD1YmT+4YYM+gQPf+jdtbAYYoYFWvh3GToxsbvvfI8qG7u5j3TiXKmH
Yj3PBhIo9o4+0YxQhIgUYSAixcNqNyy/vUgZMIbK3AHIkmdxwWtk+ISWtpXQKayOXFE1TzbMQN6H
/v8AQ6Q1YFX2T9LQQPT6s3GTgJQucUpD7xLoRDhxD/17Lpu68/HnrxIbKIXRvz9vVjQBj+efBBOc
C8h2taOYSLpiVuNUIsMAf7y3h1cTIaKhT9/cZ+wWA2mVLz4p+2aObWo4Nn0QfaY1My1iLcXo7+EG
NEA+AO06zY6D0BkOXVLiIsekpHzd3oQomprIOwcPr3h72fxfgtMtVWA7KtVO19cbxN7CkXuK3xs3
4HonMntX8fmOn6QsymS7YipgUoKuMRMtHzghUWDdO+FWzi3QmwazaLBL8RUgibxsq/YaP0RgCyB/
e4PyQFz8uJVhWsjKoBGUwWjNfnf7EMhNvW3jogcWaIz7qOKUUBDdpCQ1n0UwQrtyBa+KamXm3tfr
o7nJ6+D5swnPtyW2oY75LhUHyYlP4rtcsM8ZDurty3AnhBCju3QbCQpKvKE9IHF0ha1YWXsmmaOk
b4elff+trfUKTCWKlTgGJVBbfHPH8VNXH/XhFWri+CEcjjDRyqdhh9z5e+LAimuXj8Md49JL0eRM
mTkr9igwtPijAzMOtbrC7g/ZRckpOiU04WGgIsIo8eEsJRtBCuYAN5DKBLqI3+dl5Ay6a+HOAhda
pRypSNpsirP9kQAtvtUoLjOXhMi/dZ8H9VQGWfxEha2QH3o2SKXh8dmH57w7AAvpdS4v9WYa850u
soH9wyxLHfK+sx7l/phFfzhrk3HfXXpBQq6fxG8ZuTj5PtfEbiLpXwe+hZxvPfqmhwepuRqSS6q7
Y65JpXqleujYlCJwPf87OILVDD7gqD4DNVYLCsc66QT68SXl/OXxFFJgbZp+ifQrgUH6seTfGp7F
aW+4B39l6xnEr7JdKX7COvjiKzm39Vkj0rtdxLd0j6EerWepV5Aq2vmTpReUjfLpyeLW3dbbi/Qa
ggLpB5R4ZRyAn6g1geJ0tEaEcZnsI2b+uQmOANEqk1UPPxrO5/ghflquW/wlUgwv5GZtL93E5PIj
UnTbmA+341wC4YgAcruLNJS2jJVTQKZP8U7Pi9zJEjw7x0wM9A1Qbz9EZY3x3YEDsPWXRQ+91lp0
vS/Fx5zlNykUmttCHwReNiZDBOX685/FAc8XZ0NTUz9WRBILhsXw0q/b3VACFRuXljP0eYOfUZO4
7MrRD2E4JFuESwxn1bPIozTVDBugFKsnev6k5k3NOtuKxwfR5Zphh1KO1UCmE1xpFwqgB7ZQbQw+
wqF1GXINLdHJ7bx0kN0sR2q7obIVNorY5IufhTDkzvyEbFNJlBMSfSCgqqxbTyvUY80lzNjQnsBP
JQ9wHFXr6lsCrEqCNU1BEczVmzzMxk5WIYmg3I1Ms7xmMNxPRRyEKN8uf0hlTEdTneX+jbjr4Ut2
+nuXwhMnJgoPX0KWuIyIXC0xWxfP1FVmXIBmtx+JQ78+SCHdlqIPCb9ttLJyGGxsQoYEom+JMHVw
+61pRiAONNC7VKqDIoJTurRctTt8rrfvwX2QZnlJ+bzeCsM6MKC+3xqFISUBZxXtbbUVH9lf8sfb
agys7SYVt0JchSV9sJOfXoxmFmpoh9Yx0iN8qvJqmF7ZFpmSlh7ptjF79pIYjvrfrE/OJJyZdhRn
CjpSC5HTp7gESuMZG2V4cDl8ae3JagtCyk7b2/vVa2i8sHn0rbJ++CquXeNukZOyKjvQ+Ez0FYCX
sTeog9fIbywtr518FmxlA8lZrAQN/obdYevuNv8BWXg5FlIURRGrfKtv20QlBKmsjQeycHx3U+kq
tB0mu/uBnrnnasewiruVAJZSyl4QAJUn6iQDEmv/MQKqnN8Nb+j5OPmNeQI57ztVJ1Sxlvn/GTSi
45msKAK/1SlfvYHqQVM+QDB+R0glUGt8XRb8znlpXpzKf0p2LXBjpYqxBFKbix7Qkv1pvLiNZ7yt
3WOhkxwMnNMeGBwyiODRjqcWgzL1U4IRuuiMrdTfxm2sjJ5GlhKe44C8Glcv9T2oF+Kz72G8JeHm
K0PHwg/2GMBHTLZMM3SDFwgz3+7V0VBSeUuz1ORkOx9iKiF9/yL+uBy7++qZdzbfhzJD/eW4uzdp
TwtxFS63AINLv3r6Z5cCgcz5SLl5UDPWR25Gzot1b64nVjJ8suGJfEZvOubV5LORvo9QB/JOT3fX
Apc05QjypNheQBTg1POqUkv9q3NNXYZ6CPIXiN2gjbL40dT7Ik/yvJvKm3PULiP6dH5vBS2JYAyF
ukcBGVKLscKaiiHmMITSjlV5pvCh9IeKmgo84Jd2SC6hbcjVQsk4LA2cSi8h6HvaocGW9faZvstH
GWsR1yPlj7clPUUZHUNSx92CXFk5ef0JXAqucPUCZiCT6UzSDFyF9WUrC7zRIQ2T3IHmtE13ReUY
aq/sYS32px8IVh4iRddNoTM29iZBywC/6vaqF8vTke0G9uKwzga7AyRWnbl7ule5wLS+WXQrgztl
gt83u+xlUS9LWuYMDcTp0rZChuIc57EwuvfoFohpZZubt84FtgpeebhNt4fuMUP4TCDpWc9NjCGM
3yNN1kwMTiKypWMbHAxtLgS6ILViwP6rsUJj/Kj0zqhf6bIdmELG6hpYEIiFKbPE/bOlWmjExQOf
FsBYlXKk1N0uILFAuV+GUB7X81YSW1F+UVEkTOtp+QdIEBjodRh62wgtL0kDJBVkuZv3a5UFmebt
S0Sa0h0mDJ0kGt9zzJwD5QW5yWTi+BkxM64RjpmZRC7G2HlAUT3huf3quAcx1Up74dNnNM+pg6Z+
4SUbYQU6jbQK1uwnxCBkN4MbV4irplS4hn3TVtDQkeBP5dyuvEJVd60v5dBLS6T2iHFdRA6acWOM
Tub6LL8zmvbxltH3Zph9lGtdiIRfclEcctt2iP4fQJERqJlnk4o3ZdwxSkzlwKOhxUpYNn0eBaN5
SuzB/TkfD0e7NSwRlfDTFni808QDgRBkM87PmS+FImUHf3q+fi3WXyBnTYp+lYw3ZXCeB2UtEIzs
nuSL1BjlxpqGuSZ9dN8zOlMSNPCJH7W/Xd8sjqCfFhVCZs9fPPYmTKp/bWSQDPtCRVFyXKIvZMsx
odzZFkQcaOF4Gt+yU8w7VdnKXh2E2baN18U2PQrMocold+oUZa6imlr502f2XGeuWQmCWASnhTyj
qahUv+CTUhoDQDgk6b+ZFGPNw7HoIP3ioJsrxaU0DkeHOrcDCZ6C4m2klni1lvCWFF3qQGKOF6nu
CJTzfKcUg256JQWl9NdK/NXAfY1Qtajw9pAEL/4UPmfqZXelzn7Mgp2HYBXoht6B9oJmdCPy59XM
QFDeRxeiGgm59Pd6bEmrFn8o4wEsb6uZDz8r4SmZoqaC+W2vMJwqSdUruJV9asQ1qpTU9YGeAX3a
rz7GW2W6iZul87tKnNYwee+wM8sh55uF7zmXMnF5Z4IDZbpTY0efm+TtkXwCLw55LMy8pElP1udV
q1tDvND2kaH9JUNLIlk8XZoSvZLFktzgceFkkRxlQTV4LhzoifMpF67hQ5QEr98mhHDVpN/rOwwk
49WfU6rVrnlFOSgaZPRcie+e+P6DsFjGl2rPJBqpWVzMOilhmgqlOwVVu5DHs/1dAws6JOok9bvw
layrMGButLqy4H6sTm08dJ7wYdY2vxTGyVEjUskCNPysbI3+vhLONytodsI4e7stNaSf3hvAaGSn
etLFvcifoot1W97n3g5yFOSaqu2Q1OdCRTm9AYixcXjhsI6+0P0KXa1VNR6/aI0Ig7aRaflnLEkS
sSa1VUYgz2n3sPlxk706XFGSbW8sNjIM8IK4fx0NR43L0hURjm1jpVkOg2QorjiOGD9DMNycnIc2
oB4/+qVQmjGPzhrhXq0Nrl/soAadErlKJSr+P6JYNF1232NkVYLEZv/C89DCqvV99/425h6Pwe4M
qmcxzLxPp99xLNOM62cJPSR4tcJUqDGgEoia2nUJDj7sSq3+tHK9kQkZKzqa/AiANbyTFJrB8g+X
xqfWCQ6eG/BDZf5dvaWUWDURPnEIrZcNJmHZjQzptfUvfmQ+/SWH62JPrTMmYEIc4643M0lmcu82
CbLeS1LL9vxQ/earcZKPJhQzUWbZ3FQwl8avWNpkD1PcSJBMQuXrGiMaZt44S5wXaM3lLRDrxGEi
OBkE5xHkPjvPAK4c5aI6tWT1tnGqtKkfBeruus6Yeot8J5WOglsnViFsKZvLHfwP7DstCCp6I+1p
CoMG96doEXod1e3AJu3mFCIghVlOMRCc/qNZq5dWU4/6BbkxvVM3LA5dUb/VhKOKAflkCd0jBoXT
zxneVzY3IJlF8dEGOBsXluPLeTePgb+NPbo9xhIBCGQH42HHmFcyvU7IDBsVmKIw4up5l2iGeToO
8cuFnxxckDWbqMYYS4gWHGpc+uC7EkeBKhJQ26EfWxxOw9WOunFEbHmdTAOoGs+WM4S9aOX7B4wP
Ls+iH/MLZBmmRwJ5rOJPaGdiEKpneUsqUTL7lBp09YJaEsEf3c4wi1BTALk4/WzJuEMRwEx+zApr
O98KZixLVWxvgIFdtUsZL29gKx1SR0QivH4Ud7CCKX77h12o9UdV0LJWYcryUxGpvYYme98omKqf
hdfns1OaEq+QJSfXSgdDU4lYDcemcDSAwHPM7pzwEf5RRqGbGRV5DQYB8/7scfeUlOCVogbms3ae
9KRL0gLgOmNaBdK2QIO/Kzwe5/PyMCQNW0h50RCiaD6umhDcyyvecxhYKDtwi2Xhr5Q1nJAtWYLn
YQ4fjA6NeDcneqoN2a3MOPMvJMq1R0LCK1l6u6yum5zqUm/6JD0RNXrHe9aIe+KUt74vf3grxV5i
DKDB0G7wsuThUTnjYyS1dQ0rRsLkQx+22QNebjrWD5vkieJTHUYoXJ6oq83I7aE1mfC1yrlmM19I
dW9B0HL2Kh1j5r5O6GSiPsmhMhkhnjHb18kdelbVuGnBwVWJBt47hMjiiyTSAATpvoXn8X15yQkH
0fkJKhfuJHaPdiFBnkE9uzpi8JQ4oeukAEYSbhF2zn9rA+q7XJXiEdZS83T7h7ahz1QS3eOYmACQ
21v+IS7ZwYBU3EfdkfnTmc0/8N9/NHhTc3m5+l8u5L3YcVGpEf3e6W5KLzHz5s3HHA61+Ge1c1Fs
saKW8J6DvINg/oQbNDEO9xuKjRwl3qHaDXRlUO79yAUkRRhGWnMRRDYlXweB53yE+VgZjxDpfNVK
RZsUA2E49d+Ggb6apPiuypXcJyAsLcEDIkmvKCTTj7pWGvmRE9+zFvbwD/B+ZYhC7xBnHTaaisKd
DRygI9oD8NFR2rtcy/xay3hs03mj4d+Fo9lnWUBRcN8LhjGXEI7Xr8TTC1sKetyL+rTJAXjBwIqn
Dd3Ks6IB0LOaZm5EFxUip1gSo/XZIKvYEnPtVUZ3ukx/dYhakYpSKXCNqiEoSxj5mghcqoitghSd
AqHII/MboZTdC9i3EoakcFdASxoIJzwJ94bYJyGj5nDl5M6/ggrbfLp1XcGZ6azUtqJoRkuHAMfQ
Tt5I90/QYBswgFbdmX7o1nDHfiUqrjQ0PilK+4mj6xIl91HHpUMYrDVfbAozBr+8i9Z9Tww7dNOD
+3W1SvU/nbnIztBp4wr2Rf/BJkuOmZTlC2ISAgM8fGAu0z2L/5506ivkpLQt3cTX3WOui1S9+lAy
oRV0A9yp/0JMwD1Z7Fndgm7rfU2xsVdHKh2VntI2RzS15iDGld0zb2hGK0zsCYbRSbWThqFSTUAp
zFTnOU6gKO0DTqKfINYalKv+d2JqTP+tIsDjgZUgk2zEDHEMJrLmYXaINuUCEL12NkaE4Oh7rDze
Ik3dvvqspciEgilmHWntmVmJ8o53NtEYFzXA+l8HqwpPX9ecyuJRZuc4nHmGdvnnvzH7tOiBLOM/
/sNj88QGz/scWYGvRW0E3ZzcsTQz3qOWCudmd020+W04SxLkKvJxBdOGg5tj+vooT147JklEfMsF
+Il39Lbx286+QNftSd0HA96O9yp5CsjTfyodUres8cQW3w4yX+NG4Ze3TWSCHlYveFxzdysjyOR0
KUZdUeMFR/pE6oFQ3C5COztb84/mX/jHK6a/igk487Mx6zyBFHaiFtifdfkYMtGtG3tQEtgGbCMx
WsEP5k6JJPgS/ARSBRTsbpxaZ5zkW10dEe/CkNO165TyIvoVzhGuS0HT2aVU1Cbl6wDD9/gGPgHs
QGoljmEzjh2vyJwtLrzhREVugRvCTA32MPDjXaYoKRB77GjE2mFeZhd6J7tKjWgl14lZjQ9LNMPA
JDyQsnRamnK6LPHsJ5DqjYX51VTpUeo7T1gEGhOT6Hjl7VDj8zO4CwCojRITxXa4FxKpcDuglQqX
WwCO1s6AG6bVqyyQdgl1Hc2CmhXbxJGmTfYZLwBwNaOqeojiyQ/yQ87irlLJVeRn/mVDkTFtyYAp
xtRZ3l+ttXW9G2M7ZD0RDvcB/yce3MsxalFouq9Ox51V1+mKKdMACYOZPZ+8FW2UVTkyZrRnADbw
FyZF9nP5XKV/GLavbBTmRBhKvzGFqHX5CYr38VH2Kk3wCLOdEg9LEmRA9gFRBNYYw5MeFliDfHlj
uV5yGC5xisjPmqW8sSDiSwKnRS4abh2p2463vMJe13eoF/r6dBxL8UBAXy4voiVdls0BxjGrtqAw
i25bqFhhLcZyxNBnGw4V6/1SQcHuhvlkzYrGYb36WjzZdIeoavDHllSRYI4Q6pg0rz0irmRzN0Z0
ZvCY1e+sehfSWOMmmG65FVoh49E//8T9XpuqRdxda04vuPSEXqMznSFaAjFQit+gRNFPM+OP0Ui3
5QxE0OJp9BXKMw7ql+X/1wpkfK6cPkDssBelzltVSkn7xVBazRm3bCnPE6bz21fVE5BBzkrfLsHq
14JBKrowkjeeifp0mqByL0KG+b3AL2TsE0ox40fXFnLUM/PN9R78MguMSJ3m0mUl9pBq3aroKy+Z
06tvDgmDNQRH4heDGhm4N3Z8OZlzplvCFYTMgycg1AbrpN2l4rFjm7LEdCWDERa+PLobhKZJ3xSl
gvxrb2cBEvwPAg3MPizbpRJwHKnQZL7h1nusvHpyn2QASnhpVcBr3gwIKd02pATnKeBALEkjiSUy
haxcb0qRcHel8V88bWaNtqZox/QmzzzLxO8lMLa9n3zpE6T4PV198Zx9SWqypsHWfxhD6ZxVVsNx
OAV18zX3PKi4uPoTD+gd+cbWsDG/NR5uk2bR9BFjfuUmjmwDCEzfwajlUr21jiZE5CQPwsJ+PGQN
KFe/1qxZ9yH/RuFRUBLc8HXTHMD2qhFBQqx+lJhJpq1pcmeD4Awc89Vo2rSO3MyjkjoY1hGqUYoe
Q1L1XzXywIz9nki3E1YmCI/TSfM8b81W6+oDRn1Z/k7mBYjDhdMoBT6CpWWooeIPqXCVtu4MVUYb
HINE5ZABs/Zk3q3eSDEOybblcZikTHYbb4I+FmJkkgjJccm1rLcnujqJVg8VEBbHzOZBPEDM0SBN
/GApng8a1NFAr30UfxSHZwZqzmJEcEZnw0t5poEcjgyPYu14rL3H7JXxqoLPBzEvvYgrhsqdKdZV
mIESTosaJ6Ssc/GcGupGFJhcNmxyV075i48ovcHVXPT4EKqLUS8Twzl8oqXT+RLXdfSKnB1SONWb
duxCVcjJNKN0rKbTpmP5VwuFsIiQYSEhllturb0ZXNK6KoYbd8eqaWZTafuGvmdmSggD+QQufKyh
tkCcAOGazIVrVmVCLDKFXHRxdvy9cJsMiWgZ7g3iVc4iJsM3C24iTuYJ/bNhBjlB9DpLnFZj8AKA
VSCpaWjiW37vPDJuFHiYXDXyRBsR2G+HLovdeHqnRaYcn9eHtkFl+ALjzY6JmmiO3GvnYBDzsFN3
ehxYzQMi44zHH4MbUkWOx5z4hBeyfC4KpnfxwYdU7OulOWlsRWp/UmSzdhe6cNtCPXJFsTuCtvBc
9XPUsrw12GxxjsYpnlmzf28MUagr3MWvjhXDy+kunV10s45FqxtaUh8bPsm2nJ3iygfkU4sCuTUh
ZRRJNOeGULaMbsKODOjq4nw1KTfvwWY802gzYnPrhdznUPXNEunXy9J1fVtfC+2YF+AC/zFs1Tik
53qe6sIukviJnk6Oza6zbYWRAfaovkadKiFPmhaGSpyaPD3eMQ1MJ7qG+O25918O6M/yOADMcHSX
rO3EI/fWoH7hVH02xrCcfn41L2yiEA+tsKk385/1gJd3IY8V4e3FjI+3/I3vW0uSrwsGMqrMWOsf
gkN6mpnQImw1qb92tqQmrxw7j030A4/IwLmwUWI2fC3N1oHNdPpauVODf7YPImUi2sGeOhikWUwH
zTmFAy7562+tUhl3mdqvRUcQLBqD78Ruzh5/jzBk0rZN6egfmBc5F4R2JRCqjdWhwEWTpZwB8ntD
vgJf7jNqKVv0KjrT8+6zBcLH+M/tE2PN3XaqDCsKjB/kULH22o86mFW78OCLlAXSHFqeB9Rtl6O1
zp/KNFfS5MXlYgHjdC3OZB3a6ZOPT5FfB4gdnbGfe6Oy+Eggl9M0bqQBooRhciLGbU2P+nrMJGJ3
ZclKzdLLxOeP5x2PhvEOu4v6SOQJfIJ0xPW98SRJQMmRNMxpF07qJOXza1Ztl00MAjlx+TYl6wtO
WU1/Qey0nl7TK4Yvo5VLXi7GDEAwl3zLQNbGwkJkgSm3EbyqHYq6I16lyjDMIe51USpeaKot2+YF
HoNt9lVUXBfmUnt5WE9VfAsAkF3In/Gt8VJV3CM3e+PoXDR40KWKuQGtT3kEctix0Yl2AFWqnRvC
EaHEBxlZVpFHf/cWgo7VF03P8LhWRRyKCEpCc3RYZBNHCfCuNS1nOpZhzktdsSZk0auYyCj7NGyT
hnygyDSXn8jRfUQTiAYI0Dh5X5kioYLKOh+IeoXibvLnkvMHwHzYZWI569zQmedZMwjbigNe69px
jcHWp7h8tMSH2I7M3TSgj7N9qkbjolswRIi+AScwUUcOEDg9uo0pw++TUJGMXVPQxV7NhhXL4PQ9
yt7BpvfuuwtxlFLTXgrWMyHcWgBh4xKt6AUuJNuFYrgW8xWQLcuCCmIoRsDDPTCnD7utc5pFFUz0
jJ21IKblxdIK9r5GuCDp8eHDXvRcD8b82rJT10OU5sNzvOXKmadCZOMJzB/9Mv437oqBsgPqLg1T
rM6KXZzGO/daorXPkQlUPaRE/AJaZPg3SrNRWOQSCOuVRAwJUR0ElOFgViDXPyvIKeOXjA1N+TjB
4xoFBPtrbOAyOzIy9xtYb8xLkY4081AoozUXygGC+0B99WqruXRkx2eIzOoOcrCPk6AujhvSPrkl
vyqKefi+byA3+6Kxe8WKV6GL9QsuQrQQ5Mm8qIB0nBHrQWxLmH5reMs9kJYfBsaf200oYbAmMx10
l82ukErgRaUMu3zsuD6Pb7S7Pd2luiuHAe3puuIO7hG9rW7zu9gfXu2iUrWqF8pWEcxYJXj1wxF0
ZoBWcFpcWwsjx3oy6rpNF27Vxg9t+3HneGyklxF8/DO47RVf5j+P5xwStmdfxXlKAbpd6hzlHuWX
oyAwsy7jCN9wFOjBbMAtR8JMXHs/KIr2PY/NepLVKH3S3NLmDbHrFZkZkDfoYus1JsQjXEdvJU/9
JxDUOOHmmfktYfCATvnvPz84aq2I2F8L4AU5aKFF932IokbBoHf8l2CEpvV469dmLf57WWGb1YhV
2GXPWEHwxqiNxBWadvGrou9hw6mk7anQlQ+d0ZBs6zMgDWbnQ4lWKM7w1if2nlF1Ng/Rew2U9Gpm
IU4+X4Eo7vYJ/KEBFMr07MtkX2gpEPFNSQHn4mjYzBD9lUt+/WNkvoWB2EZy20lrtFKqyLSomhWZ
GSOGr4/+OHAmVUeL4gKrDET7CJSUJZ9zxq+HE6EGPpDatxc5oy5vSVKF0oYmZGXeiY3xoc0cU8NN
I5drKPipQLTnXriL6gvGGpvhHFh7f5afnbXKy7UFKhHR6GwN1Ee92rx9u0RDVO/xLtmHEozijnuE
kz2lWg+Y5Kn6OsqKvO5GA1tK7SOQwdD3cidjQULV1LVtR5mCJwoQhooZKAZg7A1aPPSagD9GBJkU
Jtnw71VstVEJIrLV0E7WM4aSTJzubSx7QYHmHVL15L8HBICWvSzssTe5hKLn/IC4obU51uAculYB
3T8tYJ3KqEzxQntUYljqMkzUmEk87FWQSLHD9qu2nxz3ZTdWd9TVVkxVTHRW+gsAkxTS3R+oP0aW
dx2XZK6mkIcproGZ4Tj5eRwkdPsPpecS8R8wjHlGJPHjV3iguCtyXSQJNyXM75fb4o5Bv1hAx5XO
27X3w42kMuKKGkyGIWw7e+RqOXDCcyuorrCuVZ6TgU6VBD/HLWZfjRjWao+s1FhgtDfMBNpcTg6+
sC+kRaHEUKx6vNSZ08ubbGCVv8Hke4ckYmnknD3g9gsJ+z7WZ0nroL98A9mw682Nqs1mNCddTAPR
DKNp8XCz/rmi5bkwU/FPpVnKSghjadremoPzx9qIk8FkODOj1kpAn7VBI7HcgtydC0E6QJJpQZUZ
8aJyq/HGnkGcLbs7LIcmOY1vs9ks9onr0NLd367muHyAS2KhKih7ynK/dmQRjYkgXy4vIJGmkqZc
i/6z1gEO0jIFnfhWNSEDlr+EhqAVR5w+/IH8RsnJgMgDhC+Q/3W/9MtmyuP0g70R8Y/IwfvhUHmt
uiRTO3GN3tcm8TERR6s5at1oDJqX6Z6IhfDZNgpCdCCKCr26it+LjQfX8IJGMuR7no5VWLYZ+cE1
GH6H3qqlvuE6TUqZOcCvWbMBaOQrYEqOh4IIMBWk/2nkpjGgecIaxxqrvteYxal3tRZh334IFXTr
O0czqLMdq9YXHy7WT3OMKLrND2k/NNGV2Md6u5yKIYRxUvm2giIX440fS7R939tlVSsOJs0MKVya
rCuKD7nKno1TAJaRdB3dkqW0tkzjlnmPaAlWxk4rHWh64JwZhtDypzRYByq+eP77EbS7NiGIe4CX
WV20gwE/7BVzx5EmuJjELdpNFEtAmBzHj6QR/EwsqvqRofAllVa6VlPBptmXWuImVcIwBbDtFkxE
UWkkWcXaLVsqI9AVcnVBE+NY7dm1tbbjggTepPO5veo6EnIX6btjK9/3fatcH//nyWMJqqS2pn75
W6KcKIW7umfzOTD3FPPnbAKA4QATYzY3OK6nZ1xLeevILntkB/sSEj2X9aJL/tx4J0H8KKeQCvrO
fMqY8szNbmo6icUhQQMknG52x5v0qipYkmuRSLaGxvsiumlGmrueMKxQyqGkq0pFPzHMPpiJn5LB
LRIBLul4NH6RBXjm8zqLgFZGvafFyPEs7ZoObzrBpOgdhmEbD166+AMQ9bhNrbboPSIwuMX7O+TJ
Ej3gkbsambyD5LxP7A00MoV4Gtnob3Zx7gfbupOnFWFcbz+GpOmJ991dIPiQtS8IJo7+KE7AJVAf
usMq6qxlxZuceleJdxhTkUhbzUw5awh9Hq1T/Oqk+8VSKDCdNe7Ja8DFTHr48P2utvZtSlmecTJC
oZKRIpRjVYcV2kP93UQI3aSGPr6ceOt+SjNeg4L5m2KMDDKQLpi65wv5qwQ1E9TBx3k2b+gq5fC5
71hrNSL2n+VZ9dTQOF9iiwDA0dSVuXx4M8dvZPjz99Ls2oEwHTxVhbUPGO+GrKgZM1QHHEnWcKA3
55J/6K7cQR/5sNabEU7WMWZzBr2mqLRqax3k2OSjTAcHtNLFtAp6Jfcjdl0bAf2gdd67nDH4G+oY
eiUZremwgn7ou1HmOpsRED11p73lasGBuoW5l3PzjWvuPaHT+dDhLS1nbNocHuFFlFxpcdNUfG3y
St5MsEApBzdd3lmmq5bQ/fO1bhzTz+1j1HcOecO5ljVfytRHTBdJlXhnEEw8KZSnoIh3dNd23MGH
rSBKsykE8FsEglY+lUONWqBpKJg/e7pfVyK7ZqL4F4dzhbBJUFoXMb2KX/DvttKYmzw0td7PYe/N
9NrVZKlMkx70qzr3/ZLtVRkuwLdev54huwDsbWIm+LR68Bvmm/1BtbB9mvcj0Da/G1nejrOe8X2J
0AOZWady8yxh3vL56Z3geNp6WIMKaonL2IQC+TJYWDBJs37VoAwMBiiOhWf9yxmSgzknYB95Csje
GyLm+wj0ic3PjiEYw2TGjWBQP9gnC93vIodh724tHabKBjyjhJj2jtEWNrjQ0COzpkdo7jw/Yi6f
yPbkdBmApNXd5c5pDIOZNNPl+qkgKOoq92M/kVwn1Rs7C5QaHMBiCXEB8M8V+beeUO18DMA6BgrW
luhXFM0UxhRp4+umH333nBtLR9udwQ5M2G/PHZhwWKKwaSHEY3djjuCRbt7DO3E0UaNf6Kt3cxUw
KWojY6UvPLkVc5gxhteam7FHQ4OAo2jNEx65VRtIYcM7s6NF9FMR31k3MMEd0TOwdITaCO/QMu9N
p23kDwO4i5ShAxDamEiIRax7UzYkkB4i0ADd2b2tm4ubxXGU1pMDrg7mGK1d0Btyn/49JRE3LsWb
IqnNUYwBvGyl7BAMjWoKKPtiQiHdI5ELc2X3Z8ERZwl+HU/r6wRHDFLEULYJrmcDMRrUfeCD0Jt4
BtgV/8d+mTq7aAPYADGQNOfKZnpsxs7e/5aUK/FemBd3QMBzp78Cs9ZLn+CfC2nBc4GZgCRGatmu
cIdUw5sq2ntofOVK5uEht++yI+evuCgD1Cxj2AtYYS+SXBxrWzfs+Yrj4g4dPK25ZAamnN+uEI31
AJ8o8zqY4sxRd+UxCTQxY/jtGZFfz02irvVd1KgVsvLZNMkfQmFQBzO1kJFIfVu5pa7BG3MI/EiK
ptqbAyYZTKfKE7Bhun24iNrh2UmzwVevfvZfpyjrmCK5gGARN+B47BKBBl0yidiU8by5MOa7qzdv
veG14xdN+kOiA34XHtpjKMpmLGgXqCFXBq6lh965KOuwrfP32MpoE+2e+aAUpz15G53eORrTf3rL
dP504sJTAV3zgnogZMbRLNqJNPKqrGUnCU2fIiaqt74HVZpDjFVsfMjADXj7JPzBAWNn5SRI99sZ
5nDnlw57jONC6s8HBDBQzsMgrOWhsVwFZg6S2YMGpgp0OaBGxmWaLWF81GRdyp/RbONyKaAEFNHn
WI1uCGxHe9kLqQBKpYR2ZkzOQkfMqCdHcRysc63egBLKNRGIzYVW1fRj6pWdfPJ5pndVDNBSxi0p
iz2ujOWnn5FsKYwdDe+bSE49jEioI4JZAH2VWZQGR9PU6lr6vMYmrqvZ0nOzfJKRFXdUnq4300ey
xoh44WfKd6WaOOwvsFT8i6XycJvZ0bkZDCot0NATR1J5JwAdHXPG4BTwEF1O6z9o5Gt5ShERHVlG
Vkfv4f95xRF8kTlTgGZ9YD29dn6J7XIVWoZ8TxRPcVvc9jBC0dfao7pkz1DIsitDQpF+ZT104Hae
pMbwiqyccmDJgYa9z11gNBV8nB/fIDLUfEFnq6CsVF/EDprOLB+cgaQlASnBn9XaXJkBrvtJvnQm
01+g2HpHFaKSjfqEK+yGnQsiAp/5he8WX8CXVr+c/IYqA218cGtArOj9RErNNpjF6bmncUIU3J2w
Xuy/9JvtTrT5yHepcd6+rhXnpeYeeJk/lnNpj/UVsm+ZlFUjOFZcuQ1mEiQlGWebtRs6HuwXRbhW
g0mZ7hrvTnc9oRfn8HNckv3Evs78xijdHC7JdIGm+R+BjoyqDogTQviA4CXsb4Cyp/PSG1PjJQQQ
6pKTmpAc2CNUHHb2Ln27BZDUib09qed2dPz6TMUe9K4+GdQgH7kg9r9/yNhrMYaGxTWJBhOLaAFY
UiJEQ1oucJlIdQJ+2DqWUSwe62Zy1s5C+ZLpVMJPRIgQzqKuwrpztuefHuhFt6UfkTpXXddLDvtP
BAOyJkwjbEAvDiwHhshopa1f1sjKUpOJva6U0C+u52BW91Gr4c0QnQVCisGDsO94NcOsXwP/THlB
m/L/vX2dP2rS1KtTPNa3CRMlGQxu+3ggYvLsDVpqIGiF0vhgQWIgHnGmnEciO88T69uXmzU5qFJd
sBC6Hws6Ua6SUA8YPQ8xFYFcQVFxp/+aRLqyTejfVA3+I3lA7tLXAYTBpIhrzF4t6BZRGYvFzgz4
IXXNsFMy4HlY67iaYTDQ/qS3bDOv2KAmebBSbhgUDWqw7VZJeP+fZZPDU9nKVx9wyRA9Hk3k8lPD
9Tb30mQ61fwE1E/KmMAa8W0jv9a20itH4jvUa7FhqDx1Jq3H1Mgu5XGK/CUCGRL34AQAqhy8taaY
fN0au70dBusd8aAT/NbY03gLGGuMRSMWWHyAHeM4ML4gEjc8TmXoXHv5aPi2YDRvv/YUnxnKFK2f
tSO+snMbti7TW/G/+mDvhVGfIumsMJpVlWjvrimC8Ans+G/LsxguHPAnFg580yQi8NVxHLGBCqtQ
h+5PYTfrLmcpCI7uJ7CYIpTeh6OyhtRlHPQgurkMVGkjClQj2FQ+ZymQgFu8YBeujCT5H+gKSJE7
fd5uMBdDFCotC3yteSSpUu9nD5TzKLrR/TTMyTKO+X35H0D0KvEmodsBG3WEq0p/BfoU1P+nl521
9NmjU1RP/JbmgNyjuyxcK2gUsBl9jOjil1NEeSQhyrvnKxhwP9OqLi3FgS9MNUkSJkJKosp3Yucl
gxOdxA/zQKQBMYv5LMHPLYlKGxGYzlZS55Ga2xQPHFwWNdNmATFaBUZFuLgfzW9lJzfdXIjZpyhv
Y6s7HfzQS/CJQ44AVr2hymoH2Y1pKTSINF6LMvwA2nLAS/rjoqdGEqqAIDBVgJJFcYgEZTVd46EC
/o8VbCe9iu/2uzJ9QL/wTrqM48CiSZl1kF0xrFS/K/PklJurXP2VuRCyZ85FiW829pfRAq0tewK8
EaqYQ6fmsyMC/dvZ9klrZz2GwaYtCQt3Vvp32/HKyU7eTsm8kqbGFz19K+7q6kJCP7ovx7m1/gxj
4l8KPbjPw92UEoBP3tr4vvWP72+yirZ/yieLFjehZL1q1qRNESpKW2HihQBFZXsQqxFgkE20rtfQ
LgMeIC0VrXjoZMZKVAkjsKTRWS+aGq7JL33rStjkVqf6n9OwI9BNQ42yO3yWR8zmqvSjXqwQp9xk
0V5HopBV1mNs0a7E6XEijwcpIC9k0rxb61wdvOlIRFG27qlTU5Z8lFITRv6JEhSINY6fdHNPJhi1
/t9isnRcxuBa/hmZEn245oCH+pfYyVUdEbdvk41jXJKea3nlVjTbK7VyAauB/zkjoK3rtRqhzF5d
BbgkhKOwkpPwfcfI2h/loQcrgobWzO3/Wv1knwDT13bJ6gy9r/uCwHo7/L+NN6Pd9lOFhvsOhzgt
iLBXXBmu8TGcH8yo84bCH5VuM7TxuzdRqvW83zY5e98TVOU1/xyiVB8PVnORVFEPIa3+4Mrjgz+b
Xziq02/FOxNiZnwW0W1SqYN/8+ktz2Z/W00V1vz3S4TaJQYZ+dE/TXh/T2jKZVV4GjM31B/NTDAF
//8ymPZ4Q+RwHnku3m66rAFHOXRmIQ2gBCoph0Izbk8kSgPFuGDeiosGswYt4AO3Qa9+a9vwGcp9
QOEWLNu13MSh/txUW1z0BFY5yIuD91ZSMnyLo3x54wB8Sf8HWaI/WiFXZtNMiEUKG36NXL8vGPKW
aJvKEXK2D9B3enlrmW+xGmLC7sWwgV+oGgcspmLgbuKnFPwld5Pjzs9fRDzJUQFx+q4bkGXeUTkh
fXzJeiknqz6lBM3X8fZB7bEoLWiEcvWbVfTfnjPXfqFoDbfb8Lzks1WX04k0xrOOeRU3E571asnz
cyoyXfbNvG54YNePxiPlnTWOpBOvvvfcFkPrkoSx32AggQ7T6Dd6oF+d9zZtokD6yKZemV9foQ6B
O6Zqd2qFcVnCPerB28QasqJ1mMA/nhy4/VwC8EpgLXeGrSu+Gkbb+aLma492cAEh5n8eMOzxj4WW
EN259j3VErY4fgYXdBU4o7uc+AYMOOE9uPWYZtgxXx67phnEwc2+UYpjUw9tkT+dZumm3GcgqlB1
XVk1skideTllKbGhgiSi5IzvnKPCUHHGWlG/rY3XDmTp7iEbB8MrQ9cFTVhojl/3r1JM04CHPkTk
0+K+kimnuR/v7UZ9SBDge/x8kyKZ9rMVzpte+mBioXdmrs2VRpmt3PqKDFaXJ/KMGyQQwFf71yvu
ARdjCezq0X9XTrv5KRkbI171MgZWT7elrZx/UkVyCvYsZNnsUSAPtes16yYNBvmZItXzER+nbm1W
p9wbyS/8aw44mqvZlJ86I/lFdcRl7OtkTosCVP4+unF8uNp7HyMxFJbo2sdBXz5oWCFusuU3t7zS
coX6zVXBU3RVnThcHKXpwTOCU3A2nRFyVDiTBcjKqAQxMMjxSmKwLMB++Yw4BOxYvTi5bXU1iLJm
U3d7Ms61E4yxRlQQrHxbHOOoXoEl4EeLr/HNndeo/vqXQTYaHGtQDxNFgO/PQdIKTvYj7LbS7e7K
gi4JwGY4rJ8BZfOzx9RpUrYWGnM7BaWH8269g11ceFHWQMc64txv0XpYm7/i/o0kT4XUNZ/lrui8
wpuvmhZcXrWoxyptw8dNrc9HurAaxs8PlU/wi7bUijltagbweSSKPy1E9XvOy/RgM1J/H29MZXPj
TjBQNMCecWluUbntYLlQFfJZe98FK1pTOXXIaniMv5GUSQq29NHhiq+0+Qyj4YM5qjhruL+9VcLI
ZOtp9AHc3dbybk1iWIL+r3aKoQ/mFe/ZNYn2Z8t0bFJe4DMzfDnxLCXZN1PLwuThZ/k37egzxGHQ
9Wh+SxnHL5IxUcPcjXGjv64mmNuMZC/84jKTkZ1obSgpOg4b1Cksm5G6wns7TlpuCH+7j9I2lQf2
lYG8/cPh4/UCkCFYLIZiJzxpFREDN3iZSmrBIx0+b5S3ZVpravlA1WaAImGlgvEJ515gzmZ6vL4c
Ex/AYnY4hiRGeI3gPAP1UbUcufXJXXkuVDrf/1r1OR97IMSpCmuiI3ZaRG2Te5wJsIeD5HjKc6rV
ZRf+5Sfd7vkm6upiZo6i5Q07W/94k1w0Zj0+DLPxR6oguVJn12SKx7xrKOUI/MGZ64gwWeQ9fTYq
Mczm1IwH4mwd9jlPA4JSZWLs3CcdRa+cX/a40K+vKMEGFq+5FL5/TkHt8r19PykexPDncLCyLmkK
cu1WXczcxf6tghB9amn4MPVvCBXthWzrGX5+lyU94KjeCfktQdoh3x45PQ8ucxxurbFVTQ9X9Dm+
hIIvDs3+O75hR/Dqf5UZOGKd6ToCDv7dsjXdWP3M/ZAwqIKX/B6Pr4FpEyG/KkdEYVlwshXHixsA
W+A02ojI0+yha3guW9qzppnIUKfczMnKPppnPG88p0ILzHU1z15UTP+EvxudKWctaWObCV2nDnRq
UOO8UmWLMPQxkLZWsNsWfrCQujIRmAGUDM4ERcRoFGhvPIYg9bLK874DuoF1tXwuDqdUdK0SVaXP
+Ant3qqSGExF+6QnFoSfFq9lBZ4+Vka8du0Kr7C0szObA9zGwQs2mSAR5jpsbN9mrJBCxX4J9p/E
WzGMsAWE+stwSXJVZj8GXFWQAdltGLQ8vIqteg+klsVUW3d0W9H50B6BSoRMRNt6pezBWTR5aDN8
oI6ypI8O3Op2FXDfrTEq7pCjfA+/T8sGyctqcLe6mL4N2+mb6qBAc0OCaMcr9jmLlOAVgScfov+V
eJbmzhzP4y9/ecOT9+gXw3Gk11138w69KK6YwG1K43NK7L3BJU9z2udha609uQJwdIjpTZj+GamB
4w+G9AgjDjqd1bo85GGZXooWdJsT1j66FaRMWNW5s/y7467/5J1eZXX1JByhwSLo/gGUx4cbmgKu
C/sxmFS2JJ5L2ufawdCosg93OPecBwgQFIIr5O7Lz6Uj89RD1lUWMfuJD1fUP/dCLJs/Tml3nbZB
jyeBtJdnmiO79TcQBKiBkxt4LCvcDcu3ditHMb6QsBtsBKVr0MeEEQ96u8/40BZH0myiHWi4Dz5N
K680tnva9FH5unJXTh5Th+8orgIjPtQjEcMX5IvjBti+Y8lmLCwNBZtOmla76Q8TF9Q3omyacnCG
J2r+SuC52ruw42EwQ4GSnEZYEoWVhXoCid+FAbRmN/fzmtn3SxEpv2Gk7hylwWwYAsaZH0a8tR8h
ir54BGaJ4Lti3Jqu4e/ClZCvlluEyujC2PJUqKpqI/pFtmlBPf0xsvHSxaVil/MnvDFaOq/mpDjg
vmBkooP3aAUaQ3XWSQdzJxV4AhczfyLxzs7i2UgXqo64z1s2GiWSVrjwmqYc/uLC/wZuGpiXrXk0
7do7Anb9EbwTr2wxt2/Xxv5CyHDYlSIM7JVo7geRYwwK/uzsLSF1tqYrAPKD8KMYd/m62StcyZt2
lo6sb0lFEQ2grwScVT2jmwSxgFIpwEjHZEUoqFIsaEcbaUT9PJAD6xJx3qGNNFZERkfjRwx/JpOE
JogWPTdehxWML9zrBeOCe23h89tceE6Q2Bm3pjd6HehkinPrymsNtzpYLgsqXFVvE9z6mt7okDV6
fGWrxPkEDdd1stuBsTvmIru4vCo2UPqEwuCTPF0SmKTtWI6zZPFuYtwALWUopVhhtE78a+YR4e9r
vYmUsQqHdiQWVfrCB4Kj66HInmlq4wm/0350zjETKMpWmlS4isoXzzUvRUzEUuywjg5YEQkEqzqG
AqFUPJKHFVNeQJTNn/1VzRk3vKl8DXByfSwdO3RIdaPTAlxHi1QeGEgsxKvGFZrMH3URYpWG9aP/
NKXarjGBfJ0bGoUmRtdUGxRtNNantu9gkCmGv1JvQ58vKazI2HQ69ob+PzwAg1jcyPa3Gv8cLHbK
0zTVhqbz6/HfpwNRt6IUMArkz8WE+nRN8wSj8YbEv16b1CgkJgtl0XYvdQr/PFOb4bcLSbBPPtoq
mKYE/iBLDJlAahHD3GvC9GgfsSM2v4XplbhZRWNQuMyl4B4Dms7jI0YnWCPGzqxDrYGkI5QQQ0tx
mkSceBeyhkNZ49+yE7GReOEzv72X/FrKlME1RKvSoWVSBMtH+KdKAn5n27rIH3U74UwNCrxqKdty
zU7KEj40Wcwo+WFaeQ56DXgXkv7cXw6d7DETKivm7Xfyc5IUlY19jfL03S7N2pcX4pVSWr2s7a49
C4jbeMtzcEi70uZfT/d0gRerXbjlsb1YYHvCMx16cU735pMkoIkjuhwVdYTB3jQjBvy9z6K2AzPB
28EFOiiqW9V2oXwQKnIIYEqnziIGgIaxcip7DwjVTC0dDav9gA0l20kGaXqtK3w0BWq9pZSaLb6j
hqGr+TW+flW7PKGI7jULX9lXKfLEKkDRoXEmvdaO3qJSchyF3uA0/QAadDIqQXXD8f4rjdu8009v
4Qh33lomHswmclJXpQVT11+697hS3fd37MvQ/oK6HUXKYGlF19H82IQ6i8Pt3BbcpMoRkfRTOoU7
YoM+4cZwFh/qgpko0N6YfPuj8ruOW2Bp+MypgeuDgwc/Lq+fR4N9eMtYumWMnKD/eCge/VVWHupj
cucT6h8cUHkIig1+l4c8YKeXh4IYg0Dqzbt27iVzajdK8wpRxLhraidFw9vFhUZQ6/466HBfXpvq
VaF2wtrkK+7faiJGvtkjTsk0/5UbkmGlMhOqmKbfSwbRZQQI0gfET+0DneVh/m0+pppVwPYR3i3O
rVpzvx41azY4PSc6c5Qfw0bKB9BCB+TFPUfTbqluZiY2aR0r/sAQa3DGT5F6Dd1+7nkvv9zZXd7E
Eq6vs3UK+zlIshYBFbVX3ZUtG32njB7Vwuenn3oXAl4F9FUshUabM7azlwA3CbZ1CUIEvtNNdDvT
OhzXgTaL4uop9hYApmrqKz9KbcigEBbVNiU3Kj6/dCD+hp3is8wNL/gJd5JaMi8PeBmlAs5af1dy
6sdv3EWd7Fz1u9WzQjkuUd5cXK13n9EBFXPTAH3FEiVPlDxrc6fuZf/7xHgg9YqhytHadZWhMare
CRO0CVGPhu1nEM6VSLbh3WTewwdhjM6KD/RuzD8/Fkq5PjGH1YrTvpA+iLB/P5mXShRioumYrgao
QfNu37oinDmvRQLjAStav5mRR8egxyuPOBG74wRZ9R4OETfEvTiAqLhEDUZlFPL2TAJhV46amFjq
vNdAfGhwLWxJvKJuZ08wlrNMq2TX04XKzR63SgPWL/QjBKZrO7NUbyv8NcLbmJlWjyd6OwgBw8sb
0lelWO7eEmG0NGg+EAXlGpXQdhUGy7xdFtkkSFMWlGyCwAUkvRnsS+ppI5sOE8keDLCPVdKHzFZE
61X2IQRZtfvfAGCbrpKgkSUgErL1FibNKHeEAUIOtFlc1srepErBil2xNNh7xPu1CoDldolTke3O
zENT1UhDYk01l47fnLqbTZZjEnDHdH6PzKansIockmE/DcLkNGPs6MLdhAGvyB7FiuLn3LampTMo
RcsPH0smJQQ33dhOUnXcHk4Ft5ZxWTnpVOY9TK8XFVqTrjlzd/ayRMP3VvLsNc5KaH5eyijGorXv
RC77l9kzoTpfItb1r+amAKOtZIAhhnx4Xun9N+xo8gIEC8TuptN7xzBN3wDvW9sJ1tXCyY6E/v6q
3Gr8drwcTwxa1hXeDsqaUPKHbp7nv0LGfwxQUw2+CWePKBpwOJPQQLGAtAwyLszEoESeIsZtuLHs
RFQqQ61lZyKTSoZksJTE2rIEdIowEdXQOFKlcvIFJ/dRXulAeVpjxHDe4yKbz6oHi68XNidxgAKf
ZGouzLTxp5NqDoEVMK2IMtHURWeopk8oUdPRAU1IXbZNCv+M8EMEscBD28VlLZd0bUIgVBtpyRRq
8VJj83rz1l2hZglY3Zkel0AOyc232913FcgMxGDgEDzjCYf0gKNH7S7LyjJZTulUmW8R+tajtftL
kDsQf5kc0gXT+3uZ8rv/WOVxlQTk+NprjcfuRFdKLWQiYerpiJaCQUUw6XSndKkQd7qn8SYnpYXt
IvEFjsNb2Taq2JA+evaL14zH3bHQvn2QsArjtltMF6Bm3zYVVe1u/Ra05mOttiXcI1RnekxOqJdb
Lztwz5F5JGRqEolLM4sSz0FWyHyqk3miXKDc5VvazhxFeiv6ip6SLTACznUv216wYbtANdvc93OS
Y2CyasBEqOzDVskCcuxwGQmeYKKIK4G6pG6VKTOACtVfIuRU5NebZrWYr9VKgopL+p8X0nUJPa7w
VV4btdlDxKQcOhpW1oprRdZPoS1D3qKHOHFdJSHHGLuk2GIY6d/4iF9U4W64Fvr3+5uCIe/8nw7I
mtdwG4BvnviZKtHlirJbiD+pWiU/3lj2JU/xZLlGYAmL+iMRN66Ueg44b0D7KWrhSBEzTeh3EpXS
cLjYZxkyaGxN5zx+aZi5hPBXDBOvoAqNJ5rt54ak/WVJZ6rfNNc++Lzvg4jZaej7Ae1KQ+PkZ9F6
O5nO/QH6wKvbS7wBvOl/KNMj3h9+SpoMZWQGv+sugvtZ2fP2LTRMuFhd+pXaJP+IqVF19auBBtA+
EKDd/L3dZBsiRWGyWmnQeHZHbxG2V18cjy3Xrtt3RSq3HJdzLjhhuVOEvvGVyvWPZbnR+gpY5I9M
3Lf8qpN6ppVkKQmThtR87odsLUWAz4X+vRypSBIjmjzkggXSx5OS2E34Oe3P2nMV2brUWG59QiJH
4Dmk81koZlds8+IkfsDyEjUU5Wdv2myHiIuQX9A4wi4Ev3dWsMQb8Gc0aJwQBXxS3pDL0m/euF4t
NFezpFkFp82DNJ3tvOboHm9W6lcN9Ah+tmIX4xewV+iYtu7hF7d2tSdblsODt2Eth1utscmxfc2s
pQsHBfunkclCG5x4ixcMViq3Vf4gujxxsZg4BB7QVc1quRbHXQLByAd3Kuvt1rjTyGHeXoIAP8bV
E1S0PGKxBwPFU3VRQ00JimgyBeOzn0BWoFSbeD9doH0Nl2WLFdi/FR2SyqrhDQy9mj5UCo+NES5h
D/7riKfBvEGz8bPbQ09sLYIfG8CGM84+TaR80d1gPf1OLL9lNf74LZRkYPL0xTgmn8l9Sg7BV1tn
JRMPO9Gdpd6jeGpRtWrPf9NhZ8aUcqBBy4J1e1e5l+1EL6n91qmXC56WFCQAi8vFuCYaGJgkVLCh
xCPQRuHq6zFXlmwRFH4nirqJg4LKkbXfN/uqq1vAn/OWVZvM16tWu5l3OCYqzfRoJSQz99HmFG39
di5GPfgMQtpTTmQQ9bAfuqBnKxjmFU+pcbzV3P1bKUdeVbG3p+Ziw69tRtT8h2ovCuYMO/WZ66tO
yuFat9b/3MKKUpKxsHVeBiQEvWuhhp4j/P/ICngfOB+OaauTTyvRz0L/XdN56w7ma2A1vGdQwHtn
u7mnWZqY2cZnWqp6qtXhMq0MU7hga+1BOf9K9wnkonMlEcFI/xnlonLQZey/THDXPtIY5ghHF+it
SMQB9G558Zaa1qANUGy44hOshMGB75pZjEJrKQ05PESJeKq27x/xcKt1KCtZQZ16LSSbFTHHyeUI
N4ilIJNFyMuDfgCewMeZXMdz9J6t4EqhYGpVd4Va/AILPBKWGjm6ZtkGsJD0SzLgLVXu1GfIQgDX
n0Io9OqfdC4NmcHAv0afBTiFzr/p3QwZLSNDKePfGFb+0wm4fTRVndgDiQ+zy7AnTuDgI6Wm5zi4
hr/nrMTpcw28DMFPn17V9JU7ljQ4u97zyJfCVNGtNi8le3oglRghv0Y8is+ooI8DzXJNnwfkSbVD
R6x9luPIwlfCEDBd51181b3aprmfNcl8p7sH78TPlJpBXo9xBI0yYeP7K8chW6+Y3pc89x9nzE9a
580A3tlmUEvZtyDF19JT+nAanUATpt91XM0srhNtEXwZQbMBVtS4N6/SRfRdJw9wv1KcNQc1xzZn
tZJWEbtfSKA84Ztg0DZqCa097CycCt14AZbC6l5POE4ZgjYWYbdsru8peq4r4lAnJqWBEGDMFWNU
jFwoXbeEuWFE/9lqZkc67jFQENC36B3nTg3UW8MG8xmznf49mwyeEsddespMHTtAJm/nNN0gLLZ/
Ouw/FFsLa7qEnQqKB2V4rfaJDo91ANFnrFHHNELb6h79SVm54sctjrw+6d2O3IUeUZFjttCr7qEy
uuYosYnPhTfk12YTQUmrXHI17MPp5RY8+kKBlPkMtFJI3PQtIQJ7KDvFLmioPv2tPBKamfwmSPM2
bAd0d/kfUwJBEMyOjBqkunSTC/Xxh03gJsV5g/9ZV4cM8/Ir5RAMSZSoRcuzECm9LhBMlETLrI4n
cpO3nma8CogadOQipd2O4d4gWd6LmIjG4QdYnZu8pc9gwkhOyJDnZ5gy8Rv54OllytAhcYqZe3q/
QT8CbZ/4ZEXQji+za8iVfoU2pMYxH5e48TfjhEAP7SfutS0l596vs518X71Avn54LSO+XcGL44te
Ya4Nwp+9YIBWlyRL1ZXdiHaNkVyUGYDouIXD6poFKNHelPRtiSrAnxxyipWVSI9bgkBdueri16vt
5a4ArIhiuUIYHSGRC2+y8cb+3NTQznZYe098HpKiTbC2qy2WSt0uT+rj+LoN01L7iqQV4eNmFJjJ
fb7Am8Q2W9PH4YnhH/CmwrBYboBjji2izihCbUEPekH4iFBdf12V8CEgY/axdRugJCUZWmOUD4n2
RTeMMIcWNGXNfzkZ7N4wWHw3Y255bTncvU9YnWtiCd5JpurVpHbnI0ENsEs8CKTsc+HSSwIfXXmV
oz6Otb+vCTVhxZp4/J/wMjWqW8EPH0oAAVuWiZ34HAMewLZU9Txq9cQ5mExMPt6OC94MTJPQWVbq
8ktuReAGqA7c1+ooX9+ctb0QtAhbKuDFrtV1owytL+ahESMWlkCbZxmXnFspzESwloi1gUspG9Vx
UCY/TOx9puvGuctMiqeaLdf405saqGJj18QauXJPZcqpOTjpSD179sJbkQDq+5NGvqOnYnQ2K4XL
/uFxS9kwYUnHsdinONAzRZH28XDWlNQsRgUxTjHPxASZsu9+iBIINMryi5FRoPTiWYwFIHiiXgA1
vlYpVLo0AcslZjPWb6Fi7aT9MlmlsJXCgMiAqTqWdhWFJRsYTzemHeAwjAWholby5kdSzrCSQwDu
3qIw+SC08hLIrFSHTOjKSRFDj3U8KKDDjg+wR8esY3NfD14eD0Mbc/ZlfrEkW3S42HdkYBN0gUWi
AgmUe8VZREJ7P5QkN6CNXlXRsDtuwS1mGZX+Z6+34PDKASRZhyD1Iz8+i+s87z27nfoM/hPB10Ya
BgnehCx8EUuvIXLpYci90CHuLO8C7SYngwhEGNnTMon5epk6Cqz4RBHSmW0UBB4PVVU+l7DgQfFC
NyCGdMADWeU0wDpyRTv7kEZSk1stLwcCDyOi6zN8ZiQHoPwB5pCNesrr62zt4rll9U+NFnXmJE01
zYcBkZQHTeNDorAsaWw09mjT2aIWk4eaxdMpoQsWBSSquwr1PEBpnCIAmOMuou/x3ggK67Gs9TuA
IstSerr3SGTuaUTJlfkig/B94ort+Q8PgRKUWArscHTL+ypLXhC9IdauDUC7tA7T1uk7Xop68Xp+
TATeXYUoAnBfImxy/vf95pkGO96AOMzw+Mf3ClIbkG112KrtU1Rw+gtmAjhfAVIyjv+IU/oXtZAL
srOmlGTuUTv07x2xX73+3faC81k0+9hf+VEMEVtldrkX4ZPd6Yozr/PYcHI4FW+87DrqPICkUjHE
dBMGfu6HqFMI8FnF6wof3VnW43T1kC1XPGcR8OETKBgp0VgbTNbWUhvbqsQGKifc2LfpOx36s1vh
NP4GnCjL4c3k1c1MLb5LStcytTDQH9pYYRAwrvlN2rshyE51PiRBqR0naD6AcKk0K8gPGhSRCi0I
YlBZXdu9HkhUunWtTilteVQu1O+qRtUGj9Z//xIAuaL43N5g3ngQvlydajgWKEY3dFIpOGzzh+Kz
nOx4r2JzBZ2Fw90SvDPaVYmO2xdUvtcvD4Iv7oASaA0ReUKDdULcHQysKEFhM8WeXa6a8J118qvz
zTO9qqhHrHWNCyanCtN7Au1lUiFaHymfV+NTjPbMaYAO9hxmUO9r9G/KOXDBE2p9qSaNpzGVTmDs
tpRXbTJYp3tY/K5fHQXTEQnsNEi1b6KTjuoKWMHy1VTlyPIKQHT1GyjssEIaqASifih2xC8tuRO/
8fMmHA80GxmMR4teXlzp0O+wUR4ZcUn4jOIXARR67cB13D3x6VFnYnvCxt8wNZ2xT5VBrkwtoLye
OZQ4wekYmkBcAiXEpV4/H/ETJpb9wn5xw6JdKWePtrHUQYqAiFYtWnLK0r3bs/mTAxXMJ63y+0aM
3edVWDq2Pk775GMRWbM9XhXMJKIoIgx+UtSANYso/5ATzB8csNmyerAL5ZQKM3rUx4hqdZy5xRjI
La0OYoPj6ldxqbBeNf1Uuv39ssF89pSsCYztygS+VacqMp2072w4k18JnrYj49C4LULYbRSzhot+
yH4ltME7wDIWFYWTtZb0ew56Yli6Ej9T/M/iewaAn6lehXdSt1MrstipWaxrZjIRt0K1MuoRl5Ka
TlLox5SSt/TZIoEQ4VP+vOptF6jL32WPf9YFlcbm4ZBPfi5FVvd35z0paCWkhIVK685QG9EJOPqF
kD+GVx59Ercxs2hahOy8NeClb0CjjFAMB0DNuPLXcQlTUGsVYFPHZhfQOWazTmL/ZBChI1QsL54N
bc4k1c6AjgKE13Q/A17SZxcwglktNE49BinBpOKGOAx3w+wqoYBz9f9H4AP7pjdJvodGGnhkYrbR
xTYTrQj7aY4a+Lo3uhI+l0/ZrAgTd6naTYwDipjaclDPAnvRiP91HGFOvmPfaq/mominVRtb5fFC
F3p8kWcVj1pDikEStAUQUikUf5FAmYmBpqhA7mfgB5HLFpLf8ThIUwmIVUPt9opVxK9zGJumXTLZ
kCgaJd+h9R50bvnzBu7bkr0NwqHEKd4WgLDrL1srtvBj3PVDeK++I623+vlyX/oXCtV41ktm3kUp
v80Zklhlg1qB4Ku8cR5MlxMq15r2tvkJoXbj/0lUpd09WLFo3yq7xxH+9QUzP4r3sNtRD99rGRfR
Z5mWKxDdDe6V+wZoKyw2FHtb6NPqabnAKRhdKffdvm3yhsglLcWtIAP4PxXutcoYVRWH+nXdWcvN
zBAXMWAtMvG1VGMt8W3q4ScvAsRl2rD9uaIUTMvuU1Cw6sdn49/RmNyZKSkB22fH8bNnXQWesGe0
Sqz8sj+K6EPHbN3Javpk3yWPZgaZ3gzjfW74YWB5kw8i7nhyNQw/G3RMr4tElRaXcZCJ4T4MfP35
o513pCwzgxE0fM2vtMzpfqGvWs1NGzQrL+OddYEJXocn/3Dms/Sm/jt0mOHIIL5pNiyHBNxDn8LA
lWBGjBsbWaeKUolibXP3+/oZBg9mi7xlL9aD9k4iQnPNXzLKmNGHXCekF+eFsy+D9rIMUKYOZiFR
v87U/wAS+J9D3eg9Td9x6lzMP5iQZzDorji4DEGK3YRRhJojuTclGNGRk6M8muITAA40IdU64wns
gywbTkJE4yO17ipmPR59C/jI9caxkVKh297rNW/FIaDwzX4to9QDLSbShz2HlY2WkMbtgluvrfLF
auzGq10PjWozQd3uCes6M0b1Fdu4V+OXUVf0EtTDRv9YxPuwY0K6W+dA0eMuRJfqJdsVmVyM4Oae
enMI4U9nvxHQvZQSIL4vnb7cxArAS3p39POQM/kjFeo1rxGnQDR/cl+WHJJWPpCEel1arfGYkzWI
NgTkbRsKWRTt6ahOYbMJUyE+T9D8/4eFIQdOhubY66a5YMZRKZq6b+fImxJHUdQrQ9BDIVqjIPwc
/bd7oOHbmmi9f+WrZUjgs3FjQ2DBeXwAuUAYC/yjp4QLhopZV2YnKMyZrsN7YSFW/scsZxXrSVG+
mYfklONS6oNK+OHkbel1u81IA7mYtbEJXmKDq0AG84Sy+YJjG8DVTlXzk2/YZrEuDSW8WU5XJaYt
UeiGPR4GPPUNuznq0wr/Dv4BgRlwGjKgfW3c4jCF1VtkTYVkzf7W/c4X6itcvLWf43tFaqpV1MKu
tlI7/gSkNFgPlO9lJGiNirOq6Ja+9AWSDYjzOpA1h+UTaG0db2egYTtz5AaLvt+5XvzbFrf9Bb1o
aMV7gAa/c6wXcKd185XbWLDo4PsLD70lDDPLi0IoHkehw3LzBtCTiU+3owgdTHX35DthPERg1DP0
yyxRfCZrXcMXY/72pdABptf00V2vq6paQX4RSSi1/UeUQGmDtZu8r8XvYozVY28CK72ViFGJzVa/
jsv2k1Zae668nE128r/cFBgrMwFnFt7qq7BS2GNNoQOjovX+VGLSQAgIKBCnBb9l1AeX+R21T+sJ
TX9kHqeBxegaBPXRlnJFCbbIG0Sz9yQohQeZ8Xqb7/3jrTXDgygDw6DHLZ7Wh8QGqRXskEX2a/zw
UQ9YwDHf3mw/3e4nQapC+ySVFQQfuLFcxhFrD5YnoTeWLZiuxY8C3RDlgVlJAOhBS31mK0RV+Lmz
EBmAbVeFVXN0YVKVbL90VWpndYsSyKtrmju5iYyzL5lWCZ28vQ7XvG7vUam2e8pS078DwQsv6OZm
P19jDYOidWepELczRBa6NXRpv9sURcYhldUHaQXYZpcUzfuUcjhQxLjfPzV0PdHHnxd+RD6xas4l
qfpAQ07e+yiLbZze9/CPJmH3L2Yk0EUMrl9g7+oIVok/YEt4eERHa+vqgpuS29jymAYFLq8Lzvsb
SgKgGxCSMrgBLB0gV6Lhvd6RGwkYuaX3ZnsFa/ESWAO+ZN3KtomPL0a5jz5CufhT4ZdC5LLX5u6p
F2SW/os+yQGDzEIbex1UC5az57s1bXnTKE63RAOfrYw+NRYxQhbpUQw5BkrcPDcE1M1HNcdtGeHm
tq18GEtdIq6IffXkWYTYsfvbjKuwHQSjx7apA6G6CmqdKuPpnqDILSGFCNWmmId504BY7Fwcjb6d
jw69f7y7Z3HPMkJ/ARWN2b8pgHdQM6/e18iclh+di+aI2rdpEPfjIlq/BQ3nLy1x3QiO3yc/cohp
WSFsq9lQ5dXga/sVwDjPJ5EPKg1tfX3msHd/NaiFZmsDWXij8bREPe2WZopHJQjGEnjyZai9OtQi
WpGTxfOd6rbVceUGWf3LOzJykVBZkppX8n51BQ3km/0wzZhW3l4tVE1HGLJsZ0oWmNxYN6791CkN
XjZRbVzr47IpoNb0ihp6XvoiJAqxPyrk51M8Uv5Y6jJ3x+FA9Iz8QGTvqW2bjf18fORSay8/HdQX
dhybbb8yx6EJFcS17pGv68x8modxZucrAqN/YJYw6sXmkANPg2S8k72EPoHr6LGKIRcssRci4U3Z
oZj/hU0H4wI3nRo9pwmRiYbDkfGbvwP3EUHIsuNDIvkqqc9JDzunQ51vGFnqQd50Z9GT4h3LISFe
Ermjp8QaN3XkeALRwX+GyRUXuCRzgpbO/3NyKuD2c7n5dEWcT8y79Z+rVO3PhnR/NXp8Hq9BhWyN
3zOWth2YrjzfBcqME3sLz52Ho3L4Sw9932cAvBYymg3RPnYNu/0wvqjn+/9R1h8U3+5mN3Us5xK5
GN52JM1KppRuqcVpJdrdoS4st8Z6htEUvsaPOSW9WDyi1rYOujPfzmqzLyLbHLFnBb6h+GokLT29
FeCS0PK3ltDU+OYbcQozHEqpkIomjiA9mYecqK8HATMRRS2b8NOBiTmbaPM9lfEvUNouGH3yW6pa
qiXRBSI776XmEjuXUE1J9irKJGi4uEM8Rhc2lATU20hSunZQLk/+VuRn8ugTUQRO+Yls+fYTjG4+
UYXUxbXQwPxhnI1ma5iZcMG3ECZCp2IzGRJbbPK9dmSMzc+ee6wpA5+lxzRU+0iXJMY7tuws/vqT
EVIbjYMNbHjZyhmHVlqhwkZV/g56Y52JiHE2SrTPYaDTq7PbQN+34jQNzdVpgtff71tlvmcHF+Zo
diUWRQfA+hdEeGeolg6Z+8Le1WBkV0/IEaEcgvsuPruR2A/ER/M3TOawhX9cdmNS9ZSB4GXgJxe5
oydwbcWd0XSPjUG26ea6M606fdhfgM9hHpecC1aZXBsifmFByFVTrMXrF8VgsEsx9Q1HsXF5qKfp
FADv//835yBbmzEgcBrYI5FcWDza++SWnBt4pk0UM+ZKUJSCHe/2RgcqTvGm3+UrT6mUaCTpAva6
aLmV6Ktr3F5C2iRaLY6CajDZ1GScSIoMRF0ixxGQPg/hXwTJaAwH7HX7g/x8lzuHEcNilFFAyzwy
9viSNP3TIEJFYHf9psSLH8nQkn4GmUb4rdiy0aCQzQEB8uylOy31voiHIxSpkuaxc0ONVh4/EKs5
X82Kx3mW3aMekq/4uXkx8a1E5npfqzrBFI1miNyFCKIqxQZUjHfheY2b3SnN4hoOVaqkHhLsdFhk
8rl1NsjMWPwRQ9EQ6omCbS1jXGvNGOyau30rttnjBtvD/5HS9QNFxol1LZ82TRycLFEyu2GUNJw3
2xO5oAPYMtiUNHY27V3xqi6fRK9Cg4GbtFRqsBsb7ZN1zGUkTotn/dmyugLfTOE5qpXWF6+ark0P
k0G9Bz7f5BLHk3yfdyDJtp8dgr9jCRfD8BS+xO+Y+chauv3cOjatZVOiKvHzMuo5sxR2a277tqNl
qnPTeA1kRUbZP99xVxDFOB07jLTIpVNazY27gcoduZQspAn2WF0w8jMeC546QzF5nqEzyqwN5RUh
4iRdzefa/q7lqEA5MJUcM7T+nQsV4ESizcnXT7IU4fCgMlCAsTTKOiDU1L8dqy4wiCyh6QclQj1O
v/oEJlJRD7hxorz6TLwxv6sc4iLXLqHOatGz7+iSaRnB0xAANaZqh1uW8d0K3PurNCIO0qfW6JTx
BPqd9VWibhPA//E38ofUvCV+sswZBW5J+ep3/uHzWrcZ4CfklzriyswQqT5UQaOQXfp/DzqCo0tS
lfMvRzwnVFiDceLHc2COfHaKLNZ86zWepReyLv39F6ODmkHeWbKDk1Gnq9CESvpXEtNGrPuLdI4J
pxasanH7GkcPHXDby0IIvr7riK2dqp1Kiu2FFEPK3t/S4L4/3/c4wk67rFDVkbC/keJxZ5k6jba0
HTh2byq09OYaKf2T9N5vIuRKiDqXowwMLLpqrNVT+wYKzHPg2s3jZwegvpxJ1rZVA9bPCaigaWh/
PBUoIBOTQcN5fZZzWC8O/1NbGGX+0F4OIw+8WBu6D9amXMGrTf0gtkDTGRxjWiiRX2BKis1R4qYT
VjBRW/B255CFTdLc8zdQWmEG/IIqACUVTQJzx0BQjvpa9PNTsgNr7JKDBDgMrK9Ad+9gdftzzqF8
Sbq8qz/cJFNOiAGw7Wsg6dYK1n1ZdIpI9RGSG1g1+H5W6HMh8wOxNndLQPEDhFzQq+HypJMociZi
WqSVT9RWbgKiqj2KJGNk9bvZkrKTcaY2nxuP1drX6+khQdYZS1FMLBUK5eew7wJkGdMxE6LUKwfu
tyWEW7Gi8ADEwJhEIxoxFlssLTS+9RdEIsfuSataW3G1RKgomv70SX69r186lOaLvVEkVH9Obquy
CmqDf6kFowtEwCzMZ7GAcc5dnrhLbQNEEGDHZFE5Dy9i8Csi8MiE27l+S0Mx3TRzaiUrRR9I4NN/
5n5y2Hx56jZJ19ooX8Gj8UP1mVnhlRXwtN/uMs17izT1mbQfBjjvnl7D6lUzqnaZBReqlTyzx21P
orvAKxgBU+iTXBXzrSfhVfOFCNHMM5SpanZ4+cYghqVgxW4SoF+2vymMSvahOibNk7Co8z43TEI1
1A9BovoPKrIq14m/+EAPL114khsR/uKnnweyLSzx5Aj2IJ5tUjCrZlQUsOvpIbbmn7TgU+8KZAy8
V2mdvYzvrHJr79Zo7+wsvPPG7nnuWcnGl52N6Ud+Znah7yfO68FYGfJjMW4ozBBHzBErTguCylqT
jTtFoE6HfHfqtiX6aLPvHzwayzZOuVxu/ONYkhkm7S7dDsP8zERQTKEIQQfFdzy/XqH+ty/6pJKX
y30aFDKY1qg5WwfBYYiMct7HPeK6QSlD2H4iOutROqiDVDWrjNaMYit1iDE8pfWdGFxDk0XAqp3n
N3lQk3eVbJta6nXavRodv3M0VvU0pjREurnfgAsEOd9Wg7kAlNmSyrFoAPPZPXdolTZg+TvouvyQ
+NAQ8P1gIfKpttxCsFUrrpzhvC95nO0JvmwTyMexOCskLyEsA4KQiuUolZE5FbJmibcCt2oe18T5
RqnJ7Ca9zvYHzLc/UhL0FZkR2tYlZVAuZ4SHihNmEmPvrXVOHNFfcpGZSXqVwtzKsoZWWmhL6lLz
iLXS7exUH2LEMUuTsqzj2JAf3HXwi3P0oqGJPp2csAM3GFfvAtsPTCmvU/cspyARZWEYiWi2gwM2
7JkUpuVE84hPOCNe3Z4on9TxYW5pWOsX9HUq8HPvZgAwc0jThqO2//Lhr9R0XzVkyeXx4/i7r40Y
u8bu3MAULHh5WRnqRPeK+ah3LsQiRX4y3753ra4gYv3oLDI371wBdbj5pjzUMLW7Z/AJsNCFXxgo
hysU1BBnzNbICG4iTVzk0GwIvMfO+quiRSpMwn1KP6vPFJDdIYNP2W+Vyla8/hNP6mHe+iBdVkHK
debNHEYA77AVJrBzTAYdVrTL+83CCBAyAd5P5C1drOOo3qBEwlVngdI8c6LxfLjUxlcMMU3xT5/m
5dNCStYJiDqJSTtI5JBEHTPb68EJgJPGZ4DOOt5BWigF1a76wsTsYNX2BjXlAzBedowx5N5nIO5K
pN14KrQi3xH0aAE9ZYRW1QJ5VKOfksBVlBooNNasvua7hKWNQ87bu1XL1QqLN8PphdJeVYo4aSbz
lP4Rui5KJc3tAhWEHvAjlfWsdU4RhufQv2nWC+flEmC3yvueQ2X1gumfQj4o31Pf2XIMFfpOt4fG
6PyH94ulZUaR0xcCL9niYhKCBT4FiElbhBE52fuK0G7ZtBRvYEarXpYI64TjLre2HJMPk1auacJ9
6VdUXccZ51FGeRplDAkAt/feU1YBY2cg/dQw3Fcw33UwhjT18tnF150Fg9Rpr+Q2XhKDKj241SX3
Pnr/siolw6ergCRqKHhB5aj9Q24wx7cxcRUJhkZES2aG1Iit9Ucty65Ha17BwmicVf17tN1b2N/B
Jw0/0ZgfMt5H9TzMlLkYgYG/pJ/fTXMG8Y1zyGRNFUdxn5C0Qwu8VeOOabKF78VCQs1bVyiLDmVk
3Pr3wH4Aln6DigPJW+YhgsjCRScBCpprMflc4KmMYTM/PdLIgN21c90wq1nIKbnyR1LDiXDFJova
LPwrlNZ93E7+DupLuL21sWg3sTHEP/sHqCGaqMZ6LnL9q7zZpwWofgaXNi71F38WltOfhz5BF4HL
kJcXdhuRmGllxHMrAuOzauDnvuDEA58EDynDtLyKaunmtW9Yqr8VQ7tvzlROhMEYVqZX6/Botxai
jD5cTgSGglwgpbnt/CKGSUQXa03Mb6hHhUpK/LBnbZ/Pd+zsbye/IM+OmvKZal2nJGQFBSBIeofo
f2UozZeAzeOgo116tqvjUc+iAwXSXUrBmIemL6X1zT9KCnn7QeKmGUzQeEkgZ6mqOU7AI3Z2pBF9
jCyEiVBl7s9w3b6O67ue3KdLKI5O3msPw3Vz0MdsgZ4glPVGiCMcSE58pq/6eworTLzX6lrWJrsW
T0Ridp4R9GqAEOih5AsOY/NXGabyd5VKsiJgxYqey6fujpsWPWpXZTznqShB7LdMoMKx/zXZkQ7d
J6xG98Yn/osCebafmqP76Kbmmcd+WbVKeZ8tuNWR2eahXyq+1DHGuWE940ayJAwOimu5ru893iVE
pzg/BdZwLO7r4KFMRK0GljUi9CTmRxSLcn7szxXGmm/fGd1rIWcMWu7mSTHDCjvaGuXzJ50eQlPJ
x87xq/D79TprwbKxtlJfOYWyPAbn6uUnsFacJblscXhGRAS9CDwM7U1DALHSEGYqwYs8x3DwdrmE
YeN7m5XSTNJFuSZynn5Azw9odfbEwN2CLS9u+f256jAD1CVE6qIHmF7ox0U4lNZNQp+QwB8xN+PA
i6rMwQpBD11xGt+5i8aBW9VC+51Q1pUcesIalLMn73zVHG4I4mep0e3KaIoKZrLnOrwffp5ToNKQ
9jcDHToiXF78g+t0usGOw731u2z7Vnt4ii+KnCMeIsJ07XYLURQWL624pwxEM0ISgb2p9YJYu2UL
2Gee7jIntlp8k3mz0DPYHSQbR8S/n1o+HG2qN0b/1fXDN4jpfhIiXiqCTckddarIQiJkyrZZp4n/
0sDgzS/e/ujW+9kMbTdW6VBhsAo5ALFlXKxK+4I/+6J/nL2PrA5HobePrOa6V+w4K8NnOz6mL5qe
29jnx9kWPM2cYHURd3OgbmyNPyZH/4zAWfnbTR/RULXIYndn+fzduV5UgwSKHvnVAunhH04yKgHo
oYe3x9IkHJ/DjCyC3pegomw5wR+WYYc3Hs7TZ9dZxvQVbsHDIYZy+GA1mDb74ztBZBfB6nYGwVcy
VtLB89XkX6LOwqJtclz6+bS69fppBfEnZrXPlri8Rc61cxS5PCuwCobG9kfq+hVXMhXiVtySR2nA
0f8HrpzAyQ0Umb+/5RBGAamT0JsPv03DnuXE2/04jUoM4ncipUrRTRKOlLA8+XMpPQs+DUB40LJo
3u86broNoEOIg0bX09fqHP77aojBxQsNXduNpBYycRu0Rq16lQBUVB4s4o4TwDP+kDPSNTic1YR2
iWIIj0fJDVbPfDVFJw2OLEmj/IsSNyRzHB8Kl4UzfR6i6WB7I0BzUqbF3V1Hsec8KP5jOHRIifKY
V8AHhF6AGsIIqLdrhFxE8a4FEid6LhXLcYd3FsgeypeZSypKrQ26EawqHTaU7QmwEAH5+LmQBFvo
8CNjUcrwYOqBoKrVQhRy5r0tOeq/zxO1gPry9N2KKoB3PrrLEOggB0jHcBWja12ileQQcagC3o58
++nkDw1dKU5QFHv1GU9hx0tcFlDMMnC5+03eNTgrXHtgGLk418r02o+Ed/OWndN3iDyxc6xBexAa
q/ENl5CfTUMSgz2I4AJDyIKKQthIwU/3QsAGWGZFl8LgBpSVO4FIrl14QiXzewHHMcdrXYW7SvgN
1afW++h70cHfKEi4rZVhqldj+USsQYm/b77tJ7kSDiN0srEfZm4omkS7xldnJPpV74ODTrsnUK7F
+6xIIyVovLnNn3Fsp95+mV0EntHJYlKnNHOHvwGpBlAuw3IqzrdBHwCyMzLPX10AZP3Dl487b+0U
437gHFIpQy/yb0kt5Fad8S73YTu2Tz0zAzDuVeumntLIxZ6GtysKcCNsePBp5DHqBQ7MH+Cfwffg
IL7v3LzOGN3kknWHkdCsUodQzzHAjnLEEZOxHxM5BRisUJX5LWAMQZyoAHlG2qdipzGF4ovKume7
3e2MWEo/AnKeU+0j8hjxyYiJXj2fERSI0QMdPMCdCnjoie/G4V3mKpcMSmwmJBnFu6D0fbGyVKX7
BTuUGkgtBf1C29Y6wEz+Zj1ErwamwnODomjOGdAHyRekPTmSYNKZdPPLAoFF/Bkwvcp47mXXnGyQ
95F4XTNS+kX0M1nw0jTNAAZT3zhcOf+KwBOMHkKs9BdijhpF+DGw01mIfy3fP7Da+y+EI9TT0ypR
c3XfW5ug0NQKQgDZbCsxzV52jIAf2keiqkwjQwS7PNJtbo+VgTrkB7YpGHV/aBO0ZcBa5OuYAi98
suoraEqQsAYUBE181Q7qLGvxHruhHIt0Hp2aCeXiQtdJ7oLxnuC05lgLOuPkpoWLowua1K6wmq4O
EmKpl8RUFvYil47+7ah4Qq0Zku2r9pJRWEVU08H5Z2A6ejuOxbYebOvpyW1FXlJvAItOH76qrp5R
o8KrClSpN9M+9RJU0tC1HjY8htVvrJQrm21Kw3TGsC/9v/ng0TvTZDbdcprI89p4/QNevuz2pyIw
AeBAUynxD+AGAgrTS+/JlnVt/70r56Pb/FJV0tIfXk31XvKj8jTlwqkYWF4sgRFUL6IhOt4HC0TK
ICEPRV3I7r6ZehqLa38ZwqenbMUbTcU0hXRROPQy7D479LrCvB8pcMcQhHhS2/u9U7/vZCrhNUAJ
rJspflGs1aFWHyxaw7kHvWl+lPKs6+jQfP0GIY4E55WA5DFRgjA06S+x1N0IQJanoPu+UkdKEyXH
d+xu8QEWB2VeMYx99iFR92/rcpBpTAIz5THF0ffCK0DYotuPX75tje+LdpEtrlWCqJfhgvhS2RtT
RVea/UEJZN43+FuJ9bo0H82JBixmEdtFn77Qba+umvTaOpMhv0YO9EWLU5AfHs0UEgrqqQgNP24N
+9UU/3Of7tBUAB1R9s4RyqZPPFJbaC2yzmrjeWewHPKsKNqHOZKbEMrLAnk6fVRjRUtGIhoNMZgR
VpHmEAbbaqu/lQdB5IYGPVcUipxzYeFL7I7GyWlYBT8vu0eHy+rLvvHzQO56801VNua+/NSp16C2
CwLEBCV2ItwgKuXTgAQhlReZ0bzhBveoUtKNUAvCyAKVYS6W1UYpi6KTtvAQtse9alnnIxKWFVAt
XLADSEkSN1BmDZpfuQ9zG378ZQccyd87k+ZqlNLeN4o5mF+fdXJCdCDFHb/u/c6Ss6R3ELiVvdkO
+NqJzNmkfCbe9eQ4obvNQ/mXBTtjalvKPwM+pRt/+G33iduCMZnn6tLvRuiG7jTGlfIxY+euaz99
d2NjWzeRGEAQgkwJs5zna2dQBHEVC27qat0l/ubiMFnoyalfVUi37tZMXSFdTjU4LELicM9DtRK9
PRQ9IDCwsQq9LF/ZWdMWzgWOTxkxiOf/EN2e1xk+BEyq/NomqKnKcT3ktXhslUiMrhbXfXaIwcxf
XFLNCiSCTKzX0XGb0LGoL4gWMScSeaA7BKkaCXcLGsG5hBelhWrirUfbT7S95Ay096ldq9oDgYZJ
jO2pbNYcIVe9A8spa2DYB9uXDHjuzhIP2XD8xRoB5iUgsmWHdJ3uqII8VhEIO3yA1kf2FpFnG/3b
WDjG1YXIYspge/X7dSDRXdFyVJcaPd4mBh3Qa82/zZ/jBAS89hycBg/ki3ia47fcq2y652nkiqNM
7qJ7mMUqXamR5LjiwGDq2WgFA/hnE/y6tjuFtbMuHm6oYqLw9CB/MkR73A5g/vPGF+Hn2Nfyy64D
MZmFoRUcStSEoVgtoMyMh/TLYTkT818r9fv0J328Dvk4QpsMKzppHUjcJiULq3es0W3Sm+TyyQRI
LptAJeEo3nW/CadnjjngEtyU6ZTIN3HEPh09pPh3TEyG2LxO5gVqH74SRybwrAf522ZO1T+qbC2D
Aoo7o9NL12R6x0VrVzhBJ0kG8XkFDp8IHk1DjKI1fv8zmMi5A+H5RVsI96Aq2FuHEDzYgMffLhFC
3ZACEXir0Mn0gO/lorUQS9vOjL5iDbNefv0skih+AzKqXqTLwkK5ny31LwigUwcbMQSKf+nqK2eu
j6eihSCGtJ0g9XhUnWMVl18fdKFOvrcdyArKfc1sXSUZJ6sTbkvVzixR8K14eieM+EYIkd3loNxJ
alK0k8s14mMYhNZ+mw2YlvzZOI8fwkxnGhxS8UhQzeEWf6sh1OnSrpCXQrcrM1x/R5O08hbPsKbp
1gi9rjjXDcNSsFwGGNXgWtcJB2f5WE2GktHc5+6kErXYhc6BxXZe6s9vfbwMPBVwDAyABkVki6aB
Vp+92f7Rms/5IabU5A8CnM0srSS3m0iYFm0NpenZrMqvuER7mTaZQ3LZ0dIVWBbd960OC6EQ4HOt
LRreaK19c/nDYTmL0w2XHY9lvSr0qgHEcqd8M5gdvM7k33oOFa/H8cR+RkqgMep36iBTb/j9gtOP
ZSvnW28EFU635NLVAY983NbWB53e0D8/O/drGIM8aI8aHuYXJDb7Yuxj+QEURaFMmT6QrekNvOjY
mGOP0ShHmMlNHpovtPBGww3VAkQBRwzBhiw4QdA4Speukdn1W558YFkVsh2gl/cX8bdNpK48Qp/B
VX5UJAMEKiPhiRsCB03gC1y9uvWTcJoZcFu/5WCmkE5JZ0mt/OAK2328rhlGAXup89zak8NpGH2V
sl560UyY/vM1zdLoym6kICawcG3tpHbFBIWdzNt8koL/6/yTYNqy6rjub9262X3LgxbUM8uoptkZ
+bkUAIR9y6smb3ZZfd+3HHO7qVUv4f3VTAelrHBfeBOPpODLMTRvUHJMMjTz8S8luMD82sYu9zVh
u/xDVdZuJ/AZDkrI8jetbwEil0f4ZIsqSYsUOp4IDSuncmWTOQFvvXahbSofDfg+iFexJyYvdAMV
sBNRpgiO6xRDCSXL/qKdEi0l0fmCIN6y/FtcU8XBFi5tECPcjCWaDu8ntEpjRa8IzFTJrUzxktsJ
j9k0ydwBaae9PBoY7S6OhgwN17LdGm4UwUYWrfMggGceyEKC23GB3E54oDfcCO3HZy6XPYGNg6Bk
CK8HLJ7G5H8uY8GlkC0s4CDLNNBC82dHHywgJPLANHTct+sR/uQJeWfIcf89D+HUQceoCCQwTbUd
ODAJAbaE0UpDXSm0kbcIZeBFlcTq3q6Q8DrUFauMSZUjCun2tEpS7scQ8YCZvNoW56xQ30Znkx5A
wgPcctXCC3f98ZPvqUGw3zyUIGL8vbTP9kS98sCF1Xmkx5m66P3rEJq2J/AKobqDQQFym2ypp4to
+Yi71UXnkp5HVgBeIIJbhywlHojVYBaNrMWl9De3cMEshb/YWBNr80K8kgeZ/W0ybCMyajcNyMIZ
lWsPm+i9eRuoKHECSVYNDhJ28SJSbZPvtctdXHKXO/WdHXphEjl0D5kcyJPcmNNN8JjLfAeqQUMk
nxyX965CjTCS5mVYjhyRWKiY7p7fv4w125uE9JUl+A1vr3mALAPX0bh8hjuDnjWJSzaAFiDUAOTD
wmVVsVKxPzObabyGM51Qao4Oi7iSTihlQa8UvxqO9X8mSErDx9n9/lkGdFLIBOnqvyzSp+6ZQPsQ
SVvJI0ei8Qp/kCEjLEMb4RPicP9PLD+a7e0Qw7fukVf7bk6FR5EKRMncOxCyKAWUlth1hKZfysrZ
VWO67NHpDalXzixPPwQ+ou3RW+hOc3p+ai4UCkUazW7fF2AgqkZOONJDYnZikczuMN/T5kHk2SeX
E5yDfuOEXHuhdNK6kxd1Uf65f+qOiK/He85hAIH5M/idNQMF7hMdMJPfaHDTn0OIepYCZF9UyrL8
odnNlneX83kDU/nZ4C0bAXhcfMFgu6uS94W/eCP7V/MG/Bq54qT+/nG6OWHzlvB0gYFrlNYFu4RW
i6mViCpAP0APKuMV4WO2k3nea5ZraI3Oa69/DVEDSPf9H/WW54Mcu1gCoKXEPKQFlxU7gU03KitI
hfzrHj0rjki67VdQ7pcfDWJqWmPosfUr5MRYvP4YffKCseYKMj1FCMTHSEwgTVPvdeWDGoMenIni
coy71xk5N+EBE1ozn4JprHvkfDHZQ3yP0RS85dQOX6pN5PogJR2vJc+9/y+HIlcbuWcAPZlFsGpu
ZDMgkXUH+Qu9pGDJnNLDTiEdWkXaio261JVNpxL5pgCD6Org2Srd6iCE4VajfXnUVXlEmwajWjbN
Kgxb4ZsQ3YdqoVlmbQgzekWclLu+OUeeDXI8G/Tia5Soyw3hceO4qG97ypfmanP7bzr9zFDeOmRT
cdjT9LJ1S0sOIdIBRSj8jQmbF3mApIgXcNt7KQE3PXtkKbkb2YXVfj00r5INUdt6ae8ilSua2SOM
B6nLoeDdIU2yonqE9llJGIWsYC0fAkf9WncKQMyHFQuzwMubZFL8ZielnOL9TM/PSJE3HMAeCdT1
WCQ3vVaFcRDT2ps5K9tCHzQhkiL7LxjIIYXOjUCuMJlhlELqS09OsOQllTk/ZregKu3MVWoDmUgW
oKc1fOsRyZcupJQavVQTmVBGWCxRsfWwZ8mcWIZreX/fY2bivCZy1kxghssiZ2x7jMh1ylmcSl6k
h5EwEFDdY4e9XiAGKgYVVuOwGOMw6FN/E7SCyCriNjkf09tMTJe2EFGNutP2EhfyCeSr96YmcKpG
HuB+EEq+a2XrD2cgbQ5B9VblC2PIuPVALngTj8pGd5iDanJj2siDxAnl9DGszHnW/pp994U6Gplk
DcyFY6SsgEVM7OGS3TG0B0wGtlWj5tlCIrh07/hVhvKXG+uBZxIf8xQBp4CvgwmlUz4CZxLQYEKF
94eg/FDutZCMTCi5Wp0crjBoN0XuVAYRNhiymv7kxOAHki6BGC4ywrB+KZ76R0pVNHWnz7mP34AY
AwfCNx1OevYWMrVdzDAi/Jqe+vZKljk7LtZbMYB0d+3rClw/J9xUAvRDxYSVwCXqOGmSKq+f+Ecl
yXppqwBXjveortl/D2y+FVIkm1FiCNaOYs+VlpUBj+GaK3/GvusqWQkV1eu35cUJJhFcnzaBdEOB
9Otle09Oicy8g4QD+ZotoZc2IGGs+8OoeBtxHp4w0VAUIy+haFD5wpLjHPPyMwTv9vQ4VKhlmvjY
6AWALMCqLLcyCFLtg/ZlTQGMAJGM7zpVgQ+1UV8jfS04XEm9alDbbQycIMaVIWvfzXOPvOxhOIlx
qaBZILzRJhe7mLsgeyKut7L+xwzZZ/WocBtziUPqYtXfZREu9tyfBuwtINPVuHMSEmvbMmg5MquV
vnOjSqBe2xxoCxtmLWKVtvbPRrDWqBbB/yMOLRxOPdovuTT3G5j5pDxM7IIAufRtOdP17qOJwR9A
pUQj58snBxA3POK22JQUmiEqnDp+ZPgyGg8/UdFMFlgM8k2sO6ylmKocdxbmlTZ4XJ6SRJ66v/L0
n9/Yn8h4q61Xjx2l15SQX+nvGaqYBxi6TfjKoE4YeQuPItmtcqeRl7UkEVl0ZivB+qlOvV9L4/sp
QKRf57RDWxe08lEsD2DTzGniuCkz1TAnF3UKJAY3v0zqPdYzSSmBQENvYpRdnhpxWyvtcPlXdYCa
uFP1RpfP1oH/ik9tMMrdi7utUwnUA2VGFNoDnw73zJy+0vnTB8t/LWX+tG2/sJOcWsbuH+SKMpe0
Fo14GCTjCWmM6OWhaurpoYw7Gwe9xKb7hxks9Ci5VhrAihSJFrX9hGWKMZ+pIbHTYSdqPYfsI6e9
HwwjBDpMfDnclJM60lpLCl62yGpBvWI/bDIGfsfxYeDiKdnLsck/osM4SkPD3YISJrbv42VIYyoz
WcgB4BA1bdEuu82KhPAk87hYSH+7MAkya5c+XmM6TQnADF9k7zaTQlBPUsvvfi9T9u8Sum42pLrX
kVWn+Fnm6vOvvn8W1k/5O4wj9vbv2AjgfzbWubGa18c8eLjOCFDQMhd2DI9Hm8LF8hGvgiLioDxX
l8gGNLHwV0ZgvDvCJfWx7MezP/6vc6Owdh9qktGnlWilwj/9nlN362V0ChcoOJuuTFSb6egf6TU8
zMuHfDwPY5lFL2IK+G52mMStDzPs0LDNmWxEulyzHyMLeoMs4r0kZ/kNE9BkLCkHd3Vb+Edg1aiw
DZ02sXxY/TrjfosL0NPlJK9TcFGuj1xpIRFYq5mgvz1AeztvpjtkmsyTR3Uag1ErfClmkt+Xci+U
usAlgvDgLqbtH9uT7qK3zWZpkPFOLH1nSfS0nSgXwCl1l8H7ZbleR6Sfk11LcR2/6FkUcYVDn2Nl
+6ZPsrMB8CFQrFJWZCBOK7qnTB+JjlA8UlIpH2K4LRAkbtpsUNNcphfv+fCDlNj3A7BQAIHpmFPW
owtxU/8UKyjxcwy1EVyyP2PuyVhr49teq5gc6aU8fXRS0Goc/+fHQsarCQPMedSSNBywd+rwMdS9
OFQ1iWgR+hdtplJ+Pxm4XXTqLGf4wGrQVIi62p75RaZZUBy2k3UmwfLwG86JviPnv8E/P2/YZkDX
69aJVe6l7XKPWdGlNRttXhAjSAFFGOUzRuNQjw4piSubWBfhAGGh/7aKu9Yq9O24wenDBYWrCSmD
lpWv2L+DiynyUJXgjuQ/rvqrlG9CV8Cn1Q81Yx+S1TOFU2UF7L5ieCbJXx7ha5y2SWMiKMvxxyyf
jg/XHAgygSrIP0knbpE2q6g6whbIMYIPuuGb/W49jlmi5+RbWeVCH5qWyJL62AB3j6MmJnrv6jd+
lTGgNKSVmAsjwhLk+a9mXWIJgTEVx8DDW2ffETd3aKkueK1B3RtXKIqdYcrssEsm/+0c1mK16PIc
w5Zkg9KORYSfpwwJRWfBEeqQ2vgMCFm7UVYTnwX/2BXgeR+9h/ptzjaSbpZtrZWSONrAfER9i6BA
stdwdWlNN2nQC+q3Aa1ZEKeoe67KFgJQq59XHdcpCzkzTH+WSG5I8JyUcMEzD+IJBOyVLaHITIkU
piBDFs0aa8sYgH6e9iZmqD/vb6d9MQ0VO1mGfXw7QMQ3O0ZesNagy4MFqOUinxa5Zsppj4IeXoTp
dTuQ9G9JTB960CnNR+aqWm2/qJkWnSYO20o4X/QMfG+FQW7ALYnvNY+Oe3Amn25uKaS0YAvVig5i
9A+gM+aEYxdrj4YtQ2wmTi4++er0MmOMhP4QK1P/PlAWwnw7wLqHDF3JvBpS6O9xDxGqLu+hs3c4
Jf4p7geJELAe1xGsOZ5vuyNRrwUh57FqiItvzgrmtzl9vSMWpnpmNJirX3lKWN2GzffYjevAe67j
VbYmkfQTPIFgQlolMMXVejTPk3ELeWO36Vy30cw5jhZ+WBC7x0UMlRFSo+3/ZM0W2ND+ISDsjOd2
/QkQeEwxQy9tu9k59tTw+bxK7JH/C5mPqg1rTOTJgU3mlHP5XTXdYoGRNZjtttBCRZeACLZ0Z5X2
+Y8xHF1ptwfhG87LjV39m1AkInU8AxmGkIRXYn8VhR9cYFatzvIEnt322V0yxmqhoqfC8ZgYe+JE
pgOIg5BAjlUcfxy0DNb35XAXWzyKCfOnRRVqbtPZwzRfT4ilX+nrUBZKITJWDZxeQUckhDY3og1o
f6y6hTdvT6x845hcWNHh7KxUze5USPUR72LbKZMoSi7QG4httMlos6PtSo18WvrHXyzZUbfjzCOz
hKBU9ocrkIu4VE642PPgMC0Sln+Dt/9gYe1BUl4HWc4rbrpHE0/AAeZT9khKOphoTghSs4XoQiCI
BcAGONpR0dJV3uXRbddm4gNE3yhBaCzLTS0iSvYSm4XeqBjfPgRsbKuUe4otWgAN4ok5jNKIbXHz
MqfVDO2DLnZq7s37AXpX2+Q5CD6/DGTYOmKWw/mTHlQh/O8sSc1yxD954zn+bvADjJYCw6L1pPEk
/EfJ7AhQLzMxJohttqSLWNifKifAvaG+UGSGfE3nyFE3UYM7ZdgC9PbjujHb1458FRB7PxlxY8iK
perWg3UJZTd3PFmQxbXiXzgIAtPW0bgxXUokGAmyxjXfac0sWiWwLsWwXCpHrSR9+DsOUZa5ua7O
l6aqrklCDQE74oDkWYoX4bpXCSowlecukug63Vpk22E1+KnhlJxPct5u069YCkls92YNjJxhZ5u3
MvPfrNcocstTau07Naao7+YbxsuXRHXiQJ5PzL+BxkeGixpfOWZZgJrszyY4W0IarammcAEkEzzj
1IRzLQAvSeUYXbcrJMiXI91uyqE2oBWwOaEDt2j3Uq72Dv8jYpbvFay9IDbVa21qaCr2ONJVzWuZ
7rOw3eDoSTsOP7Cmf+ZprHPmb29697R2EvQ7Hkgb7TMCLpkES+2ovHc0T0/0Ro/absfM/MExuyX4
Sp1QxwwwxbaN0gGVyZOo46HQIRldmBsZKuiJRrRXM6wwhgdtpgYt4H0r4COzCavPOzOddd4WeTFq
liKKSgPMq7+8LZPEHhCcmv1WK2+Nf2Z20XvPKIfaskdtuSap5fVQ3B4mQT8695rkasCN1TBVSU4G
3trCUNeUTEOBaHryF7kVf9oGFI7/QypiKR+vj4P18CTdEk4R2ucNPFv/btqYeI64S47NXmQzzqPL
XTJfOlhscyQQQ26S3ytpITnjH+W9iJnxCVPPM7SwNujonXhIsNjJmAkfaTkRHzKOcHZw5/iPJbiv
3vYZhA1XahtHFsV/TXsL73LD01K10G76RK99L20B0fDf4+TodyxIJb6zcsip17cya0mEx+RJg51l
epah5X2vWFzsUyAwm9ICO+Q4Im8vePcGHJdlN3qvCb18+IQUqNmQFMQKmuz+p8yo3skkR3YxSqfl
p/5dcYCrgv55sk6sSnOMG+esOzboADBgaBP9GmvW2MD/ieCKtps312o1BHKXogNtVcnPT57TfE8Q
edOhQcBCugy3VDmJ/VxcSfBxjUF+FrlVd3zv+EQ/eQUmoAvTbC1N5/PZ46H0SQ6rPDKHEKE0X8Aq
AjksA0GWmgZMsUPxDt824msTDOjR0dgflMubFss+YkCX5UKfNXjIfgGejEt+yW5yifbmNnBp4Y8A
N7QF3uHIKsENb8QKMbsRW24mBrbfpjTlSOfkKSTCM3syYkdZFMvZ61+4p3bhDN6Cpbh0TMJOZCIM
5qf7l2jv+vMLXdLi3xpE87ug+pW4dqj6VUVb57ZfeS4uMcU4OUObzZVnDUMtzInCtfmuG2aJCQtZ
IeRhzFuYJ5023HOV8qRZK335ft7zV6gbGEAnnv0dW4nZdlTpAe/quHLd9ENolebz5v93/8aMq9y+
xe52tfaozNvvXniNhEKzUsJ11MjFnmZ3A2C/YdoiLOh1QG5Y3y7xB7/o6HX07naqWu5smy3N55Bd
6HuLaM+MBumyMhJ4gDQRAAaqZJ2hJr3O3jNMmE3QvX9sBKwGFwGOEyLcFbUntdATzL/99pwy+Dcx
bWvys69Q7ZwLPh1re/LEBEYmr+EB35RCjVf/gzPhfJlLT697Mx4uGvy1yFdps48v0zSL/Mh5mkli
ucBXEuo/yT5v6+VY8PvmYL2IXyz7+QAD97SFngSMPgf3V2S4MFP2u0yIDNCt+ax30eJceGUbFsTq
ZFT/aNpMzz6ysUb4Rb4a01AIB/Ahi40YjzoUbfCoP3GjLYPmeYAIi+ifV7r7r/Tji2rELxk8LgNz
PkVzEIxq4nhDvjvhuFW2d3if7/jZRLeNEFcNK9hKbaV+l+XJ++OI3XFhoTjKizL8glekAu2vrcRI
Xgv7+tQpmxCk5AqSGk/B1IJFK7Qv4deyVIp0sr4rK3tJT5XQnwNpHMUIGJguNqTUPqwljNmZxV+6
G73b6uZSP5lqz1aT1LWPUxIyhmf/VewlCmKvWOuZGR8ZmifrSK6MJ8WlnM3ut8nk/eIOBjMEf9Ff
ZBXXp9iKdZ4190zEtydoauRkuLLeU7hQwtBAYn4G4g6qzPPmuLsEbMQ7rOH2b1L9wKOa/el2BPBj
xC6X9XSbWjfcNuhAVfan6HhraLSZX6vpVXXhalxwhQMSW3ki2yRsA11scxgTfWX2QcbaKIhypo2f
IQutI2FNvl80tU7Fg9g6/XfAVMbS2LmJbvF7jfSo5e6Ya+rgMWsNcQaXzD6ATRvVedsd7kJt++Aw
63+AD3RBcsDLByaJShL1khc7Rg7cyNmNvoC6ABQqYgXPwiEpX/2SujlzLl+bHwLNsUUiQK7xsybY
3/i1PwQZUzFJZCM4Hwzul+kYqXybuD99hLVmSQglYG9Rxuo71BJV/KPhaE96nMzxVnjJG+fEGgLM
buPgV1R3pIY+ECmOnWI7aLChtV5bi0UGlXbrX+N9z9kwYKz3MNG0RL81jIylz6tvW1XPO8tSOhi0
nun+9bhqsBHsbVzr2mB4J/pl5ZM/lZRrWqrcSYOJdp00yg713SJYIIjPv4wuKx05D/zSkR+0iQCc
pmPmIypYQrTjLGRZFyt2oEYhO/tQl0I/t38T81Bga97Nf40RmXiHwM4SnTiVIfovy9HJB7XigeCI
TZjfj4e0v2avdRuZqnzQiayRpXHVnFO0bnZ75DiX9QHJl1mBYUMrlX9ToxNb7gs7X3MgEHB/o3o4
rVYm4kix8WJ2w/1zxrr9mgUXFYkcfLaSG24WexjYXm0+JmEfXj2yyb2WXxYNaGzjbLYHejXvawK3
0CscPN7VCc9BTfWMM0HyMHz7oGMVAdF/RD1yJ7CUN47FZBOcPCTA0fNM1Z/76YYG06X4nDV20bzl
Rz1ZAnFX8gteTH+z3LOnfgI44okiti+A5XB0ongg0TKESpm2bGYuxn+mMz0huxb6Yxk+9KodtxfB
GGyhT0tK+gVVSZB21E/UQRkK3Tsm8V0Q8Irc34fQth3RyLnz+KtOSY0FN6+FtmJZuPQCQCQL18D0
xvJ9FZZSMFUSeLOpY8rBCzUko8TVTGdNyLIoZqkP3XHEx7PhlOvY6WsuhIM0gzdlR0kbn3tdFKaY
ZmjejKw7/p1QqUmspghW5oUY7tykS1rL6Ugkso0wkgbLDs4WTRD8ZGjC6YaHUixrG7VL/PS5aF3H
EMeHiLLceqFTPF4Ty9g0I+peVNvtC6cMoyRkV0af5BFc26p+NyZPtcKjNLKv3bzTxepLayk1ODBN
AkjRjhc6SzkiksRZOqh54J8hNOyUF/kYL/0C7xVGT+GioDCEfsPLkTG4fYz4HK/ZxShVki60lK/3
IpQFfsnuqUFiPNhuQKS+Rx7OGqBnRjUq1LWWH5aQsPyqsEifNcqSlEq96P0MtX0vV/zI1P0VN7lb
996V2ql2n87atZcITJAB63bZx6vmPwVeXjseBmjXhFzDtH902f8MZeqDHqFIcdX5drBBvVnhveQs
5XD7ZiOhJj3UwhA9dD7ZgExCUxxC+WAaKUDhMlz8+iOJl/FTUKXD3Jz+qYj1fh/urnZy5zUcDORQ
ddUlZ0zd+9W80t4+2oDhnbgFDzlqqvsFVLbwU70w6SqDSUb3mTvOUTmlBGOFnBZElkeoguTnkQHW
IaJspqHQzKI/0qAZPws9+y9TseazQOBooAVOLcFT9LTX94ZqSKT7oKxgdWaAPS1n+a5n+H+aayek
BvfG/bhOZjAVp6K+fLRZR+lD0+XmyeMGkoI+QfXqVGpMxQAozNU1UeaxqTO9LViMZMhqbhlELo/N
S7QN5dfsnbKVO1tMI55T6kjwEps5znMQjo+8j2ufM9dF38mAJt3mtXtTTdBwvw/d7rt6oSOGvJQr
0GgKmTkAg31C3Wp0u+fYh8FG591XP0MlwVddAVb5PMByDC/avkQKEhrXi2aiX6yo4x3guTt5VYjA
ww4n0eUSkeGCpOriCsAaMGdj9aCvp0eMFRJ2o2jJBwf4mmnkn36q1wZcwYzvYajCmIefHo6NllOp
S2QoPasCdoqX9QAvrsGo/8d9sixs8s0Xy5BVexli2jHkvvJZpZS9JnpfX8po0JavG23dBM4Xl+Pz
9R2x8GpR7TDsVdBXwgSSjqAGVFdssQdM83IYrRY1qTiLuoACdZkt0cpKJ0T1M3vp+HDF1+XA3lRE
LI2OwE81y2XQIGZlU4Rno3FcA8TdnZxCWuK38lwFH400v3+upQ/1N3zi7PwJWc7Z7Ggb1f62jTra
aMCTy8bhoJ3IHAoed3rMIILA2xrwxOc4Ku0k+qfw7vfcuXYlWfd8d+6K3KiN3g6vhSz4Je81x0a9
V3HAr3WMVcWMklkaROY8a2FOlihCEugQD8QxZnx3YaH1gyXwGAGuA1bnbq09IMiRcpQ3DRAWV4Ab
g1Y6Gqcc8MlveCWeMD4wQk1vnC8ByUVg3nW0Q6faH4ONvEOCyow3VWNW/SQY//KDBwnXWXSBvw0p
etgOalOcn1aJbqBhbASKk5TBniSAgVKs4TGOKadTu8rwMYJVnFW+6xfkrZ7r/Vtn3Uc7p+Qs4VdQ
jWF26GTJJ8zaAXEs71Wji0kFnKumscbxLEdFgFHgmLR1RaqdyK2gYjpJ31jD0Q6U2aSYLw1zsMQw
L0h8yCTF8EUO3m2E93XMPwm9MO4jL0WOLbZHvAwOBL6fT8Zge3vaiTco3l8QGaZPl4woHf0v+vOi
HQGMyh66fCSjDqb/Jsz/JXfT3CNhNOVxlEqfTpzc+7dYEhYFXDGBxJyvMYShNP1XZW6Ym1tbNOQL
Hfaqss7cbXWGXyhE3eAz1Qt0Z1hzV0VV0/MYIZ673FIgMDvTD/SeddmHQzhhmA5ZQgYa2hJvKQOg
WCDKmljPboUxPxoXZzuLYEt4gkmzp64wUHfUZaYAOIW0G0gCnZYBfUBQZGZJQcuy6AWfo1DPbVMo
MIt0QWxg2XucNZbJ5sXnVhDNj0iDwimZk+z0CdppS9e2juU/nG0BqIWrgKl62RgPLrBk7ZveMvtl
4UQ58MlqgWHojd3bsi38Ef2CPprdGo3FwtdfA/BQBygizI9oMBFFhCYcQL3ZBfqwC7226NWtyjez
Yhks8BF4Q+Ng35BlRoqmQmPreOCerk3IHP5FO9GPMytstqdpCaEnCQB7Pi4uD03gDYiK/ORAV5Hs
HS6lju0mzMPMIJrMQ/hgYztajmAZFggM/BSreU+i7xg9E13J91Mj5sNJQfarZ6dpyIs/5YyqOYqX
kQu66tdtsY0DE8XtPaypyaUfYJt+MBe2+jzDFNETEz6WqH6IxoPIZVCEtvwG7gcxwLERDX03bfhI
NONpxlersUFzFG8HOJdnAGmLMj6XYoi4uKFfV3cal5AVDzJKQ1HbErHe20/VJzgYLi0WzUtxQpw2
lKHhKDGuCWe5utfbGEbboPN/gKnV04DHZJ3e8PIJTvw6RnSngyZes1cWuoV55leoFZngD/4NfoXu
cmJW2qu/dmGJRTEVDkkOErUyoXpC3JY9UABFpuCS8+LCa+KqgP+hdeuuz4Uek9dBREnisA38ir31
oiwALiPDaV2GxpEbj++oWpykPmwC1fqyEG8jyW042eZQRUfqghSEVg6cXFkqCX6kHiWGyjEklcVN
t23blQ4fPBXdUssEfwsrBJCV31xANFPlURyCzshLG9JY3/UKH1oN5eXouDvur3/FHa8W+aKqUZqD
mKQRuv+fJ2FleFwvCcbUsbnXNC0pK5vJjwmK0MxZQWI3mtHECNoO/sZksm6vGLremAU9Tq4mIGPD
4Ee8TV+0/yF0WV5hqUxm2LuBXwfMJjkqQOVsKn3mzwJs440LODTLwnlZVtfUsvBX+wCOYMw10Kf6
e+1CmwmPanaoHFjLyf5rKO7ByaQspY2K+6ouQ7yyWvMpwHrBs+e5hfDSQ6oViUMtixV9X/Rz91AM
8sv0GFe/LkX5qWLMO22ZsiBZ9c868aT+4henV5y4GDl7bP+sfUoqGK/K/CPawv66+4ez/mLA19cD
kGcC1MJ+zCfkVBG1icmbuBMrIuqY0mxe9uUbUip4k+Q9vP56ZgrVFyjhapVxSU5DNyV9PuUL3YnD
ObFxln8kH6moYKmpRU0zb8C4tJ5tyhfbN+OCUoM5FlhgMYoYRNWPSRCp2FB1KQ9JKT8HMlARebyD
Wzhdw4wNBJvqd8YvsC39MsWSltQ/UV0hwQo4L9mn1NzzfOotsc/mWkZHlC6nhqH2MnAbTTVdJOgc
AwhqOfrRucSOxPmHIExuty+DvjZb2sxESZkGxVvt0H77d7SxJpY9uT/72V9UO3Bp0UNDZfdw+NA3
JFn11snBPYyOxYx3+Hu0Yo5HF8QbZe8MZHgD7RcWDgayLoDphuzTa7ob/pG5z88PG8fkcR575Rro
rexDbFhQzUqukfdVB9GbVSBj3mkziiX8LTQ5vJmANqARRHKLWifVZFyn4mMi4bXOiWnSnCejx1Rz
AYT/WnFfDTDeqg/a+sjBfijNOQXIFjU9wCMKz5vQN9FmZcBNxEEihJGEoP9KFIItZMUgQmBcViaa
LhdgxGJQJ6h7r07jmlTb7pWY9KNAbWywdWAZOr869551BkztC5wNFjJcB3IVJdEExmXgwrBvtdkR
OGwbooVxgnVBmuGemsQQj8HVJ6PIdU7ZPfbjkjLoPEYsVkSUw6B/r+X10VhJ06ueeYThb264szL0
L6+Rp/wHE/yqloI8tLA+wlzaqDbVbh59XDMdTXMgBTly/+rSC+Ghhmjshaq5QiQpWlpBoocST3lJ
MTRq5KuiFs4D2350iKCQ4EL78tYuUxzhyy/GiW7NXMwhcdoFO3hKGuWkKAfd3SQ8OrV+paeq6Cvy
qhoxQO0cvCnfQ9agmtr/Np5FL8ZJGgmOI6MoyDBS8se8ewdSIoPZNyHn1rAfQvOUsKGHLFyYY81G
q+xVycnqYYOvk5ZDwAj6hUuyylILDOzRIRhE6MZSIu4KPjYMhbvemJ0cMVwqYadMgfGPiHtfjHCM
wcd0nwkSC9bII22LZP+tYoA1Hi9c8A6Im3UBAIr7MYWTtEHVgVJxK3FVc1eEVlqL3twrSpkjQDCQ
wF0lPvFNa2/jQZAXlTKGq8QMDzHV4B57OUolxkcy8XyO6EeTzv4Gy1mc8ChcBaCjUEi/9Yf3yhIf
2jc3dQ9XU3gSfoFN3wBicQjv8W+1XByJUp2J3QxFqiveYDmhV49aDGXZbXgS4ZmiA559fW0K3xjY
gyRdbY7xAYsO7RKzs5HfPb5qxuU5UMcdf+Or89MYhECCuf3CJCdeR613Cgh3bIWxibGVTPLlU/ZZ
kwdtUCsS8Gth2QYTnQtnV1fFo8M3zjOf0n3l1Eo6A2SBaXLsZi1YQlGZj4cF4jqYQ+ZYC8ENv9+N
gyteY7IL7NlBgEHZvtkNUK3ZUOjcjGXrqPh4s7vO/9eLV5NaXdd2nGVMV9nqpfohr2cnBqjHUbzF
v6pbhaGvDQ46O3BWEdptvtBav/XQW9tjJTjPzvSntaqcRSlOAX/O8eZka9hjsRl58PSlzRWV0jHl
aAp+ZNdEaEdaDGqBHYN8m2e6X0oQbse6wGPsGVWAiItOMSm4YM9qaUAGgZmIxfBC/LxVEC1fxUj2
t5pkewjLWFoI9+ue1qBxZelYHAHUVskBkqwCiuCU8KN3Ycwr0xKOY+UT9ogpeU0QFfZxy15XRr0A
M+i+WloKRwZ//J6VSKV2ZY/kap89YjOiPhVxhkJEw8icMlhur7rQ+K0yIqy8JIbWBMwCLP0KTXp/
yRlsUvn2ytaGcMAhQRJ8Cekeo8yOGIrIm19Pi0lK9jljkUtaqcE3qO0VopZmDx9oV6jKrK2v0/aG
nU25EjbISoSOseYG9DIRRgco2HxFqHBg7PCM0o0EnlYNgIke455NqSNHmubqrd8cotjo7RF7teqA
OWHncMCpQgS/HXDI/VqSPkrt99GQibo6aROFAuOj8W+kKsqIkZX1COapwiwOERz8caY7DqEApuDz
bt8XPvs8j8If48oPCRLVvsFC+4l3Fez/WPlktYtHH78V/tkxDaYB/HRpTvIATNi0ApbGTj5lvygK
hmwluOdRoEHt1C2cQcl/8XBHMvi3TcWZtuQQkk7DpUijMQtnOQZXrX4s82El0KEbpTxzAw5eNHRb
j6O/0+7FftYffqkK1nR7v2aSHISZZ65jJo6fRpI+ALQoUnrjc08Vc1DIHAjuhEAx8IxD5L8NJ1Ye
WdYVAx+BFkwBaJRGX9d2l6AAJv7zqnyXawG0ukuzrNogUHNjArgqG8D7yMz1VEU63BA0Vsj44HKR
0aHC/uBfy8jH0n9FpccOuWPtI5sYNLm+K+EgZeDmqangQTkvM0hHB0Ep+2mLyIgcfttZeaKttnqf
cDCj7UL6ZQtttx65znMk8gYKTrYKIR+4ywVzBey4O09BVzsIaysbZscfXKf9JxJCctdjfNTqoVik
8EgWgL2ID+CL4+Xh/KCJVvjjuWVWeZAMDkYBf5RKy0rcApEn58gMyreh94RgPQofvbxZfRntJzT/
THynwkXdjpGhJYrp8oJwBlgzq3O5GFKF895AQY9Qr0eIO+d32VhK/KidSb9stdp/ju0GJs9GguIj
oyTb/aM2Lm1zmIEmzbyt+JIt6/0r4O8rzFbCMtWxnC5KyT67SgWuNj2aTGexH2ynPHc7PXa0PUYv
Pb3L1yPPD7X99awyUajw4yQzXT83ui4uktfZs8l0zgBrjgRq7+iHKbGAcUdNzOH5SYHH+/stmfUU
HAZLl6mkl7v5VJdpAaKNCemUr1yxtGbeOcZRDbEne+fI5xoZECyMHRw84+wvrcUS2oYTO1uzBDmb
FQyo3qdoe1XXEPgz0iCJO5mVIs4PMEhFolqI6ZMxzhDAP1Iga77dNf+6VcEcFR1iAUprDQUo7wtg
mXrK26sf0ksh5eAN2Rx7SH2vKIc/ELaHbq1MSi14LjWjAXveVBmccr38vMHzqn1iyEF+KTNSTgUc
AXdHnGo71G4gU7LpIAbMWWAguuRj/fsR/0iiMq4x6oj4O9jKky1RdsafF3OQhhTN2xFfec/y+fop
qcD8OMChw8TU1QtZTn9lCH+NMyp5+Cm1C/3DIYdpjaTUtjzuwdPP3a/t+gWBmtNGvpv99rz0i7+S
gaPMsevJ5vCrfRbBXIWgH7EgQd5jMwW/fIP2eAwzSaplYb323DWQwpEXmrs+OQl+gHrJpj7cIyDY
kS2xbv0EOF+IReTuCUIYVmqXdutLw/xAcRtd7+2vU96V2+CBhFAC4JHGMycETKE2hd7qoEck0yOT
JaAniuGnbwzitnnfRdmd331dfUhvmoIvb7Lt1JRb2hAZKN7EZsvzXEhr3kNf1AtG7fK/kKRVVNNI
rgW8MgSzOlOVv7ytSJRh8hW2Jg9DsItZGghHzqE5+s18ElgNbebv8cQSxXSRHuGUmw3l3akIJq2H
HDekpbLV8SFw8+fBdLneEyDbDtJZjRRtkQC4BU3YVbxgk+AZmJEoCNYnzKwf+5qeMMpmyOiWnfzJ
lnjZzgDehIuwMKHR0ZVW0U9ekpNJFvkll4OJr0UEWF570lVowsxepDSh6RzkFrRVAWaH9WjtNFQQ
e3AaMqrwzLptLi/BNxde7MXPyAuwut7olU3U58T6ms960NReEcXbp5Zcg6tNPFynVdlkCFOnHlEi
7PxQ5lG+49T68PKV+NGBqZzD3p3XKsUabBjbD6aD6qNqmTuRYaKww6brwdcBsbUEs3JlAfUq/YF3
yin7GB7YfcbfZ4KVII4aP7BxduQnWB1nOPNbeOv4HBFnBiMdZkNb3Ffk8fB8fzSQkuDqX2ae6VO7
vHovmJJFQoNDCxc0y9lalTSYpBPghQk+9D8hOj4l4Hmab0thTEuwpv2DM9kGCU+U0pb92K8nhrzO
+jZCiAABE1P8Ta+/5Fxzrb0irn4t104cU4aHfRNFTQvj9rsaztjtlMWTCNIwjn7oOWJnjzoMbuC6
noixnO8RPiL9wL78sA3cIzQbm9lAt5B27GLp6FL+UqucRSCWFNsxJm8eyb9Z/SAF2mDavbQHbqq1
CfpTn4XD8YQw7FbA4KFQ9TndEbFuEZUwJd6P9IxxP0wYKSQ3EV+PnGvw2A9P6wcDemx/LtNSMcvH
+4Jue/luAYco4a3RpiUCgP/I4mg9mDvLik9n6XU6dJbbR9mnYQJEVR+uX0Fec5ivniBkTnBCJ058
xpJPEPmgBJNFx539yfrwsKsnBMX4tCkGBlM4bDZWvJjZ7gso+u2S0I4Eku6n1KWC13yLsmtWVqTc
M8kvEZRLzhVSbloL1vYPr1NNEL3bqTlpg0ATe2LKggjHuYcuiqq7pVby9/Foib7A1MXiHvHSsQlT
Kme2la4RAW7PCV5GP/ExSeFPFid8VdkPw0LXt4oHvbDj5BtSpTxS7vMKE0OKcNMVHxcXN5QQmggI
/2sIICfKrlKjGLZRju4C5fZEmgoyd5JysZ7KK4qUG5Y3OW+6KPTOhUsHjQcPRb9PttdJW6HFhvVD
cEr90Ef6O9N/Es/TVMUN/qZBuXdSOA0TYTnAti0LVFREftMGL+B43uqJ103A+zXXlFfFdgMr7yYB
StUS0EXhecD2UZQIv78mkfoRC3AVsr75cPmYQ3D4fN/jrGTppgZCSNZjEVv6ygF9Xf8ZOMTl7ctW
gqnTzpbHX1Z6aNWVV2gbO0qWNutlD7Szv/XqqHnpJ1WtUHyZj8D/xa/zVPj8YswmogogkmYp6NMb
Pic2vBZQ8ym/WQFEONZASOmYpXy/V98VjXVkoC37np7ji+bZssvsyAwm5pVqM86rTCUqb+87RODN
U+BIjRWv0CY/ZjtAmTlQh4NpkdhLfMgtfWfUB44VHcZzwRLnERKelTm9GacC7xSY6SzGrYGwgDYB
pxWhY44QC761xiApbOJC6YfQKT3OwL7w3/y5qJygE4DL/9xIWM0tbK5BtQ376cSMW8JJQboLLxEO
jSkE9cAkKFBgI/L1fiajtAhlF+C3JN1KRPRa4nqQlgq/GAqqSzThK2iN5INvFl0LuOr64f6jBkuD
rc2cD/hoJl9ZUA7NC+k2NE5HbnxSLE6VZ2gRIRaSX2Ub7ffLoOJEWWA/0VIRsJ0f++vUPTLdI6F7
m+loh5XOrK0rRCGBBDxG1ZiKdEG4aG/FSy8Y8xkFzRZ1+iLifij4dEOkVcGUpTjLkko94VSrNvp2
NDqTrcGdxj3U9+82onNUfwHmDo9ewC/paOmx2Nh1tr42lGHBs6fzYeLMyt/mWGChD7cKl3fHg74a
ct3CVZtcFbxHGSYiPPaOMwowZO9dpWhw0KOTbhxrY8+ibPOLAo0Z4h+uhJBVbYFh+N0q2x5mtIWE
zafhdUbu12RfFlViRxVCT1PFc2j0CS9yPMgvtM1GysCm31eOAd5TZ9rr7vzEm1vo11fgmEB18/dD
WV+ao7MjDIxFyr40jUzQ/gjSgv3r8Z+Bjs5IEyFOZceSC+pjenI1qrYIK0Re9abuzbABzB6FFYk+
gGdkNetPWE4CDwgjwnF2zJGpMVrBKVyZQsJNwfuvhQ/XV15hBvDO3sjX0yOnDnawqbWRFbh0A9+f
Xzkwa600AQ1llhUJaN53zmNDCY+Z0NYryLQnpR9lvz5NbEjeeeW4S+J+vjf3oz036wmkVHTV5pS1
/Ssw4Fx1sNsaBmL5wPNh3wGx/U16Kdc2V4W/1p45ja5l8KfVOTzKfL+SMJSxGYqpHmUzCm9UNTNo
prz9V2b2KTKl/ArlN1KgXqhpR/zVrQPkUZUQHFF7OqzNyqJZqAOAU2xUcCpt61ZWl0eAehUQpvK+
Dxl2ZCOaxhYId2YH3EaB/nWNLw0ouwUU76RZrpiW0c60YUfwB2jjNTQYK5TT0RE2Hcn1B5tzrmUy
Z3ucoNrGioYDqLHCSF94pyfvmNo2ztKdHdfIVbX7BQQWuDa4va4ATz7b06M91Y1VdxZrI0jp1cnc
tfm37DqrIBFJQqzvLHSYsOoFl+60ShLMpJ+48L2+ZVNiEoR5pbw3ELBjXmA1VuNsglKAafgTvUSF
i/YRPxV9GQurdWHyp6HnxhAQ4SxPdckrbpZd87Uei+zcw+ILczCl41VyNYAlttQABv/HIDb10pgy
UWwan4qwNyvMB/CkCAO8g6bd+TS4hTs7xyT71yzEx+52MBrzqhBtXJ4imp8O4Jh93CvUVtjqPrxE
A5ke/ily8mRxYs+k7q4G0oQ7syE5LxJ526QrxyGsMSlvltf/zp+v5gpx13/sdWnTgKVGqMqLHu5q
xsY6A7X/5P3DDpdUjO7ZSUuS6sVIViLZfeCdDVBthcW+V+cRuT/MPM2jVDbYXZ8A4KOpXSUzkJgD
8FSg+bgAaeTb4F2EjPRrZjqY1cBqn+GHdmovX2zDI0smgWQSseT7IgRMTEafDdb7sXLWNKojK0ja
eroAVWxsM4MeCfX3ZlRbksxGgsyiLjVjKLzurRgP6lYWo38B1kRvdj8aD+D6cvLzevVxfF4Ozn+j
YF6MMMgFRMZVnQI2XR3ntDOPQ0CFhH2w+J6rj1qR3RoB3mKTdsPCLGBL0hR1RDD22JPjCYSgaZ93
9XJUl4+lDerfiWyp5nj+drYXNxWBgqbqidLRA17nh/IIpojMghMZHp152xoJBZ28X9RA/o8GOfHp
F5nlrlD8xmMuk+SFT0mkfdw87NnBMVvWt8ztdjRhytuiCQdbheVh4Dnbo7XPP9+YqfwMKfawN6L5
3neHiVMTC5q/ephxwf+8MZRfAYHl8vQkAHtlUjsaFD3DWHi/TjXxodejRObDumAF/RcIku/NdXeD
Wv1z+BvX/lzgO2xQkieXL+0qthai5yV4UfKcEGBoBNfmkKQOOrqf5SvzqtDMW2mfCCoaf5m9mGnm
/4u9Rjo3yVgDazpJ7CMXdb1+SQuTpxAaseEu1+sLMWqI46xqNi6H2nmEJ7Am5KbC/IlrFotDdQHz
fzKCopivXcxWRQsp+yFPBmxTBwABb8U4goJmTAEMOe40Jsk1Lcz1w4ono5Gahp+lxtxIACeqdSCg
sJOHUaXcdfN9wVAaCHd5WKgpw5fQuZ9oJsMiGAX2YY/0c3ws6O8Yk8KCwLsFO0rX5Ip8PgAtQNDO
KI7xzPY4CpQSwH/idhJVPlEBnGz1EtFbUYvhC2rvXV96Ocuc7O78Yp3w3QdEnsOPcqyPo/OLft7G
VxygYmqIk97KxWPSddNu56FJvXEyV1M6H7n3dXjYhl0acvfVid0649VBbIuqi5NgSpHmEdeJCNzF
169c50XMQe1A6FAz5jJgeoSjeiBDD6HsWDRrBl/oG6b8H2CgKxiz2nXuew9fMnCAC2aPlpYN9SGk
hWNwFOF3AQbJdPqgkKbqVkw8O75XYey20vBfjKviu+jHoqeZFeNFC9ks3GbczJ9J68ju58wy6Ygt
OyVGJyac6QpdjzNtWTYMq5K7wT7HicrzPnTDmWrwHDOLdPHYCr+8vCERkAryMgIdUSlYpifGgxoM
cZ5sV6W6PlQWUsK34jktcFgNa3HPNUq3S86bjFX0d0VViGzb959peTkxOhICe2K1/CrLjdgmD2NJ
Oj1dJyd69+Kh01Exu2E5Q0IqMFYAKsKbBhHKc2+R9rRl+/6nkgLS5GZL67XeLj0QBZxiYHcIoN/p
NDP7LRfnt/DToNLd0wF0J7TdxJrYl90Vnch0zPi1vopPND0oL76Nl5Gp8KdUNyukznfoKyBh8u5p
x0Uv/xXj64Q3TEXFVmbtsvkHc+KRIEbJzZbo4adeD49i+S37Ykywc3U5vEtOh449cQqTihLanSmW
TtKWjtzaQ/b3mFu7fcgtVz33++gH805zZi+RyLc7VWa1nYDnwikav6+QtcQwGTfN6kO+n7p5TmwY
jIm9awwOcuaDEbWYmcrtEfgIyiZwoyiFKXlNNopypnaLS6h+6j5e96i2y8H+7e+hNBPbq42uthwE
/YlI0GDUKo0t1UpnZ47jZUKS/AatOTD/oBcJBshnQYhAUGW1OQPctZCxlNKD6gOpHLGU3a0BQnA1
j7Y12et/nd46AqJn3fn+UkE0KWxeZM6dTzZqOV4T35d+MV5b7elfHWhiHxsAT+d5iRq1Vx4Gcxu/
Pp4hszwAclIGPxg/JDF47WR0U7bXf4VIEHoXKcqz5SqENzIO0HRCzyNjD5slh5fcU6XvqdQL5S3D
Z0rRJB5xBeg1rAsBqhgSfTBs42kCtx4ZyIF3Bp7NA08pa17ikD53S/0ZVphydB8WeY4qITdkYTMl
cyh6IeR4rlsUnfcU3HgLje7BNALUNCiueias7gWh9iYlqGVxeOhyhf5ntmy9SDZ2GoRFCLnUO7WL
1RWogwbLzEcfahRWRaHnBRs4cB4yM3XAOFocfx0n/xAtWb6q+Q8ATXs1uy4XoW0aLB1E7VbCqwJ3
D3q8HtepjMkSye/3TDxrYslcdVGg0xC67hRJ6G5npmgyXKmMzp4Hf4Qvw+KcbtvomcuxXm06XeyZ
Ae0LxZTKVHaCBKIkTlKL4ZsNuc3/ZZL28k0SIbGzHZyywvejmLGzAhorHwHk/fExlTqe0ndC98/S
aDLYQ2HqmZCm9dGt3fIz57hsPkH6G7bRfP95fQAazaOr9hJ0T6x8Y8ae0ShffL9W46/zLER6+pjv
GJpkAx+ZqdFK3VrEsnIxCk0jvH94ioCHcRD0BtU5mx31pXgFyliCfrN0FYcZgGgU04lD0lFVEiHL
qUUM8WOKYOLe33JoeDghXW+iuxOzJPb3Mlm4+ElY4X88mzxcJHHdxPoQJwWVAyzFB1KF1Ofa/R4D
a1Wvsc7GY5eDEe2jfFvl7KDaRvAh30yRrSscQHe8bHAwgKYgld9yioSLujanon1REXMdWeEBI4O4
sNLWv1deiEJW+b+qhHpNqmHdC+grfUK/QQF7cSqG7bGmTvEDH0/6TkZz0UsRPloSTA/7fMj7NwPt
4IcNbPeZC0dTZnuSQ8m/jd8EOz5ViPrZp1fA85ATuWsW4t+riKqRbqiWwI9GZSTYiWt+IFMARJ12
Zm7uUvOLaFrwvv35VgmaEuf+ZiRHDkhH4/GLcDT+NuOwZaY6XQExTDcLowELl5tE6WnG5rJ6d2Fp
UhX3/iEW5WYaBwQzN7zYlem2+MumbOND9eCnc61n0v/q+vz/1HHhreFGVS2vONhdy9Ib0ErfAOj3
PSaO+ywe336oMyP+Qusanqji+YX1RFb61PVm5fWA14KoIVVsVVHM3oPKWHsfz4YPK/ECtulNpRYl
2S/WlcLTsN/E5uC1CWzxoEtWcnsvtTEF1npW5R9yZySh5p9pLCWuyPi7gHc+9Twm3e+ZXqEBjbPl
NL26gixMVKqGwNx0B4ilsMCojLrR0BuwFYu+flERO0idtfoNDBlx8lWk8XNnKtjh+3IKRfs6QoKK
J8x5eqG95mHMl8z5pVB7j4kzzlpgng6vs00jB1W92Mh3PCmlVsUSgotjnR4OSuqOcPlJjdbUe6IG
uQaS8GXbwLQvfA6n+99cBanOkokbSUTTuya5PV415cNALFXbrIaRT14aHk510ulcGibOvhinLUae
1RbEe4n7tFWfdGzAgk1c/2mcND40ihOks6Jg8R8alkTNIJyHp+zh10/jgwqExVY+3x27qKNpktLq
N2S0ivBkGApNfIWAny3WKNC5CsZ/qliPrdnCwmIvZbK+AvCW6Y37tDQfMrdHbf3atYX2h79InUSL
mU+8QztG81Qkg5akP4aDslRr6oh2xqym3yGvycdCmJ3X6AU1yUyzt8dBq2H4W9MzeWeIdVWToMUO
cnIbw5vX7Ap1cO6LCkQmnEnG1sIFmFIBBAk+p9jQ93a5C6iOJqdXyrTdpwkkp2uXGH8fOFGrlRqp
9G53rQEbsBKx9UF7SXjzspKkzNa3luJFwMpYMAtm/3GgnkbeYXkqrHiVjkoVaMxUye2pujFZC21x
vbWN/Qk17zczfPaig7cFgjNhgHRVN+iPd/9ftjSEhUC2WnUsoLjMuYKysKtxGkRdvi0Qfduom+R1
V0nTCtUoTHDgKAv8nMo9JMV+lIZjVyAPGx6xmBU5PCkT2CDlB0//G3woG58BAobSjTCPNt+HJFHD
iXOelav2PNKJShQ7s7omKgggnOvxE0KtdQEDWO3oTvuY47qfDykc2gBlZz7T9kGNIzWO2S+iOAvZ
hFOq3LIuWKPSmHdip3ieicD34wIxJraM0SwfBA0Mvp1ep6zM16RhSxNhOVDTQpN3OQjupKc52YCO
FEwQPuYXJGRAqenY8Um0r3AMPo/Hxg0BmX8O0055rIkyA3PKXw7GQcu6qZ3GLawEd4FiQBB6A7lW
/y5nUvqRVxaeixhqtaRWulPbWNZAhG8MZ7JE1Qx6CR5gVdMnO+oBZL++bexg6Jh5ELSV1XagR6SD
K4/GA93hIZyjkExsbO0fUIWpHHq9gleYBZiKxEwzpT3eMNz9m6X+zhRXg45dXqGyt/MbURoByuP3
gyRMGCEjykwOk7tKKPnXZSNPBjU3C80jqHB2RReQifYmjg8kX3QQcrlcSFngyLRXtwmj+rqROlgU
359wN18l16D6+78RKeKMo9S9exXaVX8ogYT+e59R7g6Fu/ltvle0UTm5M1lT4TvNIWHmCWI2ORe3
ucJbAMa8nsdtHr20Jb/wMIJzIfAieS6a9Jo/nAepOe7j01wN1NBzqcsMDw5hVsGuYHrbIxLFeBiQ
F6lqAi72CeksDuA7x9zwpDK+koROosFl148nL63YxfoHh9kmCSSQc/qLNqb9LsMSZuiz9IM0I2Dz
KsIUVcCMTI48Kn2unhKteg98ExJGYxn5BYa9rMCJMqnWvLWkZrZOE2TBkTy3XdUbAnPESEGRzbfY
XrmlMCN2teWaz5nzlTuI4cbI7uGxKdmfNJlblzgAolviAv21fFpamdt3epaGR1UBo4+ZFCFdqOyh
glyvxFK73fWrMYO3RPA44/do3hibidpvdunnFJ9NzJr9v6JBiv723eXo7F0Q0BCFzdfQ06CCilHu
WZvPSRAuxfQLO8CpL5EGbFxibLEmYDge7JUGAyL47gSLKI1VtEdpTAgrDguPUGlNu6qc+okcE19Q
qoL+6/jobyjQVQ60ihAr+M8pCnYJepu7rwEoshwfUtN3FtBdCuQ8ln70YdRvNRruGrAUtLavtW8q
UcsXAtzjRXFzWIqtQSBwrcTgxi5/AcmYB+tMSukDjV3Qj8ptTEduSb96jZ0+tsh0kse6PbTzUlVu
SbatQO49oYkGYAX4QwSCmsIg+4dNAEO30VXuNhMuavREENoHf9UxAwUvSAyRgiEi5nqDK4LPUwmv
5JyLrMRJ8dY21eQDUCn8g+ASM5tzsK4fp260qX0EEy96wGZgn7lbFg+zb6OWzaVtTnRrXwIREqc8
uVEwu7NBBlEselnir+U30pJAU6N3WF3EfPBoM7z97AIo8AS4sn9WGswOUaQAUjSz29zkiBzlKEP6
WQs+G/mROQdmmfDL+ylcI5SOBALFgsXkyw7MfBwvI6vPHlLp7SfofeXzK1FfuWIhAQdjsoDANZJC
GoL39qNHhdSDEHg01UKLf6sh+Ju08p1r3rhP0Vaf7xY6ZymXSlD8Ge8dv55iNvj4D5Y/Sa3lQb3k
LH0NFEN5bzpy5Ct+SviL0Un8d0ktLPVmFT/sc0YueelOJQ+I7V43NHFFVNjg7Rk6cVrzeiIaAqQ4
dFxpfRsaRMJ9inm9UufxAjhJwRnz5rWvpXNur4ZGob9EYjaf+CXXGcqnW6OtlIkCmuziBm3kBqtS
epdHvRd77bwnGGvbeNFN3S8NzWIYIKDp2XBiqpuNora1gQNiuOjWkxMYKDeQB4CiSVVnEVhzceM6
1zV/gzVVoCfXzscR2PH1FuazBSo1+edfnbvVdKwsrXXmgEA1Tqj7XHswE/LEl4Cta1T+DPZ4tHEy
EyhdNnngiXZjsNcI3jJO3hjWnaJL7/qQx0fW+yfTvAa5wclleH2HVtyykeDnSrqJ5ciJPew8B8Ka
VSdKfyJgC0K+PxUWoFT82vB6w0/V4fK7WqI51bOBSWzrfJcPQpwW4wsXnRuTJxXb/e5lSBXqIDR4
f8j5Bxio3TASi5LKIkdKCC3v24b/zp8spBtBy122or6SWAxxD889rlAOaqEWC43M4nuyWSz+NRXA
X6iT2UZEBhSYG2R3MgVaFJKiUhoK5M8pd+3F3J+kIYQ9ZyLGuhw6G/TXW001z9fZ50YFXk1KnHS3
3TwzE6nN/iZ0xubrBVHOUBOdxwbLLBwC09nnmHefmj4mvusJnQoUkOnpn+DkzkROw/6WV2XuMqC+
oJ1zWvB3ZHpWzvla6qFI4/QDXBkQx+Rpbuoarlb3D98cIuSKMW2OB5dMRTG8RSMnzy22rbh7bNoG
MQGlskDwlQtvu0Od0ojl9p4bulqZeYYR2Rmd63Q3TYqAcdbtEGjfjOwQ1qVgYteLCo0cII2NEoX0
4arC57JbEnnOmgfiFVU2H7lS2ichO427sR/Vm5VBKNeZMT+ctQxlsomwSZ/lDFoDuZZtrTZ7SRya
CGa/m+x1R//Zgx/GFTTq9SiV3ywvMdmMej4N7UHMkcUavYdoCjGsYSajJ3uH3pcKQ0tJBiihhXBJ
+k5byaoXN8Xoo+krNgWTyQ/eaQu4J9tK26mXzn/1A3gWWMvN0qtk7/hu7lWzKAWA9iLGZvoJpwXR
x/qXn3jaX83vox2HOeE2tZYxNElykZB14hVDT46JRqAD/c9B/Nj5+xj/YqYno3rDx2ReqBrm9+E2
tpD2NthZcIAdna/XPkAGZ3i4NdX+z46E0JamJ2ls9UtN3sPNw0VwpSPIXnkkWIlmUDAkWqJoElad
F90J45cwKIyTq2ZHjOaCT/FXO9Nv4RB2yHDL4iSiuKE63sRZIaSRWRUwCIqjZrEcrGgNu/4PK9wb
3fkWmoGQqwTnVMihhglo+B5f0CshN4u3WL63CRfOCWtp1y1kdAcvX5+pX56Aqw23Ud/1+fCNCnTu
ItN/qdHbuS+7BkqDSwUpC9u24V5wS0fppr3jXi6kzDuN/OzEHtzsQ0nlTBoDMyEaZe9WVH5qnPgi
p2CQ+Dm9RxuI3UQ/AVpqm3/VhMscFERlMj5wYY/QaN6L7AApiKJuxNmHGpsUH6MkgK3QKyOrgiTZ
lK30K2Zr4U0894S8FLaT2cl1v7KrkvaVTCms6n0G8jw+bHxOe+yTf6rKj1qpyhyYQcVSCsPaha0x
djQjPf2aWdsUBe8+r7tvykvhKhVj0fY1XKLzy/rKi2N4WGXs9p57TZ1KyrzRCXvb5a3cxbaSQ+it
2gjWr6v9E/Wzz4PtLCH6kecZF8qHgF5tpyA05laDQ0pJ0GB6+ssstMFSK9QNsMf68vNUXweMnh0H
LsUOXomNTx+YH/OxF/zfg0590pzE1dyE0CZ7LlAVLSeuprEzNiD7/EOMBJ+WOOW6adWTjufIw+Iq
LuOoYqHgCkEFzbg5Ptae/+/wd49n4o4dducCHXoGbuZGRrChoP4IRldKFxwgcM+/aCfmv/+SYUBK
NEDxqms2BufyW1z1rOHIzzZz1uJl3pUxk0zQyPmmlLxFmUmFAIyJbPR2p+AKEkVtPji0dLqBo8Gt
Fzcsc/vCqCzhH0i0tTeHD0yUf5tpyGZRDE2E7MOGJp5wmVTbMeR2p2XaotFPplo9JJm5FvLbb0+y
69d24kFgx2ILEdzjGkpqMiBYtUZlR9xpiwu4/ij2QrHV7HUkoxhvdyi73cRKIDlQGy7x+L9f7Rlb
tk7IrhTXdm/WImpWvXs+wwVR1sfbp9pJT8gebakLcCsqu5OCYUK180IeLPSlTUcsIxvUAd/74T1L
9oh4NW3qRr2NUA59QDkcT+x6erp6FUJsV/Gt1uugBmHBCTDWoem8/t53eXMVUR1gyVs9Ps7Ce/Wm
9FKltvRnbzNgSisddweiKVK2v8Zez5ZV+Y7T8GmeGifkkWD8PN7CxtIqGIx35pogpDJL8QL+R/Aw
iP97ZqSZfqBTHy25f3pFfrLncR+ZUb0POeZyaQR0Dxc9/B15xKopluH4iteh/JyIxIN+NEXEo/zo
NXQx5+dlqOxmglksowKDubmVGcTjFRzUmUKcCLhXKWmonuojOSPF5Cd7CnjJGCq1X+Ln21fZPawa
MOpC5eNDtw1j72RJ/y8CY7eJpKj0O6QFFawBGRn6Qm+pXLSgOqWZJkXTx9d3K8kPK2RJg1dhYpDg
mKok1vv0um2xBK0j7ve+dVKr2OQ29JYzgl7BwvC3PYKTJMmfyVmJmNtaIYuxBV/uea6hjj4mFYNl
3B/tYS/GDM8pHCtENodeoMdM1F1parqaNyOhhannDqJV4MBTxWXfqHAKYA8nQECji5erx5swNk0C
iAXAs6UWQz08C2DaTOpQ3vYnUMVe1/V8qljBS+dejLlohH20uRX3LtsJPjYe5ud8PczqZ8i6AHan
rvZlGN/m1hQflNqhvqXowO4Tar6AYtG0gDsv61mNIlIrFVDf1Z4LtiSOC2QyuDjlbzciiSeYQIrt
Ksw9VmY+MooQI7qAWH0cZge2rre5u/D5aX2PBnJvn8DX7OqUg8iJlHtUZQTJDpyPzwZVHaGiAWrN
h1C3KPUs2fO1pQHmJqUKWmVtNzIZy95ld/SDEvbRajmR0oNVeCwbypJcqgOlVJZUuEJVs6J10lAd
j96Q6r/HC8gc6cw91+njkTc33dtNL5Xa/zn75yRT+W6102ySVjxFnCVUM9Wo2idWTGq1kwVXInWa
LRYaFZScPpPdI7A2Sc2bEC1SPWVfzS/qGcANMyPDnCoPMKXy7jvP1yM29g+0hJF26l7YIPZ5FTeq
SWKktFG5svRJjRvKk+Jsss+8l9NbHhlYza42dyYETnZOzPggvWcaiuECsb1ovn6kXXafK4Fa9aN1
Uy/sQjjnW9ZzuS5hURiDaX0rKcLj5AeQD5ZGTBd0Al+k7rziIkUS2UAiC2bABzfjbjfeD+gO31bV
ITGB2/o09VQZQbekacSmRyv21P+VgG7JlDeXAWSU1qh+eyqVQSwK5eZixued6SRXhIC/jUcDswUU
sp0YsWKCQSmy5qSpLNb77lDXx9MvoBL/F34eO+s5IRtCr75YQEClzel5POIePpSBTagDMJSiwFoT
CR+wBb3ESEzZeLnxrrFXhdKFw2NudrIpHMqcPQXl1vH0SwIwKMn7wBnIlZKQlytzBJu83+5nERus
0nE5PVtrjREQmynIX7gV/Qst8WhXjn/1dfHdhQAcP9mKwtBDpQUFvnoi/yPwXtEZztdtSLCZEFNY
gM+W194aQP9a2ahAq9fGywQs0nqKGI3Z9CJ8GodOZhDrsP5PVjYjDXx8kqaq9usU2N1kJOjsxi45
hVO5x3luXOJev35bbH9MKf3e9tAAav/GE72X1iSnd/kenZCeYEt03rf626YsZTzPL8n52l8Y2NME
yLfr3mv61cJxig6e9IafBS79BLNsn6mFyXnU3WaajqZE27FFGf9sxGUgHIHyTjKyf2/DAjMShDbr
JEfnu/9S1Inq6nZqhybWZOAQVjyVoLOCohCJIto2woIIP6hOeCQmc6lUXTeWBw9SRfOZLrpcqA4o
VEBtBfenmySUNpQeznHLW71KEWtz87vtFh0Yo8W5WwgFMI+4uj3SRsTg72MgiRmHhyfN0IGIeXga
yO2TBneyRKlzCEEbPW7l4he1AI+oQVkBncj/Dem9WIWTxGvgX46m9BD1m+xuT9H24fnuc4WJgIEF
CmOj84kbm+tYu1Q2L/fGqR7cAE7EC0oXthpclZoqza15mBx170vaLRU8eZTm2ahVGa8PXIwUGXXX
FfMLml+0UYew89Ht9UDz7fxqm9z+r7cDuUOAwnrJrka7Px/nUWRy/w4VYKU9puCC0E6TS+Mjsopj
GI0vo3LXeyMO6X0bGs43xyiYEmbQjSjB3EQYYUKg0q2G/O8OBQJJlHt3xDOkgP0KD8t5VLrmZzFO
ohRJuA9rslPJ0O/ExF5W+WCVlK03VUGjEFyAf7gkxr5e0ci8EpT5MCUpCzUjS08UUw4/NFz0C+5F
/HrwXn7iHLT7OtZ7XyKNg68jONYIXDHTgssfLj2Lyeh6GaEb770byTkYLXg0PmiBdo9dEQo3wHBB
rs7PMuypF5O+RIvKDn/RC2Aoykp4LJwKrO5e/1Z+QikCmkpCsv7qETD7yV0nzqK6csnW1Aew78Sw
hM+dj/GXlctDJB332b6iqDX0jOSzteL2DUD9pVd/LBwigqi5DK4Wk4aJAysbZL/uMDK2RDn+8h9M
zF6E2jiNmCkNdNic60FXku+rg/VWGm/A8yBsAuLJcRMknwAcx+VKXfBlXQJdkacQCbkl1unXAC3O
gA2hsnPXg0b3iMS9uZV+1pDiVX0HeHga9WBO9JgoXkcM8IOLseBviulq5fJ99Ka6w2uGvE5nbCIS
rpRNq26vvl6RA/DorpG5cM6PnqbqYU2HUf397v5hWGCXT241sMDWCsx0adVy2ZhAsPMsFOXj/81B
w09JkwUs4yUFN9i+3ZzS1hHzESwojwXuLrRtg59lek7yR2Z9epAq+OyHr43roN0YyxGWqbefh8s1
USe8cu/0EIxwnVfAXs1HcoA62WG4lWaVE/fmW6mcbNLvORX1o3lNRERNka6VI5Ik2xzVgbGuTMT7
NcDkQQOTYpL5Ihf/qEMQzXTHLtTc+kL0S9/2GgDlsBOzWKH5VG2oPKP15R8PGs/Zi3DrjIIZ0/4D
5fvyRbzS/VOkeg7wvnklL20lkcVGYU6uut4YIMHT7XGNXxN852qFxf/jsSgKtvKcDhiQho/uo9GP
630+qhvYOgedfKN+cJ6dH1jM6E+OJmWsJmiJPRaTLZ8cu4bHMRrKXk0FSx0M8G7jz5yF/Z8UlTtm
viq8/BRuZtpmjHo837mA61/CIZ7S9730QEcHvkOvHzAEtKzZHyNjSv2L6k+kw6dtjZGjZZYaviS7
XvToGoAP0+LOdJxoslVKZ4TPttm7+PTGxi4Cc/DSl7ydliS0cVhv90wmndKYs4h8zpGGMi2sUMvG
BhMNtg1LIvug6HqesHr8BBq8eNDn6aLwaX/+E3xQA56o5zGFQf/8Ee85ZgrGAvt/4VDO3E0dX0Ym
9Gi3XI1/Clyo0BOVxYLX1fwZ21cvVrteECbsriBdngGdpDDxcT7+KyOLDZCjYbTn8tdLLjBeNgSO
HqbC4S+amn++a7vMgpQkLeuCMqimJl6dMO+6akXb7rgV7OQwBo+rhhK5T7NVNriPsPmBBQBj4X8p
TcFaGClmh5BZDt+gIitNskO4qwWog6a+kk/i4i80mCh8rkDMVlNmBv7sX8Yo2OH51hmjHjnb5w8N
81EBYINW6iNcLZ2jnqJLSFUvnr2FBG+JaIzRYekRMKgt1GPoUcC50CnXqpFrqITzLJ4UgPliZ0bN
fbLV++aUleJUryXqmu7Uhp4xSSjDyVNhJuQajxwvPi3lsN0tKDoSm+hWYZpAW6qf37iUYji9cGHB
Td+i4OsTJU1ZVlpHx7T9LCtyLTyUF89IlkVJrVfULJ1PwrF/N7L50ZYpvsoGYXG6Cbs/HerXzTv4
Ht5A2MBSbF6qKB2Ky+rsVHw9lJBl5AKH3sXjxqdFviYHIHQPI3E1uIDipjZf4fjFmZA5388sc3T0
E1IgaWb0B2+bBTomXjePKXcn5GnUWDklm8a8F9ZTEh5itbwbAnJSdho6pyo4tTRFtf/+jSPyG2iY
WIi29tM9fluPi9xXnc7LVsvAKjtPOD8Js4CzdrortE171RURuSvftS11V/3wNetsBLJGcGqBTfqG
euvv1FFmC6CQ3/LG5qm0iBAGIlUS2V5WiSZyBF8Skgtnk+s6BE9bqbIJdCK3bK6ZEp1DgzfXboo8
v5V4q4a2eHPTyZhmtVrhbFeX4Y6FIIHYcisGHf/h0RkmA4is6na7Ua+CXbZjhHE/GQjzzkwSweWz
Q7mHPPcki7AvIv3dzDlUYWghk0qgbFoXj12tBDOCSkdFheNeYzTQmLfWCBUEu/AEkUF4HIP9aavI
Y3dsBRsboPJG01KvfXACIImAXcfeXgPjeoJJWbQCHKpqi29jddsIbzuPxdaEb1oSquwo/6AqifwM
LBreI5KL8F7dJgHAK8jrBvYC66XuY2u5rK8/kc9XoBaRtvKUxJz4y96boF0CKi187B3jlizLutts
I8MQaOxEtspEmr1PSwdcqr0u7wu8qU/70qP4s/ANL9q8+MPRF0IqxZElITh0uG6U0ue5rjkvKRAc
PMJ5Kqmr5ipicWvSZhliybtkYF9lby++Cs7ebRpyJGlzRI9nIzelD2Ov6mURwetx67mKR1AyiocK
4Z/X1uVyWMQY+jNGHchYWxjxsPxHQXl+PW1JKGX9K3MpfgVH697YjhiB8+/W7VfHmORNf983JI/y
cOESVcVf3wpKHH1su0MR5vUEa4OP9tUcpXb8WGJESj0rnsZ3t57Q5kJOvzOKTvQ1LW9QwK9cE01j
ZgatBPWxRfXMV2ctWFWNw6UH4el+nb6nJOep+q6OaAthskmxBWwEWRmcsNtYlaoJURvi6X1bCWiQ
36gY9y1QobM50MU73v7D88AhJ2A1ptsoPj4JbCaOZ+hvKjM8SXpTebs+8a3hdExhrh/rZfMbJ7Jo
DzZEPtOQrhe71+QelQ622suIuP0N0U1t8I576WWe6j7wGsnav23ETHxCR/9/9Ssea/6bIGqxWlhB
ZIcOpEWnEsBwY01CdZspuJKU5NeR89304gO+Zbc/Bb9kQP9fieXeIh7x2eXQrKj0g6Bsatg3YBaQ
PUT7v/Ris/Iy+soaFmaMgcPENc88KsHp+OGXwdviJCwFzMy5QzPZKM1ygFKG2ndwOIATvCmaNoro
wVb8GVIG6hM68O7mUa46V7k0k/Lj4EzFOqeTx6IRcuhdeq+YxrxhC5r6CwHsnJWA36Z03rSE2TyC
gUkdN/TB+pQ1lGdgY6NC4JB9FHaTrxWJBrpLrMFlVE7h8DggYLykH9VWbmxDGu1+pSi3mTMDqknh
5PuiLpv7aQQWyvoV87Vz3XPACkTTyX1sS6cRz2jWhEPfOgAVRUKqQa0d56uZy88zhbbcF2wd6zRT
EDtspO9zC5ksb42htZnhMouCfUqSRNcI62RzeLEv74zshkfUYlYHjhHblhhRO/9gDrky2Jz9Bio9
Uti8pqIYR5YYJueKPEzE2awhramIgk+cxhpjCIwusEFLj0LBsH+ayGCG/UDFN3VS5N7QmI12t6Fl
Umj89PEK4kfmbdMqHgt6iR+0HSlQMgf0/iWR6HXwbwmdVRGDgqIPaYf65O8EcqNkvUA2sNad5Nn0
SgNt+88VNqfLb8Iuf+9c9mdd4ibYJMaONtjOPLWgaV8GlFJzyC8xMWh6m3ZGf9E5i7NN/nIaPhm9
EE7CojL3naQuVP8cBc9dv0UsJVClU77HYJmm6MdGh/Hng8B2dkS53y7gTEKSAmOWyoJiaQujE1W2
vC9b+kY851JuSN0DE9eH5nCfZQh+zolRQlCC623NkvoeUT8OlONy1PqK4mjmax0BUDNIq9aR1WG5
Eq+RUWz03Mtx2PQNGt53UKNv+VHiH8na2bDajnxklQ5jmus65qnzRDBoyLxJUPMc/QiMXOZmSMrd
oF1Uek7+KK7j2RB67Z7/A7FYt4mLRt3TUQFoJGr/hCF9+iRv0O20fkBcRL/h2+5XW/F9w0sSpuyH
mc5mscpGp+Dok6zjQPjXGJh1KslN1LoLuFttR11iZk6e6FtQadIe58FE8CdvbV/BkPGULTkGwZYk
5SKQ+/P0YQ6979i45syfC/W/WqU3YbEMKOb7erJm0TsKAIXqNK0hbjeppq5lxotcLcbRPenKvvDn
eve1tZXMEL+tIWCRYtjeU6MTl0ankEN+/kYhszxTXUIEiW1ecHDjDD/q/aTQ7eeQPi2l3z/p9fFT
VdNUxnQHgai7EQQKJ9rISkv0LZctjKzM1GhD6N6dUCKoBYqQWBJ9Tt9+RKIgZsmPBaV46Pfopdl0
obXdtiYNrDu9bn2xQtozGfVLk0QnsZ4DRFnV3wjQemzg2EFPZ16QMU9Orz1Tr7TfUHEk6HzM43A6
VfWGMaH+6sP/v1Ngk5KXww1XBzYG5UBd+t5+oqUGbrq4RaOjfk6iWUqD/L0Rro13k6612Z0yTb7n
ESgBvEbBZz6ilbFcFeyZgZVsqqjWgZpd/CTNzVzPNzQSqnn1HNPCwfCA9JtaQ7kGaFI0yebFC+yx
eHLA0cAfnIh69u5asZt5OAeHJMnlngzsLXvZq1jCVayN1srREc6b7uFdtaQ2tI4fOELd35K9MNrA
KwnOA+ZIJArdSPTFuLXaaaP2Q8smN55dXKnHhVs0Hn9tg3CCXHc7tHxVAu2PWHxGvLbOMOzQTwW9
VhGTP72vPSpuegEsqGQlpPqQnh4IbkB36jNQRhGZ4HnrzVNEkDnjoRvb2n75n+8oWxsQ6qqZVsie
KceLjxFznzugpwnrUe9QvWEkMx6iy9TeuSzaVdkq/xzBCYxq916xT9N8QG4dChalE+8ZgiTA0e62
XJ+X2wxgNpMbPPxrnsUoB/Fep9ZPehuuJO9L2/acYJPha1Qh35t461D1VqjpTwWkQWSPGhdsT7Bm
3eiMFNZtrLuqZIJ8gNlE/ZVD6Pbb2fsuFf6rVsRyDx4jk3LLrIxlkzX0s00wc8s7sTGjRmLnjvtZ
WvSL7jY7PB6mjbhxTTG6PzYaKQhMxO2a96NtuMOXUSMJSkXsDQGy8dIMFk45wNHReis49/25+HCb
f/NelqLehfCiu4SHZ3tk91KRyZtuNOCYfb2gKc/2JRzUzf2nDCIEisg0AgG5zmgrd4z5KCWKLkm8
iEE6tHuVxpL0nt0bhYgqv5j+qK2aglYw7G/TdEMOXXGDZo+HIKJZ0zcahASWQ59KA5TjMmUKV/qB
ewTkkqEU22zeLftA8MlKZVQhur+jM8lk3ELJX9gleCe5Bc2c5R5fl24WOPrKEnMTv/w0uaqprlR/
NZd4zNCzY+R3qovw7HuwKH3xkWIHkDBaV1F6ji29yF+s1wKdGIhvq/EQtBsr3nCjS8Tmf9H70ZfG
TA8mlePz83GdA+vlMuvMFcjjVEZWJsdd/ILpl6eXZkBqZ5L8Dy81bwYcd80OsYevFb/mgB/+2zf6
zIL3P0PoK+TWtmL4micl8fEM4UJdbUzawWAiWAE/gVzZpcwmLP8PJS0/X7oDYAKxZiw7adPtsSkR
Prfw8y6TU2aQahf5x9ajwHDRhmdM6BMFd+vj2Uz0wjXa+EJwCvi4LLihLCprQZOdnqTTLTJ6+lR+
CV6cs+9OF7KfEcX4pYX/VtDGaB7YyXZNUMJj/cZLjJMaTYNMCdSqzxMMD407LLUWL99jdxBKEuMR
HHCphiVJ6vTwYQqQNyOnWDOi3194r04IBg+wpzN8UhyPUw6JhBn+n4kkJkAt4owUFIDsYDFmIU2u
3+vFHvFlVaoGbC5/3lubEqI8ll2fI3O7tbNoxEYa1g3m5F7244ABNxg90hwSaZ350Q4N46UZPX2z
m2P16Y464mIMIDrzEcxBPMfTWvAGvFNC+Szkk0R5cY7ToZxN6XwuLnuacMIS2qUBZx/3nG9h9mB4
h6Axzx+VhTduP+Gzs3zydJQx6h/jxglE7/cqszrn/DVYP4X0ZnYOUQoHc/klivYOsRFUy9s/gUfw
oLMokjmh4t0rJwp561gvbAs5CPwJZy36k25c8BXFaN3GFuSp1qNz+uhXXuAUqDPMxgsqyX4zHRmo
hwEpDw+s9nNvUnG6JpeXVGraVEXMSfLeE1h6k/UWa40c7vvjbjd1Lynjo0MVX4WfNr8ss84kAE1i
O1Sz5R/Q6HNraRUO2J3oP7oCU1o5lcT1ZC0f7iYU7oYDvNcMWDZeCnjKk7sajy9V/3W8/pwv4IUf
JcXPZ3hvVSRctR+r7iOX275LmhB8D31bctmFkTTwuHJGN85XoGulO4fchyX18DOIKorzm4LMC+c1
rt33OrCC+iaefvRZ4a9mEUpLsEEX2H2gctxRj8ALLOZhJtH2gKNxYnKVZ2iSXAZR57Qfv+L1xaS7
hnD+1DWJQmUfbREJHOiaK2Bh9r6R3/r1nLolBTGVfSpptCpLrU3unXXBfSCsyN5kyd0zJhGftdr1
RV1kASJRVWDPZlkU8+UmAeP3RjG6BDk6HApn0T9kAry59B5r/70U9jfNSdAaPxowJkOk5D6IxMM/
ZnGB92BaSgeavIFdpdRaGx8SikFqXSE7jiWe/huXSrnLycJW6r4RCN/+HjvKkp/zlsJm5447iZBh
V3jpNZCvn2ZOjFO+sxqJ1hKY9xKcToT9SifPgvAeWW+mgxesmtetiTLG75H97rkn27cRK6Kvd1vf
2idvRYkj2UHe3r1nIOxkZ6/Gjcpb6T+1AQIJ6N37bqx73yeUxkdjiO52/aGtBPwYF8LoCA3tcPj+
bAlL39nYlegWNTwFduC/VY+ZsSaN1y/9L1b/67FSop8bTDhwGppnjIvZKntRJSCzRpJ3QT8G8E80
MwJAt+ki6yQzy4CKQcHRlNs6AIvCfDf0a+iqCxkEJA+qVNiASLsVpw9sX6FhmaVDy0Qaqvyez7S8
cmKin2RE5uJNuqGJaVoOXYNUTWpZqWDfMP69aeqwsj3C0ZKEMyFyvXJsJjcL++F+yC/ACuYoWHnD
uD/+F5eU6ZYp/5Njwi5EffG17j5YkYPod7pG4kvl/MRvq2E/Lj3nvMz1xwl4GQ31iSaQatxxNXjZ
q5Xh478fsB6k0gJm3pzDR+B1+wN3vCITLMrIjSJZeZbACNd1bcHJNWjrzzMLYg3Dq+hi7xPNLcA7
5b60Xwlt2OLFADcYSdHpl//FWFbDSq/gHPPEl2jeMWM1moJ+1g7qCh1vK37XCBTlHGXhZtArujTz
1JCUk+qJiJgiF001apv5hvMwFjhBTgkpCdQJpeKF7hzQ5eC1xJH1v8PEQd0jKidCJL9VoQpc42OR
k09bOrQ8sir528Hetzts0N63OgZa8PDoBOTiQQSbRpvDxTBCKIndPFnG8XVLWUNuF+Z05NO+BYRR
9dU2IHVTVC5m2bpveQdYjUIZAkyU739jRDZBqcyXDdARM0dtv1X/S5YD2jLlfnV2S6W+xx+h20q0
bD6aYRusgP6SIZlazZbFTk/PpUH3BLrSc1KyuxqEJe5gb5YqwewCBra78zVIQd8mmwdDiWp4MuBP
+9WMiQ3RafijGC/WSCvIPtZXhi/tCMyxbYadZ9pOIU02ZjVj3naO9MlVBw1K+7g3muxuyDWjBvEq
4NXTYXcveQcKa+nPXOcB56F7wDf8yh1dIPTXEMWV6UN3oWQW5Ky34/1N1NWNND1YXANwGye+DhVE
bmFiJtKWq5+svpPXWRj1ISK3hGNR/oXoPTJOHiDMkqCcEbzKN2RrlZ6ADvzxyuL63kDFdNOQQGwD
eOg50/pNKajyVvW+Jib9coGlIXjtILPe9VsM/mjvNkL0OqkigTHEZIAyzZZMIXCEqd7LAMtT0Ai0
rfMlhIubCxEINxDxmwBPW7MJ+2QT5ovsqsGMz4ouCAfQG2HhfmuqJC5/6oh3vrDk72+VCNu/0FlF
n1udHrTCOEwBng7kJAz76XrNP5ycycDQMesThj/EPvCttq8kI9XPRP60M55p7bz2PsaT5gb6bSWL
z7xEP9QgTbgzAy8Nh6YV0ffqvrVrKMOYzHhIA4zyAj+qMHHyf4Ssh4EBWu2RsBUbXXEesOXCMr+q
SQcknjOBI68uV7hkvxLej/7Om1CHeayChW2rp8U+zaDOlxPg3AKAu7mj6FQ4hPaYB/4pBictpd7Y
AEEQqKiQ8tfIg7OT/Oc75N8+fa/4cH+4Zc70gxXSgwBBBRZTdhBhOHyL55P3fka1S0BsNcRIEfej
kYvyOKOzSI78tcNDBImlg2JpCJfzLDchyuHXvzh/9SiNPBkMXbWdrSzDZtHH3mSi+n3vtbtCLHo4
8hs2Ze+1wcd/hzmpG1dVvB4cfz4cbNg1FgryHpkc10xHqanIa2sIDaD7+qBDbqFwQvas4KGL/TKA
/i7kQb/omCD0hSUXvhz2I1bVyOPdC8ceW/8FiYKug9Bgqej2TXn3wcQAAm95wbSqMGiFvDiMGicG
4HG3upW/RY+ftuKTX9hchYOOU4b9UvAhs2HNv/h2jATDI4a5DTD84+P41ionqcIZPBWODxfDKR3n
JxHvYMo3kwfWobcF1iKkkxJbUfzyNJLYNE7g4LdNrk/CQ/g0t21QpTWPT2UaZGlz+J/ij9ciCbZJ
jKN6Y1KOSAta53N83ot/+P9eBwz5sqA5b5SGvS+78Q3pb6Ga30EoCWzy4367UXRyZe5IldkVWVOZ
PhYO4iW1oOQdndzyqBSh7AV2O90erW/aEqWA194FEprzffTUN5oKow+zjjaPXNAGSDuX+jJ44JQ7
oH9lah7lY79o+NUoP3QOI9HiEo9fEeowgeD3lS2mlMKRGrUJ/W5VIL7xfSBEK36Fe6aL3AelWOnd
4hwO/Tti2nqRGHJqrn9zJo5eSwNkLk8vLvnzYh0Ui75fscLqr4hNpG/7xh7KxHz+86/1A6NJZYUk
pr2etNxBofgvzuH0KxdLU0R7etzFmj9rVq1QcUI/sElLRecj1e/Rjs1zBNFLKaHXF6em+xTpBqlx
g9VisPjW+Sq6OSRQq8aJjk+fkCT1mwMbwWRN3BV0xN8+n7ZKtx9Pjg4xwpqNCSObFk65vOFe9DEu
npQVnK3ddiFK+eUOn5zhc+Tkh9jp2EIF5C7263yUM8iytT662x4dpXYfA8kMimWkB07trj9L/AvD
XV0eEnas09Z/R0mGd5G+CdZEaM/f87UvVzlF+ZXqrp1X04fyGDrMaAFDQ6FePKRsuRrlRLUNPWaO
aAgLdwkz4Z5L87fUFGvoK4YpE7nK5FDn9ZAvsxEMqP7SfdpBgyO569hxE04eBB2g9peDdERdD5mr
p/S9lvt/H4TDq+HQxCfug5WdXlOc8OIB/APwfYOv9d1THF5kcc6pg/4iRAwvep5+XF3V7XgHTm65
+bBPEuhRnatGJ7aw7HefguhOUWUn+q1iO8oL4Sidy3NgETHvXLM0HEe+H/cBTyl3m4dczF3dc5qp
tauiNgIhIVZTIALMp82a5Yu7leK/yyhUvssz11veT+PWaro8vKW4NUHLHHGpYie1GKsP/Sap5b6k
iSRg+FXs4fuYKfFNLdARUPv1pwo1FPhD0jcwVdCBqSXKDV8hDgIxfkxmnkIO/Wtv4fufk97C1f7l
doqPX9rgqxjpNORZtqCsxkUVF7+qbi1Tfz/BOWLumlOfi7jljAEnLf8j/Lps/PweaEZyXVSAs8On
PvUhFsJiTwAq4JCytYQJpn+KLjLd6ZZMWUzWdn71px4SJsuq+TEGhOshiqJzio0D2k0OA6D4BRik
p38YIuE5WWpmc1PqCFxDYiU6JxKQy6v0VFPUAXRpFGeMijJKF8LT7TyIj1qHo+O2WKCYLyjX6QxZ
SjCRNHQIl4UB1jJ+LxXGp6KjZMWER16Q/agq1Y+kEjPlEi/zeDJMh0YQbmH/EXB8rchnPMeFHH/A
0lVBzLelLqncMeC17snzXPnzaILzB/z26l5ibty17cJnsjLQZKKvggVs4YLXZITsYs2cT2ezLeHG
LAOHEBD/cziY2vsFA5CzQSw9sDF/qaKEDC8XM1mUpL3SjbseJ3UqI87MT2vZPJpXwUrv4Pa2+AYR
sOGUDdjS6fGlS1Y5Pik8ilM1k6NkQJ63Q4DiM17Jxbth/I9JLgJEfOQU2XmCDKT3V7qdmR3nqJVi
Y8lF91c2EwUsBE3rL++2OzYGxlmHng5t1Mu21uQFaSq/n+ShkWuQ81CpNY5QfI0R81sM3ezbsmBs
8LhHCt5pRBu00lSEFDYYu4VykHV0z73sDfGyespMNc1RhC6B1mxoYtsWNaWHcQju099MBGBiL0LB
F0K80FDQUlSERKkpj21fduqJHEO4SivThQyjc3ehgk0Yyv+T6xl+Wr5rKgOADkHiAmBz5v5Hl70j
T3Rru/QsBzYMybrAA5R7czfgELk9V7BEpoXs0qpAE8TgVVHQibG3tto3hQryadgFRvUKw1e9bkh8
E4mTGGvC8BGC6nXV5u7rqQzFAZlcSknXg+958hgFwL1dYxzJ44/MbVNKscy5UqwN4Yz4F8N8K6mb
phYelvt3sSFOyd8A8Np3fLHfUeuJGNrBKjrHTKxDWTOOO20jsHHz0qsTDBd3zwdctob738NXbweo
kreVAApPyS6LlxuSPTbo9kCTlOgdext96fFi01+Ug53uQnJi7BAAThKwFbfO7OsBm4MD4EhkrPdt
dwpGYZmjDkrW66p38/wHBykSzoKEOktuoG9xnIMEAXLnVwp8TsumxZaUwRJnp9XxDssTfj1USdxd
fPj0bCfFMI3B1OeBc5ADFiogli4xVbkuOPU8aXDi7zYvJJBtDA0qPRx5uiUBt+jMjjoex4ilPFCF
hLhCC9qGm/SaA89uvQdBBd5sdCknC0FMdogQYPg/MI2HfGjaPNA/GqQFVRZ8kvlHVBEdf69VYOCj
8b3FzPYc/f1aFxZ7KkGB6frFJ3WOAThZqjfME5Tt2A/xyTWuR1qX3wCLKxEToBkVqpBjFmgcchzc
J0Zuch6xVdT8mubt/Hx34Z1TDG7l8KarW09NAh8wxuwIkO48zZG4fHM35phC1vhrWCYUWGf4+0Gs
FqCJED6L4p2WF9d8MEudvqrqJsr2925NB/kcyczkgf7R0Oj3O80ha5q0MaTU5g/sg5XuX5kaSH2L
oEZqbrUpep+utd+1SVpog1xigXWV6xhzVpufEVFOtIXrA7h8m+fwQ2siLEceYOXGt92tYeNZZqGZ
F1CEUvTqPAEXV0zO9cPaHlFoTMdCvMd8fCrThQF+mySiYV6io7NI6LyxZSQa5Y0LeqRR2zfz/D4j
GNgzNOTluBLqtzlfxizmsF3GOYZxeeRcP3ToNzQK+cRmYoBO8eSrSvMF+gQmlS7o49woKgIsAyMi
9SfwcVi/SmAfk3+T+TGoakgmTROyhmKb3XsMO109c1F8G5vqGzzLDsZ8UctTt1rGh4oWxIlsksnb
pF/9FryYadmGJs1d6bq81CuoZAl/vwP6k4M/UXPfM3s18Y+sw9m1vS7JtUTC2FHWuASkRdmmfjPq
mvI48x5mBtDKE306cjfzFO99Y5f8xMdvmBF1scvE62No7lD2rGQTKwWgp8mhUfViNQ19BXVJGeYn
+id4Y4RTuzPqXUvYlZMADkJie9pCqtNoGKEwi/FoCc8HEu6Ew2TJ7+XFQ6/KG09ANDradmqrkXwr
FYmxP7E3hmz6ALfOuYErEM2xy/JUzodLbZwKURm/WoPH0b3tScvef+KXVHKrE8Nk1Db0CyrMyZqT
Zeb1calFivaERGyqfzCZHqcXWbaADLvr4ZrVbZ4MyhOvTitabYjR7x4Om6ytZXpxWL+9DjNguKPy
k59i/Yc1pLSfDNFLX9254ZnPkIvSdPCpkuH2YXAjZb1/7XN76n12QQtlytcn65LCtNQrl95V593f
6KQcR5EEDJFDqrXKYOwlg7XrxaQbfIXYGrKRsy9QhtcKs4S1w47HDkb/obbRkuFHSPgi317dZVs/
jv39IcT89CxR/LmFaCrhoyKbRwzXCjmwz1QnvgicXdSO6vE8fK1Va/Tdtf3vNpmiREUyinQajjAC
W5QfgGLU00d5eG1K/NoAuBugPVV3ktYm27nIBNENE/+/HahYO9qLNc4PD8B9+ze20NAWUmxdiiQ+
8unXt+MNMw52JsZ3Mm1Izq22hFrBUlbBJxxUxHdHHiKCwZBlH+82CLRUptZFj5pknJvkgV4Smc5U
uVMO0di4fnsA7iJNw9lNd5sgq5ajmrSeLBHJkUmUabq2zB2FSf8psuLRrdO7YURmzQjzbS7z7Rzr
3vnJj4xvjRI4bCpNlU5yScGsa3CDZpqGB0CTb/JelNv8959taMYPQ3MuswRuxwvJBImzT08PEiu9
nLmMazyz+N3t9AfXCGgj02vMXqIHCngYZ46USMPXRek7lRXzH09azzxk6jffWps+/jb0HmX5DtRQ
00B2YzjL2wk+lzRaNNKJH8SXTsIc6iunjsINSjG3/afP4FSDKBkzko3SFfuzW7Is1wXDELnAryEB
EFuMCyBpjEp1hopbzZFF2mizPiyhLiRXccjbAgKJ/sC5m9SxQMobaHsg6NU5lsRPCytCTsIXdtnz
VcVQ4xYCX9CwOxkK94zHsBtwnww/m03A+P7CMOXc1L2WPNpboRazxu5bp6UpxF20IqFLixiqRsE2
hYBG8ssNXzQhruLE3aCQpn5oaML6h7NxB13+xQiAvazeVgGyVm/HMvebEAnA56tmZw/s7MSnEj/G
asA1NNWTW4nWsWKPrlcvsHNIDcREu0iser2N6rMpCSvW7Sxp44a+h4nIcre6sr25hjKEoGWUt3NO
NJrjpxRfd5jDVlhIgEWyhtd78M8j+ZTKgiqLPFOsVcil1iggQ0aB4sQ2htEDOmHdcNr/F6FM8J5i
5k8Mt9BGs10nh/CQEse8Mv6n86bFo4K2JsPRo6u9/nCTSFD21Gv6ppSMmHskZwprKusn4T7zEbWk
AJ8mxDwcTvy8S7CNEfwsBNoIEPQAn0Fg+UbbIedPs0HxWM/y6iOObdBAry72Omlpa16vWUhcYkTn
njcYCSXej/vY0KdeGNcFPjaiuoYeBBNQPgWQn1x3/oPyvTe/3XQTeCxafn+aVQ8eAa1F4NroaO5s
NCbnlpsO8cmOYe+qsSh3QxudvtzW5fS+z7znSrbCvNhEqZOr9Pa2GlqKLn3jMJtMCqoucZD8vaq1
tu1wgPwspwNLjlD3aToDQt5HmyNH0yPv1wkmpzg8TayDESzAbVwgMhb3FvFXC2bSrybZ4inwU6PJ
q4tOYKmfSK7oa4ofxT1CHH/GC1gKbIy6mFaqnLnn9Ms3Sv2qC/ZUSlETg1HFgB9MWs3oh6lRjap7
BKTs5nivAl9Mrs+/soiEggBeaHi2zUb3Bidke22WUnlFwtXFEy+78nt2qQcCE1GyYjCgLxU9MQhf
8eHriaXt5xx48aOLOMRiUm7b6BPRA3/P+gm9crU2pLogX3m0OSKgPdaUK0BeITLKBiKEWV6eXil1
dR44VyKWdhCvgV82Sr6aJFa/4X/oLU6U6gfdDURmNt9zOSSQfP3+F4T2tq8Ag/1WBiDMJ01IfTIi
1Jw0fl9rFiNLYeu5KN6tQFFPrbpbjUXe2eba1UZHujDMtVwzTP5zci+n7rdAtoLEn/nh6/OJStTB
gvQ7u0EMPVoN4SzlEUr9B2AH0FvFEv/VPwWK3Q5P/YKcYsaleDsjs0E72osDbTZPn/eZGi7QlTYP
1GNYAww3gcVlVR0e+Ec6GSYpATBouaqNUHvELvmJddZQu56ZbDKV55FKJsG7YMUytrkctS3n5jR2
OL+Uxv/j6MusZREB2AVCuHoJkzC/k4zK8xJ1JTQFZulknOTBYiuU4CR++k15er0EZPivvQ/nJNBr
OouStBsMJCzv81aShKCUZnoO9puCLFEcrlkIXyPJ7l4m3OQdQ6TCoq9/PTWFRkwtFK7potSqgr/G
jICy2vx7G9G8yMRhdl4cAy/8/H/RrlXkF9dtF/p/mHn4i+nrEoR6RKutWsLo2fqxK9KacxdIUDjC
PA00V4+gRzCDrCL939vvK0h/6tRQq5t9H1x0ntsTWeJODpmgIl8lN6ekFHGHBJPKY5Vq6/dRrGPx
91IjuAU4gq372VT7WhaEpqQkrDxfmXiPAp+WZQMxULxcL1dg45fxRwTqmfd0u0OWL0cwYrcMg6Z0
bRFYnUDJVLVncVWwLl1RZCXQUvfXtvYhhNqdTKYGP1oBd5rUA9VcjbYhKbnS+Zlom3ChwweiOxMH
n7Avzet01rPfCnsqRo7SpYR5zkTyerBOPY1PXYXGPNFM9i+P5yQBbHnDVPXUG8Dq/9iQblpQMIMP
LRBudoULAYyOEziOi7FODiUgKxwqz8LWR9JsWxQI62XThDBD34HERbeTbeeLhd67XFpAJzXPJ1ox
GutadVQlV9B8pqEErWWsiszuageH1sW6g70eHWW9xok4l4/oiEtcyHazIUqYotau4Y1V/QcAchGX
aYD35W0/zs54ub/2DCO11DyoChRsuqCNO37wq/2+kdhaaP+HqAEvUFEkJ1RHLagG3mdFkOrxEu+C
LP0SBoxoau7l7SChdBriPv9A8amOBhynyACuSAWNFrFd04+toJHFZ39fEM/nIlTvdfXJ0sEWAoY2
5lEH9ChCzOcH7PWI8049SWpO0mKqk/Xnt2Rd4W9SBM71OMoVbu1OHVkrlrPakUFYe5HzNb8IkvUX
79ClYHO42nuWEou4Mx2bJlvesMOATublvPDVqWaJB+Ye6rfq1yrW32+33+VKSi1b3rm8u8kFTkOx
GF776LlBniWV4KpJzDhqODno/AJ6VD2SP0omDmNzTqYUEOEM7tHCiZvtIJWsWmhL7922MdZRodXP
AhsYidEP1PEIz7emgsb8Ef2C1gD6z86irg4olrSwCEv+/+PdoPdEQtCQWvLGdtdtjOZWEiJ2YbG5
I7kBe8DEn57o1iPe9uRMXVsnzqF7Vh5X84Y0zQqMWEjiu1d1qsupHCqwQ6Gz6SJsZ5SxWidw8Vip
hqUHzk6AiyXJk36KiWPxu8M5b5RqnYnGZWNK6Ydpcsc1OcDp5AkovPEnKczYxM3SwYhIuksY991F
iKoXm5F1kUA5lN2sR2bD5Vdhy7nwT8d0jzZ2cQCYVjhqK8VpbHntVFCjslq8f7A0jCDr8WewtfzJ
ErrNj+Qjvu0PoBwT3eTM5MmbKQEJkeW8s2QN6XVggS0fclMs6XI/pXSlXTZ/bHzLmuadNnAzcjr7
LtM+bolPcXbRZBXtwVy5VNPvuW/4QJvu9ypwD73SeOnC5A8CbZkK09BiU5/htR0ea+VJFjLM/4B5
2YEBKvXyk80R5/IBWczCFD7aH9zIixnx7ybvOJZHFeStwCYWOZMNPVpMGe2Z2AWrcW58TkOttjrY
oO/anM6XHHm8DO893ensn+EZGYCybpeKTYKhJQc/IHLpHSAgDTUU0kEABAlocoUhZrz/WueL9B46
uGVEqOe1rly1jVPSaqIAuO67Aen03CtwPP0B4/W6gbdntMCIo6hjngmy0Cu7m3eRZUKD8rpMET29
KSz+6uxdt2NSbTe2IMVxt0W0sHbJ//o1m1rsuny39AxjcqBg9b+ILfd8s3QGMryqIs0oq9ZZKC2O
mRzFgAcXwgQs/IaCEJaoogvPwxNYp327af/PNj3ukRocKOhDxe89bKF2SPK4ZiQuB5tLBstcBd6a
fMMkiSiRmFu81kdjJX3OI+cY9ymsBxMjHE7tCbvpxfOmfeITMSiu2q76QK8p/mEwGCkHWRtYoT9/
Eh1rI+kgwr/HF2N52sRjf9yM+VfQNGKS+9zEiCMUtix0gma4tjKx6iYtzt9TVRTT6iCB08gvwYfw
9CMqdS32hy5x0vCAea0acQSTYF24XILRfy6q1L0UUKW3qmNLHcp+728E7HEJKJ6G5w/UHO5MbfUG
3Is9HpaxOzCej4J3PswLzMK8Ds+GCT2s0ziht+lVdU745RMyZLb82WRmuYsj47r6eBNXE2jCqsqT
ERC4yDHq3J7VLKHKp9iqakqsfCp3pypUo1hJGcbSnYhBXrwRaDNoxRIbH/O+DXbC+9o5AtSZ2Dr7
yxiLCqgOtYwd3qkm5ae8aRpzJsEpcuH2ICFwSqB4OmY/lq6QFt9/0W/1zwmR46ibD4lmeokXN3df
L+TvGa9CGInokgiFkvH9ziNl8Aeo1TBZBG4Z+CCYHYU0cxOh5MK4+xtOSGH/cIrBjtHv8XCHUTog
SMWifnwen7N7ykCNUSjIhGENMhD2rkCktwFALJVElptevnmXtiZqeXV1jXGU370T9EI9mhpeSVFb
yN+MiT35sYaKgnMknk8WVFfMsMrKZ+vchT6QlG2XXPTpADfVJpbqhQc8YsuKo+u8LQ+NaR4CZyjl
2hqwe/nzgl5UfGul07GCNBwu7ZMT03mf1WUTlUOVZgV3mGIgEJA1NNPeWt/1Pv0VleQKg4U0efag
JQgu6CfCTojccQm9KirgM0bU3F4eY3VNPT80i4QjcOc32w4EKAbkCNjXV9f2DSePWta1yHzGYIYc
yeoHewbi5C1oLiW+eM6PRvt9yel0iTnQoCj0cCGe8ARzgS5w5g9ZkBPEBeY5BWQjzbgkBUxe87Yw
+Y1URXiJ1IKcMO5tFI0T+b7Izl899WGVw2iatq0hIUd9ZYR928Bnv6OfY9lbHuzN6msmZiKP4eTY
3eWTFGEB19qQKRXLJ2Gl1oxmIgHnFj6/ySlf/DH1ZxHx32OWHZo/Zg5VosjRAmqe2vfDp5ugS0x3
5FesyKH3S81Biy5CQ2WQXJtssVkpaa0tuYiIW7Dfce9Ihng0taDSQWwWvuHL9Vdb2QmZT8yduyAe
UUuaxmxxxcAzxw0/7OPcu7qL6g/Lu6HI00lO56ssG85zIyfOpAdzvzVLoLLlZZYdffaCAu3DDN2U
2a/9EtZWRunXgLelo2O87MCBTjDPJykNRZguySYEeDidU1F/E2JfJ8lrZjSpR/w80glNuePfAe0m
4ydMCBna6R3/+OTIdog8VlZXMfCwkghzOfFVV3DVRjqvAa9lzQlYKdamNzldlfe6+9A4qN62RRBM
IdEV/uuvL79dFQb0XSQ5vErbSp5t50xgLDbyCMQqDQ6H/hUGeXVw3uY1c8NIijcoEIA0hNyIYJoH
9K6vk6IZJp+oebdVxsuxgN0javS/e7PlsN1b1n7bWWjANy67PNFmA9G8Bu3h+qpFxOg6kT2VJQgn
4Q7bY0+hSzudDgC50apk+7nXD8XIj0ZhBVf+BOdksSK6byw+mvz5VUeMhvarxipyhNHRtGmxtLUG
WFIo54xHc0vh+hfyxHgwHridpQDlrNvYvNiZuLvRa7+foRFUKHIO4R9M3AfmFY7EeIL7YDMCUh6D
ZJC54bHhI4o0EHll6Ecl22fG4IafWZBdd4Bq3Gl4VlPEqrsDo+gvOKf2YdUTpWle9C82Q3JH8qWB
UbKbrEaDsnDnJm5Uy8JVyum0Qa3dYFPpMoQswm/bRWp3A0Xsg0F3AbrjNnXXZcV8dsPmck5yICN3
SpVia+x0SsMT++11YUpYVdzPIvrWo273I8Q7oPS67Naz9hOrfonZGjw4bvSP0yGqWv65tLBeVLxc
R6aTVIrWAlWyBp2UsbWoLf5N36YvewnH7nWzmsETwV6XSZlLBlrMjNb2LPf0QoHWq9sC2SzUJbe3
Nt6SlvCyVcubBT4B8bhtA3gGQsimzreImkBRpQAwdderknzb6fVfxJL/e6c1XbaLrFUfYS3XauXp
1jBReftzqIdatqOiNd05ivko89IBBJHjWY1U5ppOdT6lYsFNdypQ9BsxU+iGmns1ffpFh09OvmwL
uuVapu4rPA2OpXaaMCLGkLoJTn5fZ7t6Uyr1ijnlh0bBqqcxWKkBwCE8ITIKg6bg48RgHQy6VzFO
QQ6WISH3S3XQqZVWsUnhF9GqjXAIMkXguqTM6iQgQWGHahXOi+cWoyVPig+5d1uUzrB268WhWCPE
mgD3ELn7PojSfsQmlLCEGQB+ta753+ogeL3dwwYLhzP+PQm3QOpf/psJy0k60J9WtWubfztKuc+V
DQwHyDM1SQC/0oHyP6UfllkGo5lZE5H6Kt7+vQznwuSq7iZpvhaT9P8HZNwVLV1tiYkCFACh0BjI
ko++06xRcgjiAzcrLvLPrk1k7yTEsj3IXlbmAle/doKzSs88UZZTG5byU/U7RikzApwBZ24WagA4
0/eXlwWSIFk5I0BABTWZwg722SDFE2IyMb4PXH34PhU6hT6liFdsAvK87FOJD7qYJzXtDa0Re+vV
NwGUCuymrz13opmgfPhB002vU8qUTPNEq4cy36zZBAB3Eb6Df8KzR52W9fQ202LgPvEz5LTC8Ffw
/ya4PZ4E8Vmas4o+oGv2cYORJBEoFpEnf86ztN8oWSPWN5qDXYFqNxiys2fJx3aVu9x1D9Njk5mg
XW1qCOO86rWblrGAjFAwdW7d/fNvIR54tCAN2kGpIx4uPTAET9ghLL0YVWRJ+IIA0YWHdxKa4Ja8
273ROfce2t76+HXD9W5+5+uxr6q4pDpHtIiMhKsaKjUYIeXYLFVlczPsUTatH5DqH0Fxwxsdjwvf
jVu49LYW/FbC15ehPdRsXf/UJCGnRkJ3amjm4TOB+UgIgk+uTPKwqEdzEee4N/f+FHKTsnJxXLCc
uhr8SYqU1HGhtycPyVToXIMPf7w6rwl8MW+jbLr505HwIPXcM/SqOhyNQoXx7YnryFJwdzmSzLcY
aWSDGi0e9oKCesTt1w/NDY4QYvoDBFYLG4zprs+UVMTBaJwGNhIDiIa0B8EJCrNOx+3CvNHG4A8i
syvWm3OkuHw5+ogHBhQI3Gr/e7xk25LDlmWmuCZV71r4BM03hFoJTnwgbEUON8n1X9yVFSBaYQvD
yrg2uJKbhEGAMTqrUdYMXdz6Pxkw2H8kZBcjE8z378TrgOU017PfknthC8oPrF73irgxj6M0QTDA
XJjq0Jat09bXTF8xoX+nSGVzbHz0bR8Ex7rpjCqU2hqJ98+45aTl6kP0fvGsqCR8DZVW81SQmtNF
zYhs5puASMOk2CiOcAqUMKrgDhumVzx4jin4u0U37ySnnEih7pqbS3gpWSyIZgIvMwdhSMeQqSBo
uWNNeEwHXeYuMBgSHMDO4ACtMG+QGmqlykpCtqAJJHnQ+eAvBsp7WB0Id9WHl0TXuzh0/7Hh2RMk
SS2ClsWSKHRsGgyCPzOfxqohBINry/euzIE6Vqfy/a7UnEnz+TUZb8jriB4y5Dls9efACaWoamhx
9pAHAfp8h+ZFT75pdOZ9BylfOrcTPYEK7n+XsC/ousSv7ly3sBp61tL2mMtB4Op0oZ+5CRRXmmjR
7ZlXaNWTzP2QlcsLejPC6OWxyBjT/Ukzd7ALBFDoQ3LWYUSZnu4WwhX6HAedzZ0wMo5Ryw/ii6VV
hM+3n/Gr2uw/kiMKHSqKvVqu+oDpTU/P5PCBp6Ol75+mAueZpke3o9IAhUyRnalgzd6Du0nEfb6T
6hdXVWXHnrTq0yuOIk4HDPAzi2g6iGQuPFteRgjsJFXSUBUISDvdrAcFJxpNFMjrRuF1gqc9Z2NC
vyfbmh8zfvRLpqXNxKdmr8x5JaJjCElG9qrMLcGnAzT2HWyuQZ8BNme5WuuhfZkfRgvCEfKhg4Az
aZbJSbLxfqFcPV+FtzmzrlOw3gAnIAoGmomhF4QukoFNAdO/o5s88Igi16MNOC3FVmc+DsmIb2hQ
7ugswxxa7yfx+TAgZs+y/6gylqXJogaGk0YAuAvUE0m1jBDq8ZB1y7UpSmpeDrG5uDcrg78682/J
Oqa8/x35hVTfVRDALoQJzftEYqJaZ0NeT/Dj/VF0SplFbPZBzVwtvlIvA3l2KBzJAYD108LnDFi8
Z8foF3LgJ0FUNQOQS6+csgTUzDqIUkvzrPE7VpGZZvAMR6nu7DNFIn8vlZxtYnx+rPFDAPh3S13H
Bs1zrqXO3X52g/dc7ycV3EuETHX0lkA/UodnFzk886+vpjVRiKkoIRZm37pu0XLwiIPG0cj3k94e
bRyyH/ljCzSZCCnOIL9kekzfw8d6fjZw0afLu6LHt7jT5WNqH4pUrhqoaOJ9DhPiDeFwFXGwjkTM
r/UGaWjYCEtcVM6KzTl9bSqVtjE3ba+MswM+GMS4CvSjLsdMPaItwl75iEmMWLupcRL4j+VTFpzj
azFwbNQGLaW3jLF3uJUz7piyEk/KZ7PCdEmPjXiB+cQ3PSXQySCCrcy1IlT0CgxFVcoUeoZW3PsP
1a8yVGHZQSWZO/rEvJefhfHV3nEdY2XenwjWTkj061hSOerq/RsNwL2hkblXWukUvUoTTCobWLmT
PqYnaUXfKtCBFSorN1QiDi32QmLUw16HrkI2AjFOBiy2KVB2mfC9RDJTIIoTKy8L5na6fWTMjb8S
cAphroPg/0wxW1egC3kENCHFNN1bYQBaneXNtbvJkEreE3MZQmn6nvySey4nkySXxCa3nnpQleb7
biqosFlyCd6mAyK5G4Ys2iZELV+7tdPU9yVLtR3dRDMWMLtLZLwNNoVrNZZgy4BsYNzftu+1L83u
0xa+fvui2v4DjgDuUnmdtH56cXKwdiFq5/7uXIqMzUvzOcojlvD9d8JjvIm43EyfkWr6iZTw2RXG
R7UzYOIOMWzrSgCuCCCFsJLtv8Xr9s3nDf/fXmkoQtxP/PzJzR/N/hd7WGzJV0j6f1ZpoqDcreCG
MpDMd6WDUCHeznUuI+UrLf21WMFAPmZCNeVBulLTFqjNYsFindC9XQEppBS/7C83e5uK5rMV990N
fboSqNtljpa8YoObaCcp7oqCS54mPv9zK5LKSZDXuk2wy4Gq5aTdtIeQe62qNlHLg0yRllIXg3Ej
y1Hd+lCU6hDzO1GHnSDe4ClSym44zSeuWrt0W2ABq/C4BBW2RZ/SMN0DOxSGKUFhUPsGNUMY4/UQ
Bn9ZXPuz3mLnpAn7FD/cttAMnwoLl0UoVwzsdfABSecpaV9dO4i7Dicu32pAMPU6sdmYBfgqY264
XX05qklndEYXo30/XZiLFe28zyQVpngpE7iqdcL9sk0vPg/7A8dyxAipJQK9xF4VAleEF8ApSgyM
Iuad0Fi/sqQJyxy4uA0tej7FFPnwHTq1NucXmvFiLsFtH10tTPlblBKRreaApCkmKk43wMgJjTB8
g/mnRnUtt3g8wNZTahZy7qFbUlTCy52881FPHXVSAHTJxNGduKdXUptx8HxIwCQmOLcElfTcEm6A
yTJq9W/3DFcWPl0SE6GDwRvVxj+9sNZ2AIIaduBn9gedmOEtgwK5Oowv6Yxa0ofAZeKZ7GpSuxc1
yECY+VUqoC3qdskrVBpcWdj0+azjQmdo/i/Ab6w9yRWp3dqk9ZXTjL8IQFw4258LX5QKEM+MMUBg
rMd45VY4hNxazVF1yB+SA5fob2Yz2htKBCOcneEQIu2OLtKDZbp9GQD9otoHiA6vDzWgZl+31ADB
J46bAjEe6e4eqYbuEvjwEOTG/lJGBt5Udm/OG32tGbtwZOJXVsXpULOB24hy6fPwZ9Te8qtg57Kr
NLdIl0y2t9bha/Ierbyg8nEylEun098tR1lIlyMKTljUPxt2iMfXSfNwVoX55seP9XOd9BZz02EG
qOVkdg9SNWyI1dRQ+2JpKij2f4RyJSJOI2q50djZz54xRfLDp9HjgPs8I1CDvNJTFGRDrSNqamJT
bO8NU6b5fN8kDTKvIIp+GLJlv0ngImutI4dnTuNqRx16rGq1lqcHagz0HhxlI00HLgqHVG3nfOoW
A5WCDLvfBT4nYPhwLtl+4gcE6fxOOkntHD9eOtJ60w05ftVGuPN9xeuRAmFC1sV6AsTitHCfgKPg
8qD7JTeviseMVw/Wz/ebi4CPFxQZvecm+P8/OtiIQySfGHRr/oxroD/9//wzOrKRsftUOlAEEYcs
Mhwtn34zvlGmYj8TOqf/dnK+vokqGDa7OVURRcVtyojAy3g0e27EEDOjwZj1C5Pr7eKrVoJU4mMt
K6U3e8ccdQzy5pDzTFgNkwEmFE9NlsFNjYlrXtF3kdt2/QuZQxBMgEwFsjOnMfyUBxR+PE3vMGcT
xV/OdMa3zWhbQTv9YdN3H3RPHTxEYJJ3TeuaCe05RCD1neoIkmA1q+HTmAtGFtFfYeo+q2t5ZHdR
0S96AIEOBl0v9Q+QRetfINqS6O6iAWmysOat8SbNtT6jEep4FFq9vN93WxJna3crwRB8z73v2ppo
k4BVmamRXggvMRdf2fQVOIE5NS1xaZEqcDzRMMQCpmAwp3dCUxyUKOBAEbwJbSGKF98KLdwYtf90
n2ar+BlNyffkvBJvEKWJnsDgMjvBLjgylZyTgMlpm+MnkLriK683lvlNXMHfYGwFY+qEYk5c8kAX
xQjK84n8IhpH60d3Om+JRG/9GokuyqY4/dz5+IDKZtDDHc/KiINmDJfGtInlj9Cq2FLYd2Z4gLk0
bZL9sqSOKC8ixjHVSmKFMWGZBAhY9n0ZPwx8+ABo8/IPskE/Z+9hqJFFjb5CSby/lb6zJD1NJjAi
JIXtF8vX1PPxvKpEk9QAl4Hi+e4XsRx7nxb7J3CNEBPa9NEHe+C7EpOCZfXLkswhCy1gnb1J8wMu
KBsgfehDT9D50tKa642olcVmKWTYI+K0g5vUa3nc1+qpcGCieB/Vpd12HaynwvwQd5Rm1NUZu6p8
1nUCBYZgSNTrVi5Mw4be1KdZ9QQvyKhAg6X4mZbgBUU38kbEKjlB7TAdr1rb1fb2blc7IjkHEhz5
YGuSbinU8yzeTJ/1aYWbtcvpVEdx/8Cgdsz+KzSJ49gWXdSvrkmJ1bzyWxY6+369KOYiAWooTq8E
cX1/QiRCHpLotBH9PJBJpV5luPBEUOnW8K1fXDlh5IPhMTjfJplShsjT4MauC14rnrakWGiNznIy
OalD0z4bhHoz7TGtK96aMQTozSRuxtLQIu1k3SU0OlWRw2b652awUB0RnsXq9Q2upo0a5eOmUWYn
MIc8Po+xTctRVckSEJN/Z1SlqLIOJ7KzHqQe61ydXRzVQm00IEPOoKetr12QYdr/3+YpK6rbzp3D
2PzrwQTSeAjMMQuZ4aYtXyZpbWsizsCg621PE3yYK9ULiwe0/r2Bttxe5ji6CnJ3pAVXwIaul7L1
TMd1mH4+NcuBRUT2juICKlWOAHihRdHxD7l6aSMqC5xb/VJci62flv3hB0S4PK+xY/hQlvg41hfG
Evry1rt6kulfNMarS/gZlOnzaNhrGe9eEGtoRdQ/S5omlNposct4Ysk4b+9EL9wGmxhWIDjQ8S07
Wa3d4tn9qDhOl5GtBSJgVZUm/bMTujofJmoYPnDfprP4eam4JoVhwycKkNGtwMEyYndOK8I5VInW
3HSf1krSEY3tNfysMMjCDFtYz7TsmpVxQYYtO4gjGpEdCPCGGHTn01vkzRfvQanRLaI465Rp6bQw
4iYuvqRdPtPEIGl6Udrc29qrP4+7KKjNMtDYFEFWSyURy3HLlDUljX0w3JCeQ9yawhrGMA3kE8HM
+eK4v0bTMBBbu38HMBZKOYpqVAvsCciqRDlYeI6EjK2+Xd+TAME3GLFgS5dQLyvSYfT5JcdOln9Y
p3tMkznWklLCd3ovEmqAvMhtYrVGOO9BEw66Led9OH8jkdDdjS1LoHiOnH2xa/Jwbai101p8NpC8
zqsxTrevZuuXXBJRGWyYk/kiHUlI4n4/rh9MXpWTSH5Tn6jwRRF1zicf0cDuET4MMtsbFpDvGEEc
OaXQkN+KHi7WZD+OvDmtGowA84H7R+G4uZpwjbW/EKUHf398owgAC2N1+fADIElS658K/wRi5B/3
D4K8OnfB3C9+zR/SC7ySog4ZzJ5zJ3aLDsF6nMQZX6rkQ+CZsQgOR0oLUalpepZH5FMfaQ3vEzUc
f1OJKmBTctce7qddLCiYe194PZmOItfT7Sujb6PDa49xQsHGcjM2Um1VGNDYj2rxL08UJ9yB6dIP
ub2JXRi7caOkKjUBnKmdb3KOiGJBcq8/dzdLGyz8+eDlaIq1MsRl6D/acNrl3yeGiQ/MtXFFbobL
AKcF14wt7PFSXurNsIUpdK7wOb06zaIbpf65wfWwH9vyqF7/YUoUIsN3fT2KLnW7ySsnWd1mhxyC
cvt/aukOgZB2cyFIqrUvkBKoErLG8DXtFWpKJFpXTnkXp0HHsVcv/OnhSlMta5wsXRfN7Ez7wZw8
vcbpXQ5LcsLSHrenDH2HpdBm3Gb/ag0i+re8NwYx0mtsNNt4rZTCmma1CGuUIpTMPZf2W+LENXyi
lN38MffOvZaovkVEzMJu/nezQkm+y+UGDIn5sjNdXsFUobgDj7mPY7dvWhmk+uYAFAJkJejvK6SO
dSq09UJKun3eDRcQ8YG8tGuOolfBs0orrne8vBn/HK1U+IKpbQUNnLB7VbT7uOQs8bNKgIO/HjLT
BuHD2Iq3mS1Agp0a8k7KHN9pfZtiInO1wkUddYwOvA4qZlhffI3Bjx4H3g3G1dqJO8DFdSCMxsCl
A4+RsX4FRHGLzCGMjLwXrZeBmk6O9heBSIK9i+cIr12+sYp5itPnA5p38FD5WaWuzVFBWof1I/p3
3orF3qWTqzofqiwxEiE9f8TBvbRFXaLdKVnstV0XHvCN9On2ggKpcdLdgELwdyxXp4AD10DWtm24
nrLOkAD0eLWaNR63HNBLBbMPc+p0/DSqcxLbAPj7EK0jz7sb4YYOLuA+XMofYazZ6Y+Sa2ZFsD+0
wJSzNG2N2QmHQ25NDOrVrWFjjGlwKJN+PMGCeDIFc3gzAR4WvjGjL+qs8acliuZDFouh2hbej0O+
fiiv9lkGKoRwPCWf5pHBxuZF47nzo4oWPiQx+W9DFUFQom5A/eqJ9pkBSYartZHgtPYQEOLVFUJQ
kWNSNe6+R1ZN7rfUHHLVsfQDGcvrH57hJHw9UqJHzEgempiAS+MOtEoyNI1dhFnwYJp2L6BN4md9
xos91yem3sdEy+O6tITSQsHto+f/znAIRqzfLLby9t/1jMejad0hwDlkKFfvv8xb7NKr9r0sboZ5
7y3UYFm24sSENkEWkkIQi8n3yCCQQLVI+9JydeQimWkNznIwUr7vrCEZxu00qyBB+4TIt36XY727
ljdRkIE9MxSAHfR+c33giJpLZcd4q+hCdM1QK3cq/H/Nvd+QcQx3kr0GeLUpf64A//HpP95c/BJ4
NtZ3B1m1cIppkaA9dwtTGwwMTQu6mVv+A9bLFySyKi1YKf1+1t8zJZ4BW7GLTI3QuXw/zWKEJ1ZO
ekWIV5A+Z2mWP60BnswcIyFhzZ7WoJp/MM2jMpErkVTRBeneHNtAgBgRIZovc8Fq2OlGALwlBn0t
UC3kdnMdGqok511nrFLWi3lfBtki3erP3VcEMgoQu3673CWYKHOehKDMRS6sudZy6X1KIkdjlq9b
RIr5gJ2vQouMU/InKHYcqGqKO6zssj8NxKdFOJcn9hTHoiFVVYbQZpIWyKQyYoxPIKBC14NOY3v5
0LY1F4SGJ8fJ6ZFryc7Dr/DYyNGpRFeqTgn8OzO/WHoOS0ovw96MIsFK4uiyH03Jo4zCRgNOS4/P
dKy+dJLutZjITzJS5i/SrzKJa5ikRGw+OmuYFsS00VkS5IUwkoofwlBnZFfC66j2zodbITimI/gu
2BkNuhRxyuW2ZTJhAqoyJebmm8AGec48ajL2xS7P7Gb+HS5wFSsV0pj8nBehl7Z8ZkOlA90bcasc
PMKNmMJsw34d9FUUJN/4xsN5bu/e5lJnc1zD6PSuNp6kU7awe81/41hlsTpKxW+o4shNAw2pGXkA
ZeQtP40octVV8EX6K+INBwjbEaNddPkq2OEjXscUf2zxtgyZQwc5L4WiCOn9z89LNwGQOpEiQ7/+
26dFaDLbpBdJ9/scG0DGEKhI4qm351kYNO0+x0toEpsbQWjSvKcO8LkGEgAM+stIf1hB3w5DrU6D
JeZqYgdSN4llWvM2Zq8EOSpnrTA14BdXKDTk8kLo3j1XY509gp7CTfRgXav7DgLFaJQCt8+xe8/j
8jbh18xw3nt3DBmsZM0KOqbIroNGhu51D9e6X8DEn6EDM+V3rOypPwueKCy0ttwsaCEIz6ISkjXJ
n6mA6lmLmpX40X9YmLt75a+iImUj78Q5ZwHLAk4CeS3ugHpxSKvlZhfqggkjpUAC9VQ8Ek99pepF
UeZ2xtrl0wkNlmcK9Fka0AkPZ/CHa7Prliripesn0MEkc63oDunhsre6AURp0+nTIJojo/8Ru8Eg
PZQkn7JCswRw5V4HrQlLNui5jmWYq2zPOORbV6pVMUtxYCz1SwwCyg/fsNx3EUeDFIpCQUDby5CL
HYeVJn2uW1Cm38MTiqjOPoNPyrw5dh9FKlE8eUJtof3Enll9J5CsKklTIMsbcYUQNwEJNDzWiCQ0
o1AgbFNrRfW8O3Np/2XGbNfMIt7kZRJFTHGe1L6mJvtA+Hg0mALuP5DC7MQNWqNPY5N/qNW0/3m2
FZ7m3CWKtwQIqiMMv5bCkvUHpI7OGavAnJoN8lZzJQ4LF8mdoNYoySwz2K2mJr+WfgnYr/T5ADW4
CbU6ZYCwJ9MO5ScP09OuFe2c0qAkq3hzey4kWU1arKUMTPOfc9M7U1WQ21XqEDvpxhe+8jg62ync
/jQc1RRQmo24aaLMnlzNzLw/bc0m8uQJC/9CIw1CvwpED5EFVCvz3hcH1uUVW7SXTqDMpAbIB2XX
gMOt9eQDQ/RY3DgIX6GMZ7RI6eLrbZ6xLKE+8M2EhlRTR79J1EJ0DQz2oOHsaZjiULrfy7DFAKci
4y0aTnNmA3q7ggjawdm987QHBpVMxddh1bL9PvpVyxOBFvlPEu3fQvfkQf11WyBZRbMkqb3u3XVY
GDWU6MYkq8dCSxsqXdr64HQ7kI2BOt5SkSQRhmJa69FQ5xcojNoqTxwAsRdAEFyEXw3zAwUTygAM
GPt5d/F2h/NTsbpcvk9k7UXuGoWFWvxFzVkCTm5Bc2uqtE0nuifVMC8jLXt3gZfz4Y84oIjYYXkm
BFR1c44Udp+TCTW8xnncpDS4mW8xKSYYH4APtQy1/5vUEbBR3t711zdtCfbXmMdyYHykWnTOga9o
lIUCIlPv5XWhA2uixPe1SP69+x9Ymh88VRkQQm+Fjbm2gZxM5Xc8IJgk68eAmr2fVslFyh0ZMjjy
OEcuYtlRyNZvmL5stt8f7TqP9/TLJQzAuAFmKA0USo6f7hHHPaGbz3hQQvln4CT5eDgKNYG3fJDU
OE1oaYPKriO7v/BkggylVoo/ZI9RJNaC0iEKfcapbSo33xRr/qNtkrnxdsjXsCjzSJl8mLEk/oSX
ouJivTJPFCwmzUwvalMEcvHKKkSpBfVPMFeZPy40ctAtsY9WVBEnVgJJUMKEi9AXYPooFasYu29K
TcxQjxFMqOTPu0S03incIgkjM9sspLCeAr7nxo666XjCRqsgX0HjmguDCaklnFSy657yW/UaNxFm
LZpAVS56jGoJBgA5xCNoZ2OHubFjxhpf0Cfmjqi5X7fOtLNKpdt+3crqqWLmwfWBsbrydgKIlC8/
NmZTDj6rJzD+5KZA0hhLriMGQvNv+TNFws0fUqmZSpfyZlNGj084YcM9lI0UU16HSZzqoVWCqv+R
CMaROTaKsu0uDt0HU6PQZoDTCYLAcb94TNkfj4+s/3+wXHNqFlmgjH8Z6yfWVbU8LlpltKR559h7
FpWlu8sCALiLwudwMo2VSfW1ZQlzhQgxoDcN5u+iCotZUOX2OtW7Jh3wH4HvDgo0acigFVkAI6sC
yh3pJaEjHKSmV+pEfjqMnAVvtfHsk7+PcuvnG0Qed0jyha3wcNAbGEw+uSPwjh9Pvz1m6tQ+VWkb
ugkQACjZuf72K+EPZdcrWfBpq3t3qG3iMOc63Ok1e4VkLj++NPFSs6mpODh9sgFoWd1tHUpqOmoS
2IIIjVcLuVKje2p2lpP2RoNFcUDK/K2O5WyqP45FECEs3nW5lIX0CQIMOOp23g84AAdb3roS3TKH
A9pn1BPFPW+Jg4VnIgbEmddr5R/9YN5x7f8hTYtHfPoQmX9TZChAYDbo34GTZEB553RmEgLuBlYj
B/egwF8r3tMvHq3RcMAtm5xv2lT7sHxxnWy0UNYYP6MnkKYxepKS2NeWX0VNlfgYr5VO3tFnpN18
oIyQd+zriqk/8RqgMH6YIIZkA7xkfy6QyElrvBfIDv2BuQtYOkTMsC9E1byDhirP7xA7odeejyft
DPOnYsgR+madUa7mOB1grhVII0NRf+PadnT9tlNw8VMwfirztxue1Wu/z2hrRxYloveeK9O1eTCo
bncQkLZNRAbNkDlKSGlczfv/VKDwYtNUJBaGUySXWT2r18aL+4H50N57O9M1E8YUmTxKd0PQk+HP
9L/lCgmx8AYIUVQaxf2iL75zq4goYlqNhgbxqDgNEtge5nIwHKwFgrRx7wpcwxHEUnbsv0ToE9oW
a0NUbNpIu3jjr+gZ03XQLLRNPbsmnBu7BlDvAKMOkMC74M428NTVyXa5GouVIP1SFAda9CbaEFv7
eAodmbZvGQgbiQHQlVlCP7rOYK4m2g8qkxdiOHFVoBw8JZU+YtDBwMVIk79sBXa3LAdDSkFRilt0
7xs1msOtqnlQ2yLUsK+niZChHxASBtJLtZ1FKEOukeJK43hvonmHGu3iv0LJFtmMTnulL4ikVDpQ
EeVICvDJg2dFikiYyM02pbWEYCzVciflBc/UosQSAUZ95h09Uo/CcCl57VNTVMrdEiJ26Dy/3QFR
Aj7NjdnpXN3RAS6Px66cGCIWeK3WIE8Fc71LRJm4dSRmNSBwHDbFMg/SUl7MPk3osoftl4yF6HPI
e6zJ1gMfDfYEX0wcZ/LMWO+HGtEIBVSRxLqZjxDQdJaD3Ts/ogyFoIWF90kg8XeN9bZW+y7FBe63
W5OGLtCgk+eMVBAUs0S8lPtx/iImIrcKMzSvW6ka8vCGF33uoWoCo7povEWyaj+HF1d2LDUafXMV
X+nA+SXfNmV7aD6g3W+FMnARKRdS/tFdeLR0DN3EMJIlYfu6A8tqfKZj+Vp7rlX9DFQSk6Yi6uKO
qorB8VwOT34rjZysj+z3zY4PoVpOu29x/5Bd3RMWo5Gm3H3i6cNantd4htZPEP3l716PN5vC4kCh
quTeiP2YfTnPf/HJ4saAKrWBXZugqa+WxOqKPvsdSZVC5e9xV4f0acjDU39pnzOdOTbN+rgIgVtg
/coyZBwicSTs/r3x9EpedyKzSOJou8g92BopHsy/3J9+0XFnnEQyFbrhYE934Sqpr2vNlNP4bDfk
+nJtMGP+BiS9YNnP0+77ucRVyGXVThklDBZI775cf+CVSuS+INzWhDuM3JzTuhLBORw7wUWqj9x6
pOnuP5SpGQzY5dXXYpXAL5Zp9q5nyLdma7cCTIp4Ts84R0DqPyCveG4KeMwoznkcGBXuauaO49v+
aR96bFoxgAcOI3Ut2FeH9unsoUwYcNijt9rLrEq/wKrvbEdik6hYV8cZIqpWAis9oFoouSaWFWBt
fNhqhiCzgypQbYOZ20gVZmHgwRtKBd2uyaWdN+8PEJUpGUrzhYlqeM8HgIL8bQDRk+Gk6Ss+QOmi
9DjXHUqR46WUNGIRCswg9TgzfzCZgQoc8TNgtdV4+isfcVrNXe+W5VowEoAou+DS2Ni3dMiEvxb7
/v5fLZrBi9ck9ZeFH0wtA72jaK2oCMlh7mO4Ej6KiMFWI6EWWesZFm63fuDKwzArGq/LXo/2IKIk
ERpfXiEFP0rnB124fQv55a8tRrGhhmQ3CBozwltfznWepYU0zHxoATlz0zgCmGUl8qfLhiBvHdEh
DZgTvl8+hq3B7pEk5zJJ5dI+gingYaLrfio183pIQuYDKt4EkhdnLiSFJcOrji38ZLMMm+bgW4Jl
3EX8D5uFeyDEtA==
`protect end_protected
