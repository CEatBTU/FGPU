`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nZFDDAe5ykc1YbvYlUYKcF952AWHnVyt8JMRcrxrpPcjcm+fiBMlhGHOfkWuExbOj/6VZMAMnUzZ
2eHYW6nFzA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YWIO/0NN1TJmWrriZROZgokhi09TbImOOa2P8+vvGd4NJ+fzBqqleDWtEk3JFhUxDGb6mrmvNIPQ
YG6gXZheNnHTdJdbVS+xEF9Gn/ZU5Z2GaoANBUFNjTb3d9v70B8VeRA4lWu1hNLZJrINl2RUV2jM
zAKt6BTAoXaltKesRuE=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rE+Rvq9lUxgaZdcpB64TBRjsnxXemCwmW1k2Qh6YjVFSsv/TlBQopNwnfv5tP5OMEs3uajU3WKBp
zy23QAyoyw53yG0kCCIcf+IlXkiRT/SY52hQ7TM1StD1FPAUOB0DL1FJaeIRkJ5yRpARfZbFjzHO
DXQn5yxt3fuWLEGSbs8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D/p768Ql+sSTJiSSuYW2JDK0yViOs3rplUBa+F9a6vI7wNSlJeyGRgmOjuZnotw17jwlRomg4/rN
soT3PfX7Ufw4RMkve6YUeEesuUi47KlZNN4Z1vV3QrgeDS4cVJJsAdur1hZEZH3y3081skVnAYYM
7tkyc3pSbUf/KHY4ybMCHRqlIys0BRP84UvAO5ks+aq7t/+FrZ0/liPzYKpzYcc21nHiFe8iTokZ
zr2tecMFjJdLu0bcQcwD46xsUvJUF7gi5YCLqKQwJCHESvHxWluHtNJCv76xTe1EH0ntNPaxO+zb
NN5Gv5ao9JylzvxAxMoPJf6lOUcM5V9m3CF2Lg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b7sUV6Dck7TsdyOJMVWqUGsvn/XYPAoTcwEGKw59gLUb+WixEkb9U8qVOe2+hewp8JL8MZdr9CqK
o74xGNE+VUM4kY8VqRpgTUGRym/zjew3A8RjWqknbZPAL+fRykH8zojuGjtMQm7iV1TpWEdnn3fq
ML6qFNsu43CyvVkqLTPcPeutHA+HKRndQagpEDgXP5UW+NfjMGx+0gp7tJrV+TD/qZq9BNbfj1GR
PDRxQs82DULS2Jas8qyFImEdp8J8tIFbVKtTsquQU55npmmlc55sypXhy1VQiLXNKEh5D4JoJPeY
7RhvTb7nAkR9gCfNCelQoYHnr7vnYVG33yCj+A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IoLBGa60diGteGKdysc5ywMV9aKpkNfa58Xce9+6i6yRWyFL4HrkUqNeIx5WAEL2tg48ckJKvO89
u/L4g34j7ImJLUVrpSjfoj1kk0GHQo7FaMcKjlwes5sV9qdmGbn4ZMUzjn0z+KTCnppE0vna87OG
/JpyoVZsE8R6OLB1WM+jSagGtbwZ+04fFewAQzGOri34K8O1oQxl6cExNqXmKBajEDotRbNgUDqI
g02DlIAdjlkzvhDp1nxo8rHkBiX5qtG50QJNfgmUL3ibAP46naDOGMiTeAGyWB+3/IrzhGLXldRl
toEAoRgfXcGKCcmoHYxjOya5r5GP8TNjP7YmHA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57632)
`protect data_block
Eep/uSlu8QI1KOuYiv00tyN2jGvK/R1q5FLvHS2QdU8JOILzzp5H658/yBgUR0H7EUiYasNzFO69
gG/NzNlDI5rponkts0b509f9f5Crw7kq8EwpbnV1gAgfCYstc6WhpLdaUXYI/yW/t5Qzs0oaRjIs
sx3qsnaP5wlSDcytMnO0LR77gt1LZYNv30mdG3IHuoIZqvFZONRddg87PNKu68Y6MPwBM2PstOnA
kJOAeu4a7Q4k9mW7+Gafh7+E787qIlK0FlVKzjjghnFgDp4BucFIOEh+pW8YtSTcqEZwUbu1YCwA
+ifqIXSQgxRZS5Tu2hToa0WASH6zcxCBLENAG0e57HDj8LJ8aXh3BQYUiaTRwN+J1t6auZq+lhCF
a8pKYUA3g9qqsQa3m/Shdl+ijpTnvmB41Vkpnvxmil8JTMY/mpypGSlBQTlB4+HzLm9aMDCuEB80
vjNbGj1L/u33kjKj9L0G+4TLuYYyNiIIa+d1kyncmZriu2t395jGDQcwEIfhSca8leek6CpBgPKE
g/WABRgUf1CJ977sCZU6xJfCrIM+rFE8sh0RuF9ymUDlDloC4XWT18IQk74fjmfc6A+PxhQ/+io9
3MNpj4TvAAgXyxENmyCQZdl8M1o6AbGwqH+jXLW76TuNIJ9Iyv4oKKxBpxV2eJ9X3FHd3WrfNT5a
r1cwTg/7zWByUvCPanyx2wU0EBhM1KB/3tuFRuD58V6i/owEcMeYUdWHAilmt4o9Tuu3gtZopxpY
bc7cVeeAcZ5fEKDoVKq1yWCJhExMMo/MZiz9TSIYbjcafVegbV+/mbJI0Ev7beSA8Ofcse58odrm
DlaN5EG60a3LxLsENtNTEJo39vNIwQDaNgsvmYUJWgtd3Xoj8e2DiLAUodc3f0PeXWCHUILvMfnm
0WLuw4L972vNTLfIkLOvc1H5rSHkg2jUYlue4Fu3lRIvwpwHDeOM2nsLeAmMFk9l1pGdTnMzfgWy
upcDKN+w4F9qLt0HHlGoel8oZ2MfpVvU0yN5SUuap9veX12D57bpx1wCZM1kChc3QapYj2UqJxOD
Q0wF/mpDtXZZ8oze7aMSEMq6UGZEZzb1P+dd089f7x4WIh3iTAfQSdaetDVWi/VMwZn+ht3uLkGl
8CN0TI+CgbkCNSSLo+zERV4ouqNgTyht+udJ8GlRUIj4uXKNipYHv8UW+LiqqOrXjRBr18YXurOi
bQEZLw3R/HK2vgSGuJD/GEAidaVgQqMRdB6dP7qPD4mTgSVoBzDV+Q1nGbeOX3CSlucEaeCjCNSp
shk8r67D0LfYJInESL2qouIszYwmJLNQMZquo8SZ7dQz5NHDecyHSYFJVB8HiAX59koZNYKTENQY
1i7Mg/AQPCWxiuoX1Q7AmJfbP7WmF9yNsoD0dGtQKetBLL0fgpHNqmsN3NVBFN94oAbevZU9SpMn
DHpqtYE7BtuozRs+o6zT0TdBlnUM9YQ3McvNbJtNCG1bLuXlzv1hO3w+tj8SsTxB29XM7Tm+DXEL
IzqnGP0fCxCgTRhwwHUAEV9H3/kFJ9kQwRID7jm4Ty4+HlvhoayBu/77ssYMtbFoKYlsyksYhWSY
vCLmmcgLxr3mAKmgXXLSYbiIdD5jwAgsNVQkNaH+gtebGoMJTMMfF4N1TSLNpxYYIIeELcPeEQ3k
PFfpxoVsr75IGIb8Bba900Qs0zwRbaSVzZP1W+qzP8NNvspm074OSpPc/oSiSfV3xrwYvuz4R1VF
HLcKnDQbL/d7+I0yO58PAAkpbjEIeiOBkRqov9bfiRGbDCXvl0XRlMSQ2Ra2GTTuKUcge1RSnX0X
6fmolxrgH94K+0B7uQdwjbB08+CFjIhwMSD/FUZMFHHALGIxJYQhbhqGgZyUP/g2hiXHyLP2MZSh
iBVMj/msECofNfqTxHUgTLX+01+Cu7/MoyQNEa19/h7oVft5vZRsA39LslZ6jpvTArIPEviqb5Ra
HZhsvdm0tYeaBhg8JlmKrg5EmNxHqCW1wATp71acfKQe8sJRg5CAUnNT5XEYbg98iROk4GfmLAKk
qsqSHXva1ksmugRdL7aGyewxrdmwEJw8S32CIMzSh4RUhQfolZqA1HD4FWtus0C4TYmqkrv7yr5Q
4fN/OJ4S+fn8/UFjRWKWiLuicruNGWO7aTDfzbB+mk9KaOmQQzRVHgzK62f250YrjBXS2CHZmsfQ
VYOj14bIpt2eqhd937E8gQf71vzvo2lUx+e6Y+pw4s8dI0hUzZhgUyTDWuxp5yWLOob3cQ+S0qJN
XFkrr6lpr9eEC/LAg4iC5TgKjPnnBWxt8iSOx74AqlqQK2T03wOF+7vcXSuXwPol+QC/1NqhC1bK
4c/6kNxLAseSTMIaO4P5FnsTrGZtKZwobIYrgakrdN2cS7r7ZtPjGsnSAS+/GIM0j37RGhPQgNfE
8fUi+fn189XVSZIyTcL/ywqMmtu18KVw4h5VogvbnFN4BG7xF2p8wYEWc5fT1jvVYGXHM5hOmS1a
lMlJ1XTFhnMUC0yBMCH1l2Sgdk6H7XzW6jaQhTc9Ng8PkL0bE310w92VsjC4uarDQa46au2XcJir
IHLxcOXF3buiGJnrHZVoSaovhmUtun/kA+4yFNRozLaAwBQVC2T00xv/H5ZUQPPSqLmXCfVWNTj9
N1j0LeQ2Z7m1Uy6eIMivU2GL0nVfA7fshZOOkIPv4MdG0FW6ixqBhURo2TCHT2V1QoRniSiT30gG
6kNm3ze48tAcEay1ucGB/nsM2L63poFtKCqDKTVzCnTqCLOCRYDzM4i8GQa3TqmtM15ziUzsYXCw
rq3VZ5ZqXMaAWkxeHbNOaMlZUsD5N8uMatKagNM0xlm+SWkRmowrDg6R8plgDQ6UZexEk/HptsvJ
H4R6gbS0Dypv99sg4d4KiUHg1MhbDyfpCrixIBIAAnyS9tyUIqfSAK/2/MQCMIaDO7R0n9w0TPam
VXexU4FbZ9NiRYbW0zbSRdh6aE80FnTI7N0n3idTQ8pb4V6ezwAuaRlFyQHCASlCD4IbDl/sncrc
cvO5+t4E/G8WXZe520GS3JQdwoz8FGilK27zq5cT0+p7v5hT+wkfYXOdP1oiiJJ9T73NyqdVrqod
zxVISHZeX4h+hGCf0f63gLdW9NHhW0WA6djYT58UrSOwH1TQz2f+d7/8WBOveRfuAFT6Mvs68xJW
+ebaJ3qJm2qb9FjO/QhWiK01cZphMgnPHf3BzavJuVnc+XI/bFSj7GnPpajLkIZEK6gbBQHkxFtM
OgNXl+5A5XqU/ycRVNVC4IwEndxL1N/Yh1KBMAT2h6QcKgPkboH7ZF26JlksHU+pE6vieuUB1o+M
3A+q8rnsPwM3om5OXVxwCYCZjAp4UtRQQyU7RDFQ97AX7RTaMtmoCO1JqhqtSK4v9xf2rDQ6eGEY
ydPGwTcym6+Vq/YutQdDgFUOU+iE0TD/M376Sk/cnvNwVoyidFTY/XHwWBwuhLickg2TnZnqFiUM
1WLTjpqTwheC2ZlKweuuPh+wPkRiq16H0KcLKldT8CzLY/H+4nxu0yyMWIZFMwQwb35tIfrargzH
VFz85mRrCDum0UBgFedLvRe5P0zvi52UFNE96DFjXje5Q5nQR2PlEN5aFAcTb+GnLwWTide3n3H6
V1d6b2sqsDWuBm1hOe9iWdWHUv2FMEKQgfkVqxAbVmFyNvw+0Nn0h537HyADF503GBnlgpC9uTDO
XPJF7suXyGAC7uGLA9/lpA29QqZldUZwWnJK1CskdjcvZTAMbHSQhD0eGCoR+68p9+cgCZwvp/Ss
CXdIHpSkIarJBA+koXvDsjKfZtUtiBWGfP/L99tvjfGLk1fEX9jguu7wli8teAZroaBi/refyFSk
7KRcB73uFsMFIIiSQGb+coS/2iYCs5hkM6AId/S+NC49GI5cezpvsudSiXeFJZeA14tNpkAQk01u
0ShhDGjgLtQGejWTwcqPnP8knY37F+d6bstzqXluVgDTXPWKVpgqMdcRz57JJf1Tv8o8QavfUccC
oxUJX1CKY1kiTZrYr0ReG5WTHW2EENEzcI1YXjzaP8Hy9Oq7A83Hx8ryD9h3pMequcS4PFtlNB/g
iAQAJtntsbbMERc+lEYBv9p3GwFFvYTkDjHR/Do+FcG+1awWmk0as0kV01rkDtiSGBu0rZGAaEFu
D7tTbbomf13qUUCKDO95o2mE3+bKZjPpMiqvUi/nW1s/pb/GycCP+snFn9xrS3YkfP40vSrtrqt9
g3hXoAdfI/4WK/GIs+ZtlFJ6GY33+CLMmIUtgXOeTQAr1kDuQxzB4QF9NwMOSlKVmg5FJRxS9HzD
tHSdjQlxa4vAguelbi9XGQv5SV7fda1vUX39uzitbzPQ4EiQhU2ksi6RXliyoudQwxkkJRAIahqY
v//tizffNeKuA76cIg4Jeb/on9pASAJvQJrBDy3airyYOXJNHbW8em+frPnfzZ5Z5hU+w1Xllt5F
ICtx2cUkuKsZ0vqUyeXHsqWyMwyQeEq6lioqu80QNCsbS5HzdOs8UX0khPWuU+siSQDPN7a+rHSL
Nobrh/4GmDZWI2Fvo2rLAM3RFxAVb75t81UulM29uZ4TxRlhhxVfA3kuEebZtIdINPVJuqB0VFe0
C6NUDor5+eJnSJQi64UKHtioS5uJ6xAQLdIRE4KGEYZzfz3DtrDDkmTGr/BgilGlnhyRF2GbP6B+
HP5GYveflkpZKtx+59fXH84RL2DfZ2Ogb83KlsHkWoWJEgIjpl2csCNpjCqbMTJFfSjGwpt/agIA
qNaiNJjpwWyr1b9CSuxxZDHXYVmmtevDeySVur+Oz3VBxXvt12TmV5gkfrvJf3hNeik6gtBiIjVt
2JfniICF2AVLX9Una4dOdBBBRG+Xc258t966baE7sUkXh3M5LsEa0184gekp/V2qo6TuQSIK+m+9
Iy7uJq32az1oFwHOOK1yCIo1Zn+9hjG2erkKoY007eAO7nktrr8OwFtiei/tfPLUKWyyBSGeAywm
MFd7gztUWnBERbdd6eUO2XRpSjeDta8jO1QhyEJKOcjNT57smfUsKVTQ/UB0++ZZCrfBKkjR9TIk
mDzXKz77KwXTC0osQMkGQJAxlyODF4TTj62d5nnKUNtpAXYaRstiFF50uQMUyoRwQq3dHp5DnfeV
lHAmnnoh2cRC3o0TxCboF+nN9ynOjgOdxpSzdoQCg8nLVirR9cyMZXf1h/wOWw2OC5d2e+7vlgEm
qvY/ZjsVvfBCwDYBnxnFoUHMIobVImyb+X1qpSDZAJPpgYE3o2bMGxkHSCInbZjvFuagaWPMW7Rf
wu+FlBcyhDxjN4IHnLAxetBea86/9ZK7ZmG0pbnZvEW1Ay8xwvhWNDHvhobCwbWJJpd99bTEFegg
yiUfR71zr3Yk5wPIUcW3yvd/MuIyMNgM8HvIzXWBGnXA0nDK5NQDUN1L4xz9inPoyMt1W33XOhFH
27SUVwQLBiV8g1Iaw287vv10kfdkglY4ry7j2ez25pUyi6H8bvciR2Vyejr0Do7yH0vLYUgEH+Lj
rn0u6+8EkPcYBorW1+tJ2kdVkaklpnM7Va/t4L5Lj3jdrq6wfT3SPSU96tY5M7bkQiHji1Ioz8I/
1T98XVkHgIhBY0HNoGlLuScPt6dlUOWBHCRJ8BTFl002yKDo3Rvd6R6TH/04Q1BWU2waVsRPDFTO
LzXjdz1Nm4BTR/bUBSiLGfSskkB772ylIhbQSMLVeUfkdJiiCX8IIqfbdfyo6HBti3RWtAw7dzI5
ZBvIUBiOH18QLGgA2tOU/Dao+C9pVlwHgPDBRyuCnIhnuYoBEqhMw4sMiVaqTjeW8L08IedqmXgW
AGUKzn/DhoF0D/mJFeDnq8lYNTId3UnaQlQKhzRLG0KZTn3S2zvL23ZYTXhPA44lwUdei5jJDctk
t3PofTF1TtoSEcSq6YHavtwyvIUoROmoq1ChJpTqEhqtlajdAEQBMleBntMOACWI14jgPiPteiSm
lg56fpU32oYxWIBkyon72jxRuW8SMNwAyQ4fwLCt8laSi3snC8xsV6SnTrqA10FqFSkpkmaXbzef
Qg+1cUlo+plbRyam4+a9TloYcEceWPfDd50pU3qNMYjqdyasGvdne96N13TSFloSaeJZmfQXCPSA
7y9bTr8y6Rwm7GOsIHny7GHuBNkh7P1hFvZXhWcfLQd4DdoEMYVTisL3ec7uHFAvK8RKGKGdqXgf
VnoygNSDFybkS9jyOpS+lQIoUFF1ZHnD3LUTpgfwkNxmTO/f0wQfcKgJ5oc3DSibFAlzfURCHi4E
iKqp7oDTGA6PBJFMvTosqgnB7vrLFa/4jY5lRWdShYNeRxGkRW3cfKQgJIISjPAB5r9lLe9Txt3E
4CBls7WJYmTJGT+wZ92Z+Jt6c0LnXfuxq54C5ieJFNyEXhu6+WXD2oRZVWGFyhnHCno475V6F/Jo
oQdGnUZdr2Y4DtTlY9lPL+xFz2KEFE/ma+C95dlsxzKoxE0PbS+ASIhsu78Jj/7FpF+9WepgOpTc
jPD+HTvcB5PMaZHDirnDkgvNIrTURD7KeNowHd4THiRs9slVsnO7/LoDPN0ZtgmnDrWrl40zOAvs
5NDrfxgbDmMsturaTrget2Q9XHDuOHr6ZQRXjbmSEUfZImE36nnfB0Y1pvyMsF3MI3olvu5VnMaZ
uza/iHQYhcf0T/rMCZu7bHcCadjvnMcBz41KOXxlezUdGzN61qhopt8SF8wo00I/T+qEZ1ya8HsY
tdm3ZBU6hPuqWXp6H24WgNHQKPXnhbBQ8ysP3dWeTvN/qn/0kVhN2J8EPTAPd5iYr7F9B0sivZMI
vKLDIPJ5Yv9LHp7UlEXU98f0CbF7nvcu26VA+N37UiXXQK5LuAvHWXg63sGAq/8K4ceNtnMlZFTh
KYXHEvMwd0WEO6kYtoqR+vJg/5mgqD8jAYfXdpfxEGZqbQubGOCerhLdBpGLOGy+Lysy8oaddDM8
hE/0864dJOzI85mRj20A1RD/JthysXk0auPRl5cuuGuqSmEPeRVGgKN8UAvBPpdXVLYVsiaH1lAd
OuSHbe0uRvrsL/Y2P3kzwv3qCOJihnTM8HzBhrK1GE50UL3pqTloYcRpFOvUiS9J5Ojc29175CEM
bdp5y1X1/bx4AEkGJf+uV2STD9mDPHMyCTZZb4LAFHOqbZmTMCOXKQXNwGqWulry45oivKG8yzON
UKm1f+/agVB62pjeNZeooFrksesp78XZhLNuQGcbjkVyPUrsKLJZcxyQuyZ+ML59mzqoqXgHDHOo
NK1Ker9j9PWXvxlZBzQqlWeUSbK8j0wyddx9CjceBTKhqia+lc3wZPe+v8YkyObrGuuSj/di6zw5
jr1ockZV8/mcdr1y1CC/R8Y76CieabvNTdI9tsbr7Vy35XYSLnyLpzVeow9+g/nxxWzSGFpZT49t
OmCvnSBFIHHUhyB3cXfFtmaBWucpwAvAeGwz72lttFN8Mh9iiQjYzQQLN5jrY08ILFQ+0k3A+cF+
N2trMRNzplbBW0a6MArpZ6+FI2ZTMb681Xmd0y4p4MzXssWroiQ0ERYHwqpKbSF8CIoQ9TvPILkp
FkV+aJceKjnV5nTVDHRJeNER4pT0fA0J5I1b2C0x0Hh1DiKdSXTY2/VxAKKlSwhHQGbn2jupzS8+
RncBdLF6ccLx2T+7V928phG49hTX9puo5uiWzR7GMKdLc2s6gYsfS1pOAfGdRjVacgKbE8GG7890
U72/IFcbKCt+ZXxAeQZL/LlISS/N6I5eYaKVeYy2rVTfrsuE/oFy9bcXbpud0N1knCpUU823NJ2b
5ZrmgZCSQ+m17XyjY9DS3bdm2eu7pvA2Gv3DrCaq9E8qVEa3217T4AmcXcRmqkoTpMx4sfWC71xh
WnH5fOqh39nhfM+e5sphZo/jXiGDgDSkAUeuTnBnOfga2dqNj9PFsDVnUG7S8xOsmXN/bvAmBlB7
biGEcHSANofDOKysL9Umpi2kwNL7pZ0bzcFC8PQuhyTD8e/PW1H1WIbqHGTgti9+2ftdtxSiICrx
0cqA/G5MPCY9d5jmi7g6XwWGAEe6i7LeAvXf/G4R4zV5g8rfUEPaQQ7NSglHWvlWm5aEm6QBtUa0
MwvTo+GxCvgpECP0Eok1HXGMnz7EhdGQZuFo5ZN1YWNawUuQDRTAjwGSgbP4jEIQtLNZQMhD7PGx
qCD/M6nUM4bdHN66kUzV1oBiFMx8wnfGwFxy0MQwT6+3kkvrc60vUsPbOc55m+VMhblLApVL7ik8
R9sG3vN731vyikBetuTWbo0Nr7DFVyauXxKB3LADul04CjTL9lott+6IjJ6gDrbUDD4QkPgGzzcE
/0g/nJVFur5cCH3pPRdeVu9geuZCoaFf37GnQUtgC6ZSAA+4XiC+Y+/F5TWKBt1wBH5obDFwL70W
7OlwRrvSGVNYTkLhMKH+c3wnclCsR2WChl9Z2BwAyCUXYb5ShoCFLM/cw8USXI8hptT2t3Z1td1H
q+0X50/j5h3nOa93xzeMYKfql2hqZ6XlFFP2QFDxDKsS5L2omwwJVg3aOdjN4D1D9XogkZHvLiIM
VJpseiduoY8c+AzUAYtITolQZu0SqKwl2H86RwZs+HQAgut+K/rQ7eC+stGh30TVnCRgkOiPmHTv
gI1mKJpF6u8i9NA5bhfXmxM9dKgbJNHC0Sz8p7Z5Hp4c6U/2jD3XxU9z8wL3MpMZCfj9ODomW0CV
LcfCJT+WX658DZHbUsOkqML3t6H8xDkANuB8/9P+3mZxmemJb5cH+/s5uiLEo1Q4Ij5EprQt27cy
yO8o1e0jTfqdFwfiEin3vA8QIwnj1tJkwOlWce2huM6+b8H6qsUtQdrC6lW1jE0ORlhF9h7bsgVr
pCB1BaBTxXCN+yOIQxMTgCn+60drH702oKb8u8n58fjGEu243o7Di0/QN+zftDMjbUgWdq06FRaw
6L3WnsQi1u8pd0kb6YJ0RLsUKuKNDR3hUFa6hJxlnPx39mjzeEJ7VDhCcurBOgEqpOLC4pX2u/qz
M5Sr0ka0gos4LDyyxqSvYjAAEUQC37Rk7pc5vjN3JaUuCvgG0nsswHWaz/lS2ZgrPF6Yg7bf7t2a
uKqWjw5GwDJ9HR3V5lTv+VVaTiMEqeTP2H3/qeWKWWaNU5WZhRUx7Emk3PoSqwgSfujBJBJU92IG
dyJLWL0QrWEISV/gkvIdTUlFunesfTYilAmoOwXyTgFXhHCuN6eKNQkugR8/4U8cKVdLPSxkqwdG
wI0wFJVGt2+vwdCN/2Lt/wl3NgErL/d27gwDDWooj6RNHLPFUMxhGbvIYO0MNwMELQKeYpuS0yvI
jhMA8LL49tGsjZ+xxggKYUHUYshgsAJmUoTUnRCrN7BJUZQu0buGwnQfADMrLWqb+a7l+IxlwNJQ
4fzfqoqeGX80DVRMJ+EJluU+WUN3laqxC3Kxf2tlnqCp7YyGW7G/bK/BY4VCQYxMjz7CZaup4PjM
JwnypJaOhZnb9PYySSBG42v1alxF8MQxbshS+GcOjFO6tMHkTddML6U5lQC1EMHXRENFqhG2eubJ
o01J6hV1ORJl6rXXjzOGfzcZggXuesXoL0xSpmm4jmy/od/bPtQThZgZbcRaM0DAc7Tv1JJc2+XG
5uoFo7y+Auck6u00sdjKEPiZezIGcGQPSvH2L7vOc0fVm4+mtbpLPBF/jvdzOfhHavwqgFWbxblH
04QsHmMKH2HbLKH/Ci7iwD3csDgyrCiX06Mli9qbEiWYprZQnDvhwhGZTKqMS5/RPHmH5WrhtXAU
5aEbEdUiSdL5Q/D5d/TDL237k2JSZJ+b8kCJNmBAVeX6DLRgo/teT7elxd9T4QEyK7VQXlcMo47w
5cc7QG8UJgK6KYKC2kJYCEgomeJZFAdFL61l4g9s1QEMk+rz2CAHgI9buiqMVM7epOgPM11+4aOa
IcJv6lflC5fd4Lwb2eJ+s+aUweaiPHgzvvUzjsdkDnTESTSd8Ds2wgd0GmTcLURxsxk+LSKrJHwb
iF4nnOYqj5R/AfiC2V93XhSgGEpLHlLYBMoN1N3UEmHdXPUtmM/WE++2r1lvmPKd256yZoGNxYK3
/Si4DmpQJYNGW5XrW6eQKZwrIoisJssy9LGy4nWfpfUvpaRlxyep+kKBpGCSWm/5vx2YY6J/Ax29
aH3dv2KeaY34qYwKXvebAPYWnpVlaQlOgXlbmM3Ne3hviqkvOSDGVXc3AjsZQP9iSZh1KQj7XDQr
td04JUcaA5jVOpvAOuE3BSyPfq3jXjn6LCohlrDLxUbIlUNCgo1GgmHQ0X5xBCrhnttmiC/QtnXx
e+bcu5h4vGB0x9P705a0XWZi5Nb7jgmTQfgMR9qMPIIMyIuXwr88GPgA3n3s+/VTt3erJFqV2zvr
GmUvLnweEi29L5qFOTfRcQufqIDzunm6dsdrOXq++O0hAXCFn6HIWb72IOfAm4qgAV7pl3zDy3ea
+beCOjn8gM96m31MqoF75AuSGMVo13ai+7z+V3ZCZVv1O+2Vao7vmU8/KH4j9G/xmVb0QAq0BnPJ
KZm757pAi/z65W2JOU/AVwTX8qJ45R/+x/HzlCY/SA6fHojjvknZveKgVJWfdxSSgGfFNc1V2dad
snxtwF9/AKbuMxXXYWAAer18EdOEXibgnCLta7deutwX+1+9iCyYKr90uf+Nk8daJagxsGFuEUQz
b+MgVw6teb8+P7GHzJ0F346AQOIPuUritThJLfvk9fR28sYmeY5GE2ihvUbZwzvCpJpvZcY/dgmH
+u0kH/fKrnMhpoadvOoHfcgqn1MO4T5D4Rq0FqwVfRiZZakPLCSmekRBko8F1Ep514sojny2AhqE
1nt6HoVLqJxw4l9FxZ+f/bGXfNHjodJxKdZVTFWcrQq6dn5Eauk3ZL/TkgLfJnXGOnBOYTVqjfWX
LbX90ZrxEHP8z1UjmVzMN2EHwFils2bdgAxtJgMMvikeF3EbdPBHwqOZ5C2dnJ+nQnJzWmW/O3mr
/oQtdlr7lpL2pT3Cm/qDXVaGLlYmxtpFdLHy87xEQ07JGtTBxz7TBJA4dh6a9RSc/RQCcesQ6RwS
mrRTbu5e3gFie6HkCGq6fSeEyJ06m1wTolcp9Mlrw/CYphHYnZxyEa7ZncZG9c0llC49w6cpoi+N
TbHSvkxuQI46+SK0fJT/NysANkdtp2ooekvLVPNvueumVbP4FnJM6eFRGNrqL8Nsc7w6uXK5/vBm
0/1QQEXabtJurLI3r2y9U2Xs4HQMQw7By1CIB10j2AMTLDerU6hzQ2sPDMpSleWhCbIY50b4m02N
wwPi/r+LWuqeaPCZIOmPu0/dRPayAAWWYb4FxA8dv8IgGyfwoaFju55tWeksD8qmBCEZaEIOReQG
kYUyKrm8ghjHqF8DxivjUQtJjK6rgJwzRzA+eIAgA7QhwHRJSwtRwCvaekow8DpVdvFMhOanuvzO
iJ0VgG44lnJ5tZQKCTuGUXgoS7guCpNXLcQFnjAau/Hoq4MsGvcoKOWhqtecepH+aSSYu7U7Cf/9
z1G5kpdiDCbMWAylNiBhV8Qc12wWMsr4x82XAy4AN2VznAwpMyOfNNptY7iFas78V7wJzaFwDF08
rvW/hy/HUP4RawhS1E64D5vymfJahQLy7QGjDv895u9Kgt7nQtUtESblfDORtrWSyVFRdAcqrm72
NOviBArHgsdj3Fk2bINjl7wZ+BH67ktT+8D0ud7atDBWWswDvSX1hcqfMvLPwHa2TAjUlp3hs2tK
R6W5ML1hRv1dJYidRY1dDYSgsInaQcis26wM0LqK8siIqG6qB3fXDuO2ncv0V4EQnJhxq6XrO0gc
NodyOSkNOanmVZqr+Ngu7fqcOFxy6C8l+6KdRUb8CZy3Lk99vDxKV6aEz0kbRoeG8pc5aWYC9c/+
eV5GcENwu7aC5MtaoH0QCLKVG8d1Z1Roe/ji/dbQD7lkAOaQT0NdhsoritcWN3I7dp/GcJUHfXBO
9QFAVFbk98Lw9Nt3fJvdB3Et2XsoVee+wvXAavEoQpB3yz0N83PUaGHfMF/2wk7DIsXeDdRWj/0d
QQ2FauBd9mxf+RIORhD6M0mlDf3F77qOYpu0RsfCviTgKqlcsNZpSJovoRy3gnFJrYXxil5dzAD/
GK3QujYNd1nqwdOfq2HGzytkakXnQJ8ep1HlYUeuFHBwp7Xpxts9JInMlSy4/bJOqtZ2nAH2nPQY
C1DrL7kFLbw1yhScNVg/P5oi+fwnLsD8dyvWrhI+hII4NHXuWJXZVeOZMAhd/Yv5G2kld40QBgoV
3FOn0XAYBSsLZWXUWBTucuN1fko6eXYgoNSWERFibEVjLyPAodmul5OtsYV5x+bNXkizojCOjOJH
u5BZjnG6giirg2Y92tihaGU36MH7egzBkTqREYlqJgaNXnOamkSXiiTBl4pZiiCgjAI1n0AxUekL
UUgP/KJW2GTdJ7VLUdzQ6IleQurSP/+1N24K+eUilk/hLvsYM5Msz1pN3UgglRKH8O9Yvp8N1aRs
Cew0Wpe5QEAQRL5LdxJsWaptyyZjQrLRkOESpmVT2XsfVdO7oR40kFqIDYcJJpE8EwsWNGFR9Xd5
hHVmKjF12pTN/zcdTsYNyxoIlzcQ3/cVYxZuHtZ31KII6vs/xUtnR+xD6WniKTE5l5uvD5Ni5d5V
OBh5R/pO3zIK3V/3/GNbFviQBfswxYD2pT/hy8ame6NPgn+shLnVxDUCwrUVeSLiSsO+TY7b7bAs
O829zZwAsHVsjSCz/x17utR2Hn2TRL80JPg19BMPKgd9K20rjScRzZKNdgO5ZPYk6dqGpLIvstT3
Cq/njdut9jfMZZFXRdVQye/Fi7FZZihsu1axEGNBfsTsAaJKWCW2QD5qxGOPHMt1MiVrWBwqj0hb
XXD215acrzCcTxBIf/eeJcmQbI+p0awofd+VVVP1IZpzX24bUz1FrDip/e6/OP2lWhAhGL4D8KZN
BLjqoqoPRCJAb53WOcAy+L6qPmjASorDSpgyG4Ifct4Ffv8MXFCji7aa8hSGuR4hU3S8Idr2RxXc
N4N1hquQqgSG7gXnDl50o4DLz1tjG/rUgHFp6DVN3opFS9jv82Ou4ZLWFVuRHwO7B3qbK6PO0fsN
ImGTRZJBVda37p96wwmNyuc88wrU+s8Ri2KEghxrA0MyZLgwyS0NJ6R44b8Ae8xmDCX4meY9CI6U
WTCv4QhdPIiAhI4OZ8JlavWv4UOXXhOUfPrP3PTmjzQjJ6N/onQ+Y+GxcVmB1qy6gDgTekyD+o7l
87Go5TAXXlcZELBjCTizEHkl6Jl0dmVmCkbTkexEXhYoVLGjlf9yyg3nCv5qu5/OkrNggKeSXji3
rdsXL+7XuOtg52xHMFqjMamj7DBHDlMsiqF7LhRVE3TbrAo5E+vAAiTUxz169StMiBe9xY8Kd//V
pv+XRRPxVB6ubAIlnmtX+tM9lrDe4qvSlf9EdlR/Roy3F+jWSCf+egdhHlP4oAenhAAeFNx36fSr
qOIs0H5SENnxxVbV0AHRm3vdQcQCbbQlJHC8TSYksH2PLaGzxjk0VswwNfK6SwUfsBc7RGatwnOS
6sfDQJ0MX41JU3FcbPiTs+j0gUnXiOo/LW063T/dTXMyLUVjHkvIbNkXVaUoUbw4T5PO1oiMD8vA
0SFWiIGe4RgDXwxHFBd2w6TdB5wunDdH5AMdhMpH6rXoZ6YsD282e50+Upan2S8+8/3BtG6rtKSo
mXL5yV8rQyjKqoDH/9ARQpzAxnS2wx6GpfMsGdvYTBTYHR92W5JntYDJKk5BYD6qblXmlvcSwSAM
XMGC4fBDta/7KMr80mfL3XwDq6tXUVXMF/M8j3uyZjn3YGWjLgvRtnFSkQ7QOwpLhtxTtGwl66iP
HtcgxlDVYwoDOgi6tImykfRpxIzahRzD8U2cRw11x/MDyzDR5d9yjTiOrDRnOyzuCQbVPahcqZ41
l1bowu+Zp9h/XhngRfSQC7yJ6sa2+9PcEQ0iQzpa7VQyU9gr2WfWahEjlvezp2GU3pC3kq/dREfW
u41wMCL366QzWgaSdBZamhcATqiUZSjon6qbJHPufUNMmU0qfihXp6sMy8Msu+YWHL7D/TYfkwgo
SYmW5iyl74Jf8DnREAAM6Zjs/bemxMAV0IoT1D16QaZBFop5/exVVaOc4/9dHYrh7/WzBXMVJEMc
oeISzdQ/XG3tzk6EXaQ1VnTdmBIufxzhvCDlz/tyRufjKlEEztFf4WHdshRgZI8kg7ezAnfcapu+
F1fgIaGedSlLU8iEFdZBp9DIZ7UG8pozoD8lK4cjHWaRgf8hizdVx+tuQPphp6v0WhwmMuopQsQR
1YsxYQIEWfART7t0Ih753CsKQ04FSmeIlUJeVRzR51/Sbr1X8RKyKQ7n/TtkL3f1uneyenar+WTr
Tr09xOZy3ytJbB4VZzUMjw+ItgxBwXMchIV63QGNnRLA4vAbG232WFOV2wlJgP4SddXK9BuJ69Wk
neCo4MpBhz4DE+o0h4xxtx4Raa/vEoINmYFIhbPpo9gKm96pUNFBWKRXtX72wdzc9QeR5X514BTf
r4jX9Deh/NrZd5tf4ebaHf7VC4U72/IrFGHNGiDOPk10ko+9uw3TM/ZhHR3T0C27ea/VaIuvgGF6
Ow60bZ/t60kFpfV0If8MwCboJFDlEZsEKjCq7Rxr+quY5I/q1PczEGEDzf+S1rsPHPEQ9nCTCKEX
XwaNYNOgSIRgQ5ifxbkn6CVlBe9x5a6SYkHnP1GkbxW115lpaNT5Jywb7RkuYku2mLORI0Q7Gj7I
6+d/WNxGi2Rv8JWNuw4dz9TM95Bre+MXf5DqUPnOQSAa7jPslCojIkmjivG+xb8ec6GWgEg4RQDb
c01BnewL51EplHgFn9Hg8cM8Y0lw4ilvQOKuc6sSFeLApFH3QXvCc+G+w7o2wzqoikn8EfLmvfQO
UQcJQeeehIG5EDrExOvJA2luCSHb1FgaA91gKq1te4zPLHqapGcXti1SCcDSZO0fo/6WknpLtt0D
hTpnZOvAZrP28/Xy9u9ojGssVYBso9JjoSFu85nhPW+Ab+cG0SHDaCA56DT2tRDaaKWR8AzAZLeR
vvouro3ztrUQpX1e4BPGolM62Vdy7LFuMe4j3IgCJX9v4vReZK8TYKe8CqqHgegQAY5CfRNKdt2x
6zWN1p8eV7UGdD6qYYdbKQspUt6R5wrbGrDHdk3UyWmfs1Hh5wzIVWZhD4rERblw2k6nQ4YcjCHy
wtFyLFw5oGozIKPxlFOSgJXyMStIShxkcN89uBNwmBsVJE/xrE23aFhpodVm9XOhihDstfBCo+Mz
rwf0I+ODntGj0e9upZNRbZYU+nz7ZVcvD5jYdauxPkU0AnhliFfL51EUItmy4teofbcp8CFkcZAE
7pSOkLcQsoKlhkBtf7vng8Iw+4OIOyNtFk1uCJEpprWv/qnzq/ImsZkDOHSuoxRHE8MM3o2YiUlo
VoPEA9Ufp6+HBsX4zgg0mVTZFfineUo1IFRgSXfBJxieh8cyjKsA/5wMy6mPTHXbGaDLl9dGCfuJ
LCOeEcAeFK81mix27TGbPHsrnAO5TdvB3SQWZdJU6TC+D9Yt1KFlD0BpuBttNNGIsJ43/JZyzhZ5
O5oDoRzN6mPBOKNuRNSMSWl1JYADvVguPpOIsNfsd7fuOe7ivkatMAU4W3qDwXq96M0xPFMc7wK8
GF+LAKC0rAhy7abHcCGrruQm3MB6yy2o/3vtZOH2K0HV+igYwjX+0LFSsqYrjyUtNSXDiHR8bQRL
/Zng14XdHDZzwOj4FDumQibL5KuiY+H9ktWew3e1At5Nudhwgpeqyaa7Pvru56rBfAI6+0zk+ZO9
OAEtCbmyn0EhdXnWnPnmgE2IWxvTuC80WKYj4WMPmp/VOGstJEbDaa16gHqImdUiaUwC8/yUkbVC
Ne4Vu6Jk5H0t97IPhROTXeJaDXy2Jhj6ofVlJjJDf50/3y7tC1drULg1tdlM6zb5vD5qTaGneOwd
l136Aw7Xo06F4zf49rDkUxjFcg0G/Vsm5KzyGE/GilO28Bd64XZI7CST/QFm227PfTJnrtVXZ864
fsXc/cinz9WxPPDz87E1tecEwYQ7h3G8WwXLNQohhKLJiOlU0/MWd3Jl9YdszKIVgW5ZsWF50vY9
63dBkGDpr36Ef/DP2sI2OxdJA0Ehr/mgrlR34wGmSCGNY1nCodtT51EBxkgLMY7B5zXDXhBGtKUg
cVBhrjDzjSOi8T45zB2bKrdoGsPySZqskvgPT7de1AvjZPZEfKAuqUW0kqO395EXv37vuw1ljLO4
KyRksGw37jMWfVovmynuWBvOHYq1cCBx8rVBQiEBDUNKoUZn89xvOV+UeRd2NrMYbUiCA7xx2c7c
o3+lfYIzN6OjixLI3q1SlAe0tTcTtdnebQCtR82wzBFOGW/ZmhKTsSmWru39fmhapRvGkV1FArs7
n81r8Mo15SF6sCfmiPguyLe1o6Sf4ALUua22aOGl7XzkNToFXSJTEigSbnJ5cR1mgrGW8v2DQg5t
v8CtW8cdiGy3FyFB7QOJtYWi+2UlNxpcOS40Sy7LbVp2Xf9fgVzmrqanRF9IdyeUrz1PxVuHqeCv
9cXLWsBcEhyqU79o10HH6OuNEQqzzMsdhltuFlbfgWESm8it+VCqaG+82/+F3lPkkVeLHtAK+ZoQ
A/D3oG2Gok7LIyDTy8Jlfi5bDuTI5xEAmM6YPr+sHYK0MAFtV/ByJXQ6YThTTPNus/tNRNP6OgTP
/98N44zBFRKGbYCgwcZAbjz9SlJXW4Urf83K/woZE2g//4/cwtFMZXeEnTRe+91+x6txhudrCUQ6
HZw1UMAw+zXRMT+RwUWNiYBx6AC517CJrc4GMRlL/Od1WraFN1/jsnUEQ5YmG6S7Ehmt/ELdXJJY
CH1gG2oKnhZJlkN32/WQx9bXLSnhqegQwku1MYcfVZuimQHXGEfcjm0T3uE4RvUgbzovHYTV9H99
JeWRxmkEwdmo36BgdLYXAz/RI2ZHxx8tV/ZAFxObmu4k/+MycubTIkCck3/HUzY5GxighQZNvgHz
ZyJnahDITZ4fD35gyyCXN06NcUujYT0UOGcg6p64Dq4OBZypNLtRlay1YFAP+x1dYoSjlnk3jOSt
EMKMejjm9EmSlEuie63w/Tdo3ZPsxv3nuOgX7tSWSgn45tmfOgpti8fkKaCdhhXKvw744fUG4+VB
XspcyBU0FU90oYEk3IlWQ78wr6zu3yRRBcBSx5ig0OjJSLDSV2EcrgUPlJDHKlveitQEKR8d9smb
Dp7yFTLz4X5aXhVw2l/NYW3Vuu0ON/kP7NwG28h90+VSgmeWFmb4bvz5B6HBZ5eWpp/XIBCrPmnD
18k0yr7lEKxnH07PgMvUDkc+ivQk3pj33I4hGwYQVZmVKgiVrnPJfCGpV+bDKtx2+qBEGfUDewsQ
Hz/U7Q1D04k8bvdADPWeDdVmU5XkYhiK2YSF4uFzLx49xUZ0ELSNQCv0YlHuaVwfJCkF+IFl3Q5p
fnQZjSschrQTXV98FpzRDvkExr1WJcRpMHKhlKOnHoQbdoeFTcjahndq7smEbDtxWVla6wkTeijr
DzMZT7AK/akzdtKxZpcEGkjbwOz0v/Ti8O/d4gFP6VnL0OeHEZrwvHPero8Al1lD8fyOtqHqaG6z
2O5I2mLoy1JboEPx6wpKgXYf9M2ZsaLykBhpM2buaZkbF9NTOjJZmM8TO6zfsLtH6KAGMyj1WYPn
OdjvE1phFudfN/FDPDxRuP1O4ya57y7c2TJp8aCFxGxD66EuH1nsRUGSOhynxXjilqhRB3qcyEd/
E79H9ye4F6CeUKoqypW/KaEfTerUie10Gu3QOB3SWtSNh2ZeQBmze6DYFGe5DpE5g6boi3hnPWRu
78nyrJ3JnXOTwS8DhZp3Qau22YiYNAAI68T3pgGaheZpm5D1mAcFjcHmprtiA4dqjJfXOtXMbVk9
CFDUxC/RsI95mWirdbAT2u4aT47Joy6myVMOfS5AepbZPJClAJO42W9dUSAcl+FZ5dJjE2BPJapd
ZORBDD/PElgyjixOBRAjh7J3+BSicedly+bzX8+++a/FJgLMOr/Y8qA8yL/ndR4KAgC4o38/oGOX
BYtoRG+7OkdwN/dLY48b/myKnRKCRkSMqmf41eOBmifpC2amtpe8qK8b/W5/LWF9fDyhWV885SSS
XCbmfa9P/7XudnTTgEz8UHRjhXi5QXh/zoDMguTZm5c4sKVPygvO2ROr1GGnEZhnM+htBGde0y1t
/2i4YFfDB9V411duq52diMH1SKx7b/YeGdx5nDmF3cGAexNufvNAGaw8i07OPqG2/QoiVSmwqJ87
tH2xqqFZSbOGdleXttNNxnZ4Wa6g5/Kz+oD+ykzWAQN1kO7eDGYFFyYAaMkjkatAiH6bgzuyM/62
PZZnsXuCoMXgcZcRNAKfcQ8Oupzp8/HIf3XXA/RtWdJMXcZX2EDnJkwBx9PU0nDerBPeblfzZoUh
QZQ2a77xch11hfZ03bAHAvjOGUkptHPNVp5uqsg/IRwKPspCfNsFr5mvp6nxHX8aHp7BelbpXwPg
wojZOWhLWPCbTYiCkgvLx+97wqel+qPaGI8M+9jYR/kU5fl0PSlX0VSutn5MEU69TwN29o0/A75M
vXQapYaE4sJDWah77ZN42Av6rnjM8zo+Q0wHNuvMfpWS6sdHKnzs6KtEaPs9dyHuZqdiqfpZUY4B
sEpoj8+Yc1JMawuCOygTD3mZnsgNkLKWrn4Ta2AAkCBtgERuBOzdLU7u75E056FEQvBoaZXanMlY
y6JoS/CRRAYG6Oh6dfIVHPqQcKYYzFGJP3SK/7m9I0z41ybxyh/vGIUXRPeiRLahNR3rvsibA8UE
eSGSicazyj0oq0wRjzIXPsFaVJ5v9TRS2dHvyiusN9h+U66+nveJg7xbN2Bjoi34CUkmRmAwLCil
qVu66spV3gjCs9S3KO1Z2Qp6DU3StO/qIBrECUGAY0QxrwULN0HvfeP0D3fgBtXZITanz3Dw4rdm
vLZgY149+lurl3mCQ1qGRN8Bwx0hTEChm/2Q8d6VT2CiLBgaKMRHxzeYlZhUxuaIaWUTxhia75DI
jPicAoiO5CNQgT9XbMy4EdfwYjxnSgA7yjoBezq5m0hMD00LS49ry69MNDECbHvPRmdMo2GPNlrW
C4N1lrbBzS4KQtqRKfZSBXpVlIDKrvXNWjuZKklOfLpqc12pSf4i0KsWmljccTPmkO4tYdTzfOS4
wk9/YWb4jPKFmFALp+xu655lVUixCuzB+aagFsx5oP2dgQ1nAmVKhx2P9XBZ2jnccRO5cadGszoS
SQYVIPWQRnk+MdaTTpS5MMB7sjEC/P4P6ymmi06aBkNtnmKiSo6XLlIltxnZ8qPd1aNDVvwr90H/
J62/m+bzRoE3CQMh2T4GhcFQYZ0ox12kg6l2sL8M3AAkNzXKIG4dYWIuTTC15ceph89Rn86KuJwT
WszE0mQniLg+ytFsxZneql7VR7rKxBYMUUuJ5JR0hlaGXycLi6jfDw8CNgV8zq6HtwlhN/rHIr44
LBFDVtVjobuwK6fW3xJzNKMByq5DsxOd/N/w4qTWQQx7YR5tImIbrlEXdIpwkl5sSGE1Wp6AaWoc
jN6Kpb7RaHkEzDvM8MJYXrjEbT/+AT8Ke2IbptoE7Qxdm0YsXUX1kV9vIl8apjlNCn0BcaMxXfbZ
3P6Uk+zVAl5oXbmCiMgLM7PPgNaMP7nI/HB0Q3I+8nkluKxi3GQOZhyQElm9LeHEP/Zh2ZAqvb0D
1FWRXZuGGCtOmylV4YIrWhRI0kmeRdimT6KHjAnZOq3rB76x6A0aP5KsjNuCy802ppTglsLHzJrG
imvPRVHgwL6fSiDdDhyihHPrGdeUDaf5Ih6b+w5+HIicivY6Zaol1r8N7z/zhtzjaVdYJLaz4z5d
PovbObJGgNK+tiXV/fBt89V156d/GTbHxumodNItjZdx7RKSJ/KbDDXBwZrS597AB0dvs69QY+yl
WPF8fNuTvII2yAntYLa6j6WDDsiIzUiynnyEQUj6At5zIJHEtnwp7oVpA2w7IPORTrsym+690+zr
uKBqvnVnnNejbgljjWpZDcKTYpv8qWiL3Rr77gyOMXPrSOVI6ebiwRDyvmQ5VKtsDjvPKiWiZPOD
1qSJmopm9FhheApeWInyOEu9Vb5WFbtMDQREGreffahXOLb5HW2EZ+1syyjrvGCYWS/OjhMTK4fy
QNqTba7kOT+o6PHYNG0w7mAxfTYs2A40tPjS42uwkv0nww6YdE75LiaB19ZSbaTIUlIjUI8Ke9q0
Ilow1MJFAv6i1NQ4BvwntJn4JVhXdsrmul0sy6HG1tNPbMiXrJWoIqRLeF9BRLJe9HARatCGR1At
VTo3bRKstV9gSHltFFh+QvOD4VPYGNXT1zjWtO+sHsYzzrSJV6fmYH6rtxPIQZSiIPg51EeSqAF9
+HZ262T/MwmgrKBWIEh3bWuinZSbep0ENGdO0UUxsuI96opr/R+CR9UmrsIvMPN95xui3/9LDk9C
2Di3OrveJdGb2MjVBRh2YErPAC8vf8w7ey1vkOa7/UVI+/HxqT68GzcfSauZf8tYGQScw2/+wYAz
1NthXa1Bxs/fNt0Aa0Ku3XIo/K2b7l7124pMqdztj0ieGZVmPJ7UjcjTmbiTmzbOtuzA2eEF+sXT
nYRCYiEL07GiNKHYD0zfahDPoa52LPBQLxTM8nuJRK8S28KSd5mXhYhfQyEoSZxFfx483ZIbYSjs
eQCeMYAgRRnYsILvRW+UcKlT0Y33kqkjeihVpDLiZBECCqJnayrJ7N0StvS+hBZjtoSnejn21aV0
g7Ufq5FSxwOU+fadhPCsOX/bx3BSn8MeDhy3lTHOYtGuJwyBZkK2GRINPGZZz08vSmZv+KBjOm6i
fYybVK+LpqBB6xxraNxwhcvz0vEggtNh6kP4tq1VHE519mX4frPezRBDFAPLO1Zm15KYO83jc3L+
KuejMgVKs9jp4gu9C6s9uiIvwh2FcLGsmc8WImF7ouJofcPogXZYfI9Y0YYXRX9D7OosQQiWLnBN
q/xPpXwACGgjJPRmprIIn0Oi7ejhQnuNbjpZsCo5XHJOu10O2jti7jtT69P1bmnyd1naPdhbfyMI
HMPwtr7f8mZ6M0GQl/KLSz+qhUg3Z1uMSA3x4Lp4NtW4bblC/SiOnLx9DtZyVvp9dKgHZPYK8TUs
NubX1sp9+U8CdRXQkMp6j6LJWWbza6gNE/L/Q9n4pJ6nkixNrLahUdYoIFShKYnL9bUAa1kotN55
aNSCu5V+VDyFqtMVseLC2pn3nu0sS6D1+teqODQbc4pruYd80wHE880I2Dd9jjuElwSaFSlyEqvr
naDPqG+ViHKrNh0iLHhWpkcT3y8O0EMNpmLj9kaJ3cpCQeMWFCvBTxLEjFknzXboRCPkRIeBqCu/
f4j8vSoeYHD6RAjIrT0CAJksDyxL3h9HNeoyR2dH+5KYyeMWcwN1zoI3/P56DiGeDhq4oGL9rR0d
7rosZc0WzzIwO2jg6NOYDoMMzlgFV2ma2BKh7a3895Ew2JBHKl1+o2F06KWo3Yb5I7/WysbbGBxx
dor5wrLOwXGMUoMkoiaDYwe38slTpfzgZ2IRIpEwZVUOGz+jcl33aDEyt4tpGAWOqAZ6Agut5Wf3
h6NgrQMhdcvH8RS89tzksv0AY+Kou89yShAtMgFj12/5QcPxjAow2fm8FBom9o4NmJfWCVHhpMQP
3rkvjgikbaOOs4OXTwJGSPJw7nwa/lt55m3iHPIvHZlqGIvCxQd56RlqCrHp9eRlw2eRsgc+Fw7c
le/PFcHOAGvhec/wJ2tJS0feYp7Mkym3IfDwtSCRHwJV0u+bwUYqPirWa1AEDLefz1ntIrv+lUcl
C6oCPolk8S63SXU351bmtNdybNeoBLYFsoj0YATrq/jG4RnvaLcle84jkYMZDorZ928y9CEnst9Y
N95ipSi7Um2oJMzwmagcQn2gfvtbfsXV46umtxDlBH1KZ4cyZNd8YuoGq3jXSjILVFc4D6ojfZu7
wqDs9qT09aLTZ/U0/CcJHoOhsbKUFw+Jl/QOobUlf/HqEfcUsYqpd4icnBu5a0ryfx3z7XIpZihW
kPVan9RZvzHwbllZzypi8Yr+HIKbx7XFeik0L8AsMycQTDnk3hELCl00njMRCY0bYkLkecnjhjZM
x3joFS71EwWQYVcvD9ScQW6MOW7rPHp2auN0cDsZj/hR28rhAmjIFU5xmlvn018JYs/xJ+gHyMqc
luv1JuRJ2GdRyKaH2K0uqm6Y63MRPPKM4xPhjiIRJXDvfJjB09DIhkUmCZrvnj6VsVxB87j9vGhc
B/umwd/rWdx0fSfoq5ug5n9LOUFMlRc28zaMf5SBkZ3o3hWKijPezNlj5HW9icdxtMFNk7rqBpLF
V+QeaMokvWC3wEpsbW4YCRYfMLX32nNocBfQVWbBn6OL6sREls4BoweRQ8DiDLarp4axPg9T8W9n
eir/6ucRUhcJBCf43dhAhOMF06ityc+yfaoLvWGxHRoV2lwRXQdwVL7WnMVDs9SpAQrSTgU8CDyL
Grb5uV49iy9YruIqEwSol4IYKZfT9cXqUztxuTE4N0q5iHd8eRh3Wd4udCaMjMhhCuHPMEizifOk
ACpL6tz0vIhhvPM2/ukkCMT+HnD6KuWdwXcb2fzNGI3cEUPeg6AEv9u5keUfw1NjIMRDSqQ3ztMd
ReYFfPT3kmq0xMf8JviYKUOe8meDPVCBELcTLA1V55n9EWXKW5KDV4FtPBfItRG5tPekpbVfF8vW
yuBtAmURpBu/txha3/E+HyO0RwCsr9avTOu2FQHG6hXTq2JE4Hb6btIEg6dR678TnXglL4KhOc48
tUSUJ8uohsq1EtoD/zipydwq4xNa33fShMNi3tZix+sPlKjBxreiSEo8YkLys1nnMbEY1KHJ3M/u
9ADmZj6mRai1Pj21ZwsquK3UNcmtzzF88qVDDz4cTtG7+Ow5KnkSIYoTo4dLUdWUd5s5qUxQWFpH
QHaL+gDSweOWn8Z5Im2vrDxoO732itNfvtmLd+fI7BN2YzqblC/Y/GIZZ13ECmDhtUVFjSn9od9h
EP2n54JD5jpK6Mr6u80JcmY70hzwaweWC+sd+bVR21PCuM4T9oCGT8eoj01PhRLPz11VWz3XfIov
P/kTylv44hBglvpL0w0meHM5nc2Dpzso7cdNPSvncr75R8oEemlROpSV/Tcb4FALl2QGPYytojuO
5BevTs1WpoaVdno0CXtXTL6W5ZmXGlsZZTOybcW5hEisPTlUEFoorkANJOouvB9w7K41A5fJKLVr
RZAy+Htp+HzfvOGqTB3FHKPdcrj1mb4TiBbhHeoz7MMoGthi2k5XIeCEm0G43l5NILvSgjm1sBhY
1Ywav0PXgoIJeiEUljXa1DmV6XdS9oBzO2wjnl6ScRWJOW7MH7s9gNUtwQlcLZ+dxp4AUQd7oGsu
Uq6H/l4mLE44SNMC1C6rFyTuBsXF5s9dq73HIm03dSvPOVtNloL52dyV9HwSz6GHFTpj20R/roMS
g7Zj6o0kZC+7pPbL7bLaBpJ+q62zWEDwXrybNO03AFjz/+j5kWszCTqm/c18BeLLIdsNWzN7W/0O
HY0Y6JvVeXVww+IgnGW5CnX8phrf4h4aj/5dcDZL+XZOQlojJ/Q7k4EcUeHQopeCzQH3iHc3OYDg
TPTkFUbAEp7qNHU149T8+ysJnqbVk2Q17+2TK92bXRpRLMjJgivsUydqsOcvanRZ112M+LrHjbPK
YDn0V/g92nGungjEATMOH+wVEP1nKJFeD+Q98HMlgLW7qVRcSQJ+8Qohrgt8AptQCZvMC+y1RcXM
hTqc5DhSBzVmw+Vmc1GI6CuzqWewG78aeCNghqMfxNBW+v+/A0JZeHOCmNvFPFLtzi4G5aleyzti
23Px5Tn+smDHHQv/Krk5hx4/ByFym2oHtReqlpHLzlZFCblY6M7laJ0HTA6Cpy7wxJNogFQd3qOH
vryz+Ch6qOIU5b8rM72cH9lFRmvWlamHtA1tW255pDcJgOmFDq5bzFrt5W+bP87EJQ521sPihwqB
oQZanIjgvFdbBkP/D95Z3Y/Em6Xg36wuwZ0Whnzixwj3Cdb7mqBjVCxkqiFYZVunPzdJ65oFaPEp
Sl5jfOl29he6gtw3rnvgVEGg3I78EwIvdAK1Vk20yAKb87CQ8wCbY0HD1WuJL/c6/KRi0oBDQs8m
ETqQQ149FbvZLGlqklOXjRR43Xq7gPpXuV14YlB/myU1ADm6b72q7TknyEeyA2fSxKi31dzt1bzM
a57ipxV91XkBIB62dh/PNs8WMD78iFjQ1ZNbSYWQhLYnRQtcNtAd8hMZ8zMDM7MuQ4X8gDcMNtz8
lWpEbh/Mo0O1K/gmMV0fPtYP0QXdBhCESNmLpROvWQRdYFOCKhnox4LTggItbO9ksWwLxc8tcvM2
dt7vO/973Mr9MMo+ll4G+u5rps2MejcP9UnMf6b7MYG/yBlQ+5Fls13ngVdgx9wjkYhoztShvy65
f1OvpRTZejMuU0MOzQ7dsV7M942+t7UxwNVjWDhO+2IMyRaEb/zBdCge1bL8jBchYDTg2kvILoWD
+qENIvezCDrLsWVwQ7MQ8/LHnCiXvJ+t4oa+BYv4CEcAubni+sWIlaIlNjQYklB55VdeV5FWyICD
u5O2wArr1YlOHHMA2n7NGj585vVJPYJG7xZBgr80kYNq7QGSV6sbuPKjYz4Tf+Sh26gYhmHMjO6F
fdsl/UyChuKlRHcTP1pVDB3s2BcKiCZHqTN7ZJgnvt5b+UeHtBVmsj3ahI9f4ril3Pz6wEHLo3nT
qsa7WR6wRh5IqikGUkBmZUzW/ZUbOs8sWYuQwH6eOeeJr+/+nMtP1KIKcPaQ9RfGcJxOeZfQfGiX
g7aD3SAiqWXie5cWbqi5qT5567mMzOt8flZwr+rvqhwoBxqr2p4j+JwwgRb7BLgahRBXgeS5hM8/
GwJR4usTBiKcnWbfHi4uP0kfssKmILk4DQT/W4H6HnVT0BpOW8G/nfdG9itQXStmgL0+WfiU0w3m
3uUajPlUFZEmn6++IeaAKfzFNbtUBoNZsxjsYO11ZIUhWDbLCCALiqQikwRMK4qvMJb5rncFXVhG
ICZlIg6TCIrkR9UltCCS+H6BGrWj45wP6MfwEDWF5YqL3V9JubStjPZNqjvJlvI0VIm+uSafWJHT
HFti5EMIVYWNhUNKh5Iub/S415nudaS3crhHKOuzZ4mMCODGD2pKKedhVLM61t+ATa8PhEsvaO5k
gvejpGzqxKTBbE0MZb+tlLNzNU+NP26jLTeJJ2SrsVnGiJgdntUT7jB4bgqBlABdbI0tMkrBYrXC
EYR64MhR43woLQ12gneKT/t1ETArDMApVo0h/YTBnkgqTxR1Z/gCMFokSVS/bPe7ANcWFvm/P/rw
FftO9RS33hWaRYD3O0JWkkxiT+kufcJsTaE1TewxFp1euyDYH2D62+g7fkIipxI8weJI+FZFNPgp
E+hrLvU+EgByImGc0Zx5+pP1DjxdJhvfgzIxJAl17uJxvBa2k12nlEl8Klc+OHD7iEwB94ev6+zN
kCkkzQLLb+seuWWzP1uTrODD0XrYnx18ORsNLkbwATvGdWmLy5bnYz5YdFNztYz5GuRM4HxMe9D/
6+icfRNG/9JIslnsczVFvXdF/fawW+qP7ko74Sj1ahs6VN8KvkWHLTU3AgcDSteH8MPDk9bIlLSG
Iz9dgAC4XfDU+DUkWOP7SPp1KP3L4tJp2Cd50jggF3lul5o2v1Fi6EjNGUeyy+i0CJwHL+90kSAf
gAE+/y+68NbGTkyR5+HoZC3XHcVbEqUSoX+LggIocMOYv3YvehnNtAyjm4YJDq5joGGQxDdliIOz
07/2cVM+/ncQbgNjzLgmwl3CXtNtZMV1MUTuz4BSbxZBeuAGWftF1S40rutAtWDl9T77nyZOkr9D
zeXSA1dhlVUl+XgafRXasbg9J5BBcBoGY46RMa2ZPIvtFQHIq2NgZbENDM6KJTw6wmQV/an89udK
P1vbdmB5r5Amd2ciJeu5VjbrMll8mslmslPFpGXwk4wkIqGFuI7oWcqmAysswzOH5ylcEJVbrWO7
SPcjzp+GuWMGhV3H+4kUsCdCTlByUYs9vgRHuqsipGDldlbzyIvzWcDsP+Ci/1+sMYf+9JGlcJSc
LniR5zRw96U//yzcelJaXbpCC7z/F+0CtLJ1Gk18VolGUSdigDvcNjRx0oli567hQKM3nXHlUaK9
zRUoAqdqbrLSQsVdVw3xAqlYCb8UE+f35r8L/loMHm/twhc4NN39zEiWBIZadoncqRYDTCjDqH47
Powk9LKcFHky/bHK7L3kZ8HY9Zw4/a53NsJrQs8Lefr6q8cWD/pH1BcW3eYNNaLSX6DOuWmeLBvv
GqP/LOdAxP7VPDB96Hw64oWlNygsO/CTvq5I4WZj5QB8/w9zvvUmWAQhQkyzQ8hvsKjbMOMdMo0r
/MmHWnrlrEuHYT0Zu7vCGDB3yvRsbEP/YjMsULPENbS3JhvkyQMeukw0Xl0saWfa0ZiKskDC3yt0
6LZRFf3hScIQ7URRM0K5K7FNrd5Jlh9JBkF5OwT+8I9vLvEZ1Mj5ZpIGQ0xvqoUAryH7/BjiaTe1
ri+5lQs2XLlyv5JQWBgAsNWnPYFEropyr/vJ9zZCrA8P5m++1rPPYc2Gtj2M62ziBmXmqEylJ+xA
i8HVdAwE1vPzaLAE+wZWp0tSM2a4O3w9kqfVr25d8D50ZloWDXgMSbHttApGZcW7izCa0AcvDjTw
Yj+X62BffHZoKDDug6watCe40CUkTrUgZcMnKZ6CyVlKIE9Gahxnn67UgQ2IptAffteOag5b9pT1
ydA1sfTGdfO07lVEsaO7hPxTryVQokgRZQF2Lpjiz/wvCDdp7nkW1ONj588edHcX5bmXmDC4gFrL
0VDe1p1pjkVTb2VM0EXpXjESe0adSL0eLV7vLfcUMHXSLjbv31UZQRa6DE3+muuAl1QO+Yx7Hm/X
gpFMNkirzbCCiP8WJSo7+ZuLzN+GPC/kMsxGIkytiHcK/keP9IMf14mDCyvZ2NT7Lqp2ZPahttDp
pW2N/5fX9/5O8vo496w79hvlbHNH96qdptcEHSajkhFnVISgvAw7qgjwkypA6p6nMKGMcF7l/0eC
YrrEWbBbxpgk5UHo5uPIA6TVn1VFpivFNQ2SpLsbSWzXqGBWAYN2FJuLEpKIIEqV/+zmRS8b5ggv
mlfH/XMvUwOIPMErsQr/diXUBPaEayyqfXEdqvk5ZHJINTnvyDypvUTrqGGtTfrOirsuBurGwQtc
z8h6uwdvbnhiyCUNZt77spBNT4xPqFYkvfjd3X6PT2cs/1E8msHeuQ/w97D7aBR6GtckJV9kIDOK
zLIkGi0jhaDoFSvUSJf30z4WtqQcvf5jbX1xe5/rg9TU48Y+vKu6HkSGrQxUEVisN83mQ7Qebwqw
Elxg8vcnhTVMMD74j77spIwXH99gAjNAZoBNqKL4OKrZtUFmgSaTed/I9sHWY5YOdjTennp/HIUb
02wlAi8qnQ/4vNb9RjVNvypjAUqywbwsXpBf+eW+xk6DNACQIPswwE7xNzPyib6Dst1j0P2N/cwb
XS/a6IowQEIadWiH4IXans8ofLVwB93g51RecVtwStCRzhVtnfAuzj1jVmzrZyq8szM67NIJA+Bj
Xntm7JQyhxuX/BsVRz1VcXa3PQVpJdw9QLa/l8WSY3R4mG2AsDXDb7NTzbPZ/KeFZRj24I5jA4LF
3z/sso9u41/dCi+s0xvpESATgtCAQOKP2gq+shBWeOB0uFjocaWvgmq9ulfCxNLIVtj6FLxRUE5D
FELFRVYh123MDaY/b5q/STLLCvVHs4htJNXcD57GIpKLBreLGfu0ucfX3w7gP7vwy1LrjiwYh7rP
08i6ej3cTGnfmhZoA0Iye5up/qUbr+5USR+Edr+CNHsnCPciQ1LL/nHKwV71WqPdUjzyA5SkjElO
LnTbZ2woJNIwjzrD8V5pKLJfl0Icd057d8dcBsU7tjHtOigq1GzcfinWdyTb5fn83H5bG020n4wd
mXLsKERbeQxOGjEdaWpnTmEs58MoWfowQ0PpQgh5j/ukcPLwySkN2KLgMfIX/7RzeA+IKVIfP03B
vQW+S8dpyxcbi1joyBryYtlFrIfNDCpvVXPG/WFBCHc6hEte411/MVuEbjj6kovi1ksvaWlR/W5C
BzuhGC6VNuhyNqk1o80HzNtq1abMH04Yt/T6HiyxE11qpKHH1b8G1UWPwcTLR7VLR3igXQM7pu4o
057JOAQrk3x6Vs69jqOmLMFs8fjlbn/ltJDJb9w+nuA3PprNqi+zxlx/npaSGmrZeHADELpmvNEp
f4WJjEaZl9jwJFdnvd8Qk6Dk7K7uPPfgDhqpRzFh5jS7IkDwsOvd+YPPzzQRRywmmjxLmdZrkqYp
Dm1B7lRG7Ibeou+sL8AXj10XrUtyhFyG4LSNGROYkTIOcLJvtLMGzjt7/OM0cJmoBmgVRy3541cv
1AHgx6bVD6O48qaZ8epEbrUoVfJL3u8PoVXn6F3czWQaSgjBSfAk3SaO+ao0TSlDWCHyGSX82SjP
hhVw7VmRUI1voyEQbXJXWUlo2on46ZY5uNFHKlftWIfKR6CwxUclCuJCpYUTRq5YDYYeBFXE9P4q
JvoXP9FuAsLvL8/iQH/WrFlPHYqqfKo4+q4Ueqy58kl/lmie5twu/sy6+hMpgO0O/lksPxTz9mPd
cdD0QM2BGHJAyE0jOVYu1Qj/x+XhYdoLNpYpvPs5ZirBakxA4lwZv9VR408m10IeULYo0qwiEhN5
nmwAu7H1SPgfmI3FMXkiRq37laRSjWFrk1wGlrJLNCNHta+Z9dzEgUzj/p/XLuiM20hMkjNv5SrL
wc/ejabLX6nK2Ipa1xD2JOMjBz4DppN2b6VE7TOBdYsE25Kb2TbcqKydpQfZVYy2Sk+SSIB+Qgjw
jhJA2jZBmObFTw8B6wjmHBy92XSTdiB0dwFCHXWpe0ycni2LtZloIjlXG0ihNvOk6zcqfaHSsSEk
ZwAJPdKdSenzovlVX/tiScfCwG9YUCIRnJ+8FOV0zWRdNmf6gir9hm2+iy8/QedsFHrooE2yEwTo
jC7mFX4NDM84xOLGT+nSXSE4jbuPpsHCfLiz8EE/EJx12WlpXBEVtdXRTaO+YNnZcVcraTNb5nYi
LQkkIGfP7tQ9YIHPjAelk7TqpWb1K1mrFqBsLXiPQ1q5dAbQ7VemVUYCxJFgra3nrNimx6WCipDY
Xqd8FV7HlI2BiCPzCb5ysjuvEfl0lQC35av+MtUhSC276Amu0YAw94foO1uQ76kq24INvP8RKCRx
LknVPatyu1Mf3V7sAeJOY+e0PzYW4VK2l1FK7AT0almMe0yeP6Am5mRFTUJZb4BXHMbBLQIJXrE1
vF/tgAVnWGvA17tHvsFzbS7Ng+H2p7Da04Nh216oJjd6eq4DCDKDMpRYd86XlEuJ7a0O05KnfOQQ
LUDP3I2p19K6/Ia/5z+Lljb/baK5WI9nFCDaudL2pDa2Y0IfAbjUp39+SJphUkfo7FvzYoRVjD+z
26spSWDoh5m0DU5gO8r2MQWlH2vOoNrYYt/ggCDYR0obLzfmPTxifc/3F91PUOaP129r6ZeL9Jfb
1cNkCRXitWRS07m7SbWfoiL4c/0JHcOKfuPXrs4nUBrsL1nA1gV21ARklKH+u8F0zlXbRUbzBT2o
r8yrjkGt7Y33QCrZyb8jXmjZvlvSwYiDQEPgW7uKGLyEuLZWoN6uwhomIQhm9SUWpw2yUSflHQEl
Tb/CxJpCmDfDm4Ed6FmOk50yH8yzx9Bj/a6L2JDzgll5Cba3Bgp6F3ribxyBHHqkOZ/WWn4Kn0M1
I9tvJeF/S+d3pmH3wqsBqPP59jibtBMsBBOX+lwPGCrp60+bYDPON2z0Xf/yFth01nL8Aki4CQ53
D2rRKJB0xy5t9TExZYrtzSxhE0xHQ/gVdGlc2z5zjFtajJnRqlQsaqDQLnA+MDxiYbAU302VU0QM
WHEYNhDrGj7cdXY4yUwtW1BDUh2wTXcHGdY9RElv4djtptvXl/HCxg45TZc+wrS/fh64UMhfd4Bj
IsP9RKvyFLmmTfu19ubMY561SB1jW6/CKb2NcfgF3zOHaOshGxG3IXhlyKOP1ziNxjq77XhEHMmn
iHt5akFHPhBKdh/AWQXjU1X8Oc6ec5ioE8sBvLQaX85YxbX/vKu+KCUW7EAnY2NDhzB3HC476vaB
H/hZFP4ohNRZmrbkzvKg0ylFgIr9rsyoU5EX9H5S0IAl/++U79CDAE0PdbdHcbuZUVUlEf/dbUAw
zj14ehBHLKuFRGbmTTp1aZzSztDPZc3A7f16w9DUTz/8bl8/SrOWZziwXtzpFM+ahhQmCrUoQrID
M8VxKT3jDH5R41SwCy2No5PNg8nk058HtG6AeuhSDVAsZmBln/XuxmOb7Yg8NqkJ/w0NxZG5L4eY
xk7D6x+SvLMTq44owfQvYu3H7bcTt6HdLab3vAeGkLT2CcCvkJ5C/ChsAIMbe/bpfiXGDDF8eVYP
ksCnnnlS5/Z4e61waptVNroM6DXYQZJtvHYxh3MEwXDLkpD4XZw7n6Tjm5qQZDd4kxszLLkAWoFk
h874ZD1Hcp9iF9l9XkLkiGQNd9YZHVWeg+dW01qvaCq3Qst01maxPV6qjtgOAj6CmpNTJ0j5xnmp
ZPYQVx1FPOGjvwL+kJby82o68tm1XXkS7sI6CMVTW9RbIognzH0+6rRC4IYxtwMSv1M580sOUZQ6
fKY3ioKYxYg+nVFAOx1QDEAdWYTmoAjwCpUgpO+keBtPUojuhsn1DrbJi5EUDA7FW96w6zBv5J80
J9s89cNaDGwJkYZpaoSsWjZ/6+IOA3YNRhhDdBtt2dnuFB1HXJFrEgpmU8+XeU15pTyAhlA/+4g4
05P6Xen59lezKbvIl3Ck9xKBU7T+EzPElq4p15piXNZ/Ig1vlgZpEe/2G7qBgLV2GcTckNKr3CQI
bFMcol+GiQ6IuOH/F5ygIZ4YPVRfdNv3x1a7yM/UTR8YfgEodvKkJAKvFl7XpsIFeSyJnujDls3L
ZfY/uHuyJQN1vvQDHaE5DZ+27jp7lP7jeZOCU0dicSL0NHgxWN/yQk54qvgGk93+KQLsn/vxuB+S
aeqztuIkxAHXmLlIviSkWM6VE99btt957tZmdITIfoO9yCG1xokt6RSCnI3bL4zSGywklxSgGz5M
s1wyHE9KQC0ch9zIswqHmTzlIZc/lGCDhuGZPPqDjA/DeGpNhfgqrMezFt/wqh/l498JMFzVG4/v
ChwW9xauWWE0zXTx+67wSuCkH3t+CAxVD61JovMtQ2Z9hTIIBFx/AkXWHfelbVNLdTKB2YhvGG69
4UY3JdNWjWdVYRquTmUvNMfLjjE4Yf2mF8Q49BaFO9SFhtx+qYMwBHn30TeStPdQdg69Ps43v8vJ
LpGxSBLwOuGfiS/CfnrLMx4RwjmZ6sYdG6L/ZqP1B5uSGRH5XrrfD6L5no5rLThrfF6LSvZ5rWwA
EHNovYUbxUpC/RI/xO3ypmXstfGPIwuDXwnbgR51XuTXNSKVAmCqMSlioNfiW0AErhdGuCIWLxb4
zFfUwZWrQ76bgY3CaK7QiWPjapcwx6YbL6AW0c8ha587Lmx52pE//t7MYwTTvApSl42Zx/BtxlkD
LWSZEqyzY0zBZIQbHGCevPicaKIItd6ixAKrrPKYK7mUs8XjvfOM/HC1hHSjZkxnJ9NJp77BVL4H
2pal1DCm84TW3tbKCDpglVpViifjWoJ0G/xKymHl7SdkU3jdDdKGmy5MpOL1LPFhk7ZUf4UGFoJr
Gujy69IBF4btSqhtggKfykgvSFl8cwJk8LLCpHYDQAfhCVX0ZiUdgbbigImgX8wU8qVB4WJxVP5G
TcwbRVnz8TG+83boSRS70hiaETEllITqZlb0X+HoSnkCeTHLXdo7plW0woC8JA3gMTQKACe5wgYD
j4X5OghUrNJVpFfOHdQAuHo8oePeVnZc80M15QCHT9gDnuPtfZZ5FEhbiCxNhlxoHPAB4duY8VpL
1wAeOm1y121XjGIQpi5dD0u693DohdeioApuIaLAxKJgIn7WKKXaNJvXmfEPwGvzDA/eFq0gIGJK
PsqjJugYYPv7JvfIGaHu7NT23OijroJQn3beNddRptVo4YPkzRQIMMqGWfqBqHKZN4Kutn35bUTu
sFgLS+yaMHeT87uD5USS089gvKubswqAiuCVe7zTj/HjvCzHK7Zeo14Hw7pb0jMyoWWkvTvGMrZi
4jECgWGgFvaQHtIwoIu2CQBB0RBmwF3GCvFH6xFHXr0l8S3G6y95sXVJwRqYPba7/T4qzZS2gw6p
RuT3s+HqIRWLgcOXaFIrXHSVrmop7BqlhllnTWWL4kyHtdnsZqOE+0TP9TgORX9WKg7wtPKU+UQh
UQm9OvEhzoi4vgE0mmReaFou8HIMhkdiCVqYkwJ2+FUII/fKngkGalC/S4AafdAYtsqVOJelgIAG
Bk+RVgF0gpo097Uot3xysXhW1+6DViyMx0yr+XfNv37vx1Zigsi8txcZWn62Njd6W7Yz/Kl088fx
CnSe/+BhitdNTxq37hylBM1HpNP8Zj5I8lEuNsfnJAKd85yqHdCYeLM/CoCQNgVp28qmdmROjyqI
cCk2WB7+VetxQV14XjR2hdpux6vBSP26v/A//58TFsJwb4HvTilBCGQ76ozdi72orfSnpquKxsLV
Jua8tuJNibwnMuZDMJ3bKzRXv/hR/F45qf32jdDXNYJwH4n49RnYsgem3XDoiDJvSvj9qFkzi6Yk
AC5vEYl2VTz+j7GQteJO9sm0ovKBpzqnDPLJM8+VZMVkt5XzcvSRNqKn46aSB2BnvhaVonG+w95G
8vuIxktemQPVZgEo9WG0O2aAf1SZOerPR+Q/R39ZIcrsqdROATZ7nrO3USULvxqeF64RHh94GAfg
6cCdCMnmu28d0rzDJ5x5NhlXiLu8vs61VrBZ0tdCPkhY5PCTggHZYygAPDLh8wKIg2ec4HI8V38C
EZal1sKHPlGogklVdrRNMpNkmh/I34tI/0sSslZNsg3UA7RhNEmOCDY+ug6L9hO0v3kT3Fk5qYFQ
YwYK9UcWt+0cjcEQMVzbMbWqxHbL3Shw7cgHsO2vkwogtDLWNGs0UYnOR1+EGm79hD2AzU9E5s4s
N4gTEgBuqW0p1um+1f8AQq3H6SpOx+f3FUmsmcvrTRkbx29AWgMuGEhNRNDbqb90mu76hUlWoByI
S0Dc+Mc7fVygfEOS8ijxrf8/76vmXNQnE0EA+2UzAGwzNzJOH6KXV6HnFpfikZX+2xQlYakrXklH
cB8NSXSLli8JTTaasRn4TnQNqX6apob9sSWlJEb+RNGvodwtqHADDQxjwwAZQIioHlIsfF1iUXVZ
Pf+s+uBTYRPHQu29OIi+RHIN5vy0SqtEP6gTgMgX/JN4h/aXBZaD/lRuvaP6d2W5zyCJABMzLxr1
oNmiTfXiXybYcGpH8jxClQdAOY+sZvJ1qArytkXJ68z+tEzhPzCB9DnrTSUO6kl7nDgmvN2sK3lo
vgaixZQ3EdOrGIDWOkRkcLqX/eijv6axSNWvW3v2FL8FxCjfKVjXg0xjKdAM7qX1sDZRgKo+4obu
LjCfPioNkdTJSn5o7A4aSPyfm1dds6Y2jwE7rZ2k2qBSq0gFr8ivKOjHrwq0CiBc7rqM44TnJArq
hBUmCVUH0mLVNYu7ZjAGG6yr5X1HjsuBbz1RKCJ8sgdO9aZO83VJoMYEoRYqPkOUP/B7mnlZeomn
GzOTwH1qCysVjUujrupzdjTAaEzFRpHuH0bdwJ5RAXtYEhbAeEW8cc9Op1VgzzSR7kfE0xwV7iwQ
3yS+PLh++oBFZ5+Q15nLnEis5Im67g+bWfEMKOy70GMU5Fq9A0sGkNQnoS3CCiR5SIkWO8BFHHcW
hbtrUgRg+LrI0q6AbRqHf9OxU9L6ycKz5b9ASSAGqlnrez8u4nas15KLqmyVRxP2RdbLfkV1miLG
g1b82L12IGcphBmvYeUFKCBV0PNPOL/fEXzZgoV2T0/SwGH9+yeb5aVWSqfK+LyP5fs1GBezi8/J
PXD6f6Dv8JLLyaPMGnbICzRKjYFLJPLnLDEtHZYfdkN1rVdT4UFskmMNO3eTXjor9QCB4qsISId5
iIoFGQc7xTxcuher/95Plc5lTpKfUzs4hzicYUCMJXp9MpSh4FwAxgV7j+aJk2ZX7rXLqLYHTTOj
idEVQeSC4xkznf+AfrTDoMnxRG4qUlVg2YlTMuGCN1az7XfXlaSvP5GM1HJJa0o+tgTz0wqh+1pp
0IRGNExQV1ec72gEPtQvv0D0Pu8YfqgsMhoUq/niNhEu9De2nuqN/5a5rbMR0ACv2So5ig75zuPE
bjR7PJ4AdWOs7nw144Pw/tn5r8/py6ByrNAsuePN40WZQJpyv1Tx+bZe7Qi0Thy2VL2gt+dulr0r
Sm4YfWP9OkR0FlnS8oSfDuxIeUv4+ffKg6rvNmfUB0BtDA3Wjl/spggA86sL2Unx68PNMrc6aWHd
F0Kv26eCfoiEwQvmvK9jiuKDDAd5npqDHu2WVV+fUDrrzYvplZ7RkQOmptFlSn7kaiB+o1m7R1kL
PHjeLS7mxLB72CVa1eXgwpVvYo/zgcHnl2b07bsuYQBhSi7GAQeThHJp5l28zswSl3leFaSO6X8o
aJLMWbRApRkkSDbMJHxRsve+U74ge/66JscVwMu9jf9V7l7PSFenHCZd4o+6EP2xNORJ/mNSGGPG
agHGKkv9AZmnlJdLqYDWGHatq2QlBS+8wX1HG9P3T9RZ/tqrbwcYKIZq+YjKB7ZyHTR/3emtyn2d
FmzhRP8GKEPZIzDw8Wy8TdwLKvQkvsdPgOqJKM9arogZm6oUTIWUr35UNAWIZoRLRyrHAgp4zhB+
CpbXqGP9i7h6Glf82FeWgImmvPVAkqmb1Yij5e3C/lS/DKPkfBx6JEIu3jRa0vmJgXA9PBPcuwrn
Hak5cnUs+IJrXl5bwdLl4Aj0x4856Yeq1wfeHEY+Yie2U5rzk4BXWt6EBMXfissprigCtVijB9no
3QaXNKoE3rg7HDxb0EBif5M6OibR2h1hH3R8fBYjPxOggmbpbHS5PrK951Inm8uF1QH+o01uPpFS
Q6wQI89V6pAkNoeTWc+hVfMCsk5rD7DugGJsP/LGCD4J2p7FM8wkZvVmYDMJH5cRvR/FevhPOuNA
KtSTj5RjeciUNtKmAZUOp7yAvzEmVmfwHbb7NzzlzL/p8Jth3uDUEux831OGUN3IOLqb/Mkgh5kW
SLhbH9DSsHLDISVvvoJF+9RFPnqmIQ9Kni2+nhWCSOYJYmAwoMqX4SqRO6Oz1ttLXHL+LqlGWn/F
iYS5gs3ePUu0WGh8isfhu6MxcO26uZSOWxjLiYHbsLg8P7mrme2hp7ehd5IA1ehainGC9Hka6eyO
BFl99m/tTCzjNL807ZvMvI6JyC/gqDaHf+3nwSmgi56Mu1UDeAjlQkHwc4pL+F7Z2fKAnHKR0gwI
aAEbcPiRd/aFDlX0kkjv8oEdrHFSMW4H9mg29VZ5hYRLogouvAuqq50BPD7S3NW2Yb1FR9wqBikj
gELZ+lFAG3P5pSgw+xb06q/adE+FI94zROU3omyjupgi8BmOS8kFzXIpboSCPfSSatOmh9qxOQd3
mq2m2A3jOx7ALFqXjOaoY4F71k+PG9CxMmnhAVawb1hhwb29R9cckxAqLoosAce/LHCur6ItiHrt
o17K264IcEXqfVsiPQFLFajIuqSb7Tm6KsxS+uNVoyBr9656Z0tuKmHYcF2E1rhdBj4gInaC3aa8
rlN6zxu1V51pj8xTDei2yt43udWRuAK+Yj+j6/E7CzvlhsQKpWzePO/1OeTvzbI937UxvBjubGUP
vocfeZjwEqPLkXCGALvDtBOtCsQPc4geTM4I5oYmiL3pfVEnQuPH6DRVJf9nCFdUgPhOQLbsLtb0
jD4LyS5hAXuRdNcp4prqzlHRizJPBGmeep+mT+Vq1dR1XCnNFm9P4EpVTrpH6VYbWfDKdiuBTUPP
V0LCOsKpDe79X0Pj8b2i3Q2u4EmZ8LlcD62cPQhBq10qMxohhrtd5SJ1kjdWid8on71fUYsZkeU1
wDFeGTVDxY8F+W8qLUXU7OWeu5dvhW/p5yczYmlri3NuLI7AQuyAsGMdv2zFZvTuK5/XthjtutOa
5e6TIWDahip9t8Alee3dEdkmu8aSuhbhzfSC6iDt9IWYS3IjS5gOvk+Mq7HXhEqCd1dzcOyqY+BC
f63WiH0+ww2MvtAPFbeId3XXYCFKWp3P4Tkk3XZtNJjg4U53YpV8UXWIemO8t3kUfoqZyx6X+CJ4
ovZJGnlS8WBi2bI87yENADQ9mBQwsM++s//S9f8hRv+B/Kus8n94rUcjDYDMfS7kdMwY5MpGQxLR
k3powzMtq0bnjoT6EWwpwig80BGCiV/PlcMdc+jf1e4K3Pqs9uw/3pn1UpW8G6sGmEDFmyjJMsxt
YNby9eSrGSHtmI/62AJtHMCIyosl/YWjpGmNAZA4ru+8Gu5GxFkdkhN9486bWn4pjevTchn3STTG
H4vUvXX9+4dMf5yE15b0xzAw5TOoAcip5aZid1msiM1c0T9oea/2wrE8mVaDzkkB9yJrTKNcC+jy
uv16N4Cwj/pL1OoRUwMU8jKodAVWZFhckweAdZIyxVwiSWuuFW2+5lOlhWPoMkdjV/e+EgN3zJH6
XXTFWmvGdc9+528eWMMARSwk4By2jqmiQjHSQHMJC+UGkcD7Uc9qLgkaOjHEaN9DyshnL/bt/sRt
YMyYgCXT+aPKU9QHZYdt7qSsLa/gvLPbNz2dHZowZqWXRcIWMdrOmsVbNyA/ee8lHC9uhhn+J9pb
6Iv8o3DQgbdRg3NusT3qmxtVcGYNxmiYCThMPVM6xTBZ7aa+fl/2OczAIIfSXJ51n3epF6jnepOy
MiQav+obukm0FXJEI9eQYaPN1ZBwjVBoJd9mza/HFqc2+bKZqllA2zjGfFeALPezSH1LcJSZcMFs
R+rbNJ1Y398JvrqM+e0+lbbbnSGUVJywyjI28xFHxb7455hX9ggYQu9eQ4zBFn9kgC+DAf8QWvo+
J1rZZcTyMP54BqpxLP78lZeeW1H103k69dFQBCc9ISEE8oo0wkFm8z0j/zNKKvsS4wdqG7LnQDS3
LYqG/7C8Ni54KCt7AM/8qS5O0TIFXo1aIN/xY0KfsbT6w1fq7/xIi11gN5aX7OoXEGRwP4n4MjZ4
K+uwrdeOl1mW6/F6/7DxkZv0ZK64MNbLQaBCDSM76NsYy8rimUikXt0mb09VQXiMhIh094SaET4o
Bjn2dp9MQW+vnZybeXF5uopOifgiKNnFgP8OKJHUMHb4gEQy6dSl7BM1piELFJz1Uk007wSRXyk4
iLrvdLB9grm0k/tjp/URd0KIKnLnsbX+VUzzP4mFfv/YCpYzlMwk0YNWSxYbqP1GeoQlwZmPKTdk
2hmWjXYm6oC7YzogRHdlbS6LJWjvPd7/6Q2qUZIHjpPHC28ycQW0hTmd6CJv2gmi6DAjjtejevbR
g74XbDVZJFJO+DUSEvF+05nCvC6OFEoD4WCA/EUu9w9L+qWsclPVdG5ai8rKxJBUbchDcjSNcsL3
TYCbC6D9RGnC9iRAOg3TFfV3Isae9vB9vUzDFUoiA9ZgmyW36WS9fxmE4EQAazG6UlOCi29orGR/
kTq4QzQz4gJALRAkS6gkVmYY5NDJ2FthHG6MS/td6w18IDMpk+OZMoqPBBDYdPSL5QgU0CMFYOPy
qFm0Y8eEGqUaJOhg8MiCXEEwo6J6E1Nhf9dTrliQ4beUkU0Oq4qUtMZY3XQHch725GTnJsY1RoyV
qZM5L4kO6mKcsKSr8ReXCp8EyQtQzSCCSKh+ZUEJ9mGeIaMSxrkNdbznbRdHtJ5bhESDoS/pzqjR
uTqhsH2b2c8/0LZ/E6cSiEHVWWDaWI5M3ydtnJK2C+VyvU6goHL/UdKT64odpKsQt2lI4b7prWcB
Hv0dNimWM5tuj4KPo0YOfPyiLtOs7JSrv8UnIiaMEDqhq32odMl6CEMG6pvqgvoFmYRY4KT4WB7n
sc7/Q5DYxYDh0DWOc8ESxpFBIQKFU7Ul6rp16OXyybI/lUtMAZLXNHUKu73yXv6DlKH/fKpJKz8b
/+II4gQ4dBvmfWTX8RA5Rr66y2SyDlHr0LO95ebsEk9sp1SD5vKkMhI6xHhDtrhfDWLdiWvWAFvo
njaFokSc4WXJu/kvzyhfYmnE6ILRoxSg8rUAPfROnk0Z/kcZ6lpQtF7Gey+3OyeAof7fL/0vz6Zf
8sVPdNEK8KThOcKv5P2+33A/VTu3mn5Fhw8Ip4rgrduw0RHbStgSO6v0CxE4UN3YA3D2t0rwMsHr
lHXi3lOJtwZJ8ROnHpT3eN6X6tMvmItKRaJezp+BVMmSjPOx8rj0yK+82/GU3ptt56tqvVL2ZDta
X6xB//+Vj3KjyhJBnDKFxo7c+TXQWlNaCyxEy1/XpxEV8YnGoapCorMaQPCF7iOGB9JRUMPNYZ3E
egPpHDenqS7uI7m8htI3uOZDZU3Eq5D9YeFtU+gim5s01h1OH1wqdrYWvpil8MeOaqXVARvUvSUe
e9V2PHkHcDhuBWUKS5ZnDfOMy+YJMPPof/xNw6ccxTIdDCsLHvCt5LgHiVrnp3zmx9yRys+kKa4c
p3m1J3tCuaf0vRoHjCdO2bq1P8BOXLQae/2XhDd5nOJpNgGt0VhGKlJ81tXxyOWZdKxiVItQQChX
5PckEn7HYxKxrVeavI4ZmsddskdxdQaLfEgM51GfEejwvrLxuYPoGt5NjfuWE2sy73qKGIAgDvE9
VT8RNfvAyiE/uEdv11eKmu77zowgOb6LTVzuiDbbf9G4PwdljFvfXJbpRMuUM2buEPV8Q5X6WCPE
hze1ZPUpK0iXckHr/bKEbYaNtNbMl89l357ZSpJO1XyYcH1mAOUWM6pj9RjoRhc97tHUF+pGoE+6
VgY1kOdoIGqptXqg9vEnl/eZEFnXqeASR3k5Zl5n7g8OZ1y8ILZ9o3VX6d4oWtg0uj0e9SfEFWWC
AFS25VTIVoTkkuw3kV0/jvi+3XXVehi0mSjIMODIBCUmBHVKemAtijSnhdS365Mf+esIY0p2FMlM
zDILGmiXqLjT9Ik+Vu3ianwrUS0fqyvZkHN6MxEXDr/5byZv8BLhZHSe+Pw/QF1jj8JlLJ0LbMc2
Xo8xG3kukr+vnZyJKXs+ktsltva6Vi4Z2KmkjzoigQ0jl+2NC5KDcj5Fen8SZXDQBy7nAPKvwI6O
2yS6YqapRx1p2EdUGryrr4+G9QCg/Q9A2Ncype9pkH1+WRZnX/444nnzbdOZhV31KJOfq+C8bWe/
5YSX9nhDhtVUnp/kc7+WbsOD8B9bkFU7MzS3odXTAMqs7mNy2drVJtAt+5OguiQyRhYsTPI4iGsZ
zgBirmml5mvvZEw1UwbuysaYou4VCFXjzhN+9eo9z+dZrhyZwJlbg0QBrLW2UDM5meyuYELG6VUU
j9GFYiMx6iJZJLwrEdjtX54F8FWhPMUkuZWbzrZo9NF/8KQIkuWomRFBP17Rbg+1VMihXXEnU5IP
NCLlHpW8M9Xi+ol+aOYmbGobV+Enivvdj4AbmToXbOpbe8XC54QYtdn703mq+htw4XyIujzFmKOb
pPaR4kesaMjeBWg2TFuy90ni8LrMjjAQl7Vaasuhuwt/JFWwHutPawUf9rzqZiXeV1XLq9PXIHXA
n1En60IAcoanC+yBmN2Ne+OfeMgU8B5JEFSrfcmD8vCOU1l+aQlSbXYEPUuEF3hHINv83+05XuDn
a0nFdAkkUm4c2pfXM9vFKTRmKLLaT4srL8YzmeTs6s0JD0Gfgrfz96XgxheT1W2/wLLpMSZKxbEg
Op495sxH/xqCB7DAZN4yjWc313Dq8xR9qs7TWDLBqOAyDBHiTt2cuz/HVcpvZg/mKf9RLiBjH28R
hyp6petZZrSsjcD9DQKDOQtfyD8ycsFTXQPzZwEtUCqgjGQ/sa/JXyL3msoqH1bsB2FEBPvyC6+o
cZZHm6X7mrj3V9EI0btk0/eAPjbJwnUNgBi6QDFAsKDTOSQCXQy1lzyfzlLgJyOfl93RgDtzxxq4
A/MyJoIcAkmcsTu5MJPE4PuljxdJR63r0Umt1Va1Aq9pYf8weo5UbbIa6wxiSJ3aFp75eafcJNuv
4jYUgrz6A5ylb/ClUNNzq+Pvf6R/n2flkvPlksfLzSGu4FJ4iIHE4DZTz4RMCOixUG0RSLjYWck9
GD2FF/f9XKUTYzs2CllS+TnREGyO5DZvpxtuiShbFOajvM6qN5bxoyUO2VgZihL3Qs0F91IO/ph/
dkeBQpfJJcWacB6YX8F9zESleSL4Yx8DVTdtu6ZcjgewQxTwZgJagESatxdWOekm039f1PIvtZMZ
BPJDYTu6twLTBda3AoDk5SCvh1BoNRQrrrpbN8mamurSNr9CGmhISy5nDR+CW74nPqSQVxGYohjS
9fbdAN3Z2Wi55rAiphKUYQnt//+yA7dT3igOOfI1CxcMdNPEzKDmo8lN8btCkjTRqfoI1YO/F5r+
YDRGNhEtI8upAQp5QzEXxHwzoue1YskQ2lB6jRSo+R4C7sq+kQd8a6TJGrN7qMEalC31miVYbcOD
FbsZrNjMMsGAuYjkUamwQEFvSdBzYGoypvnk8gvt73sJdmbh2WsrPG7yHezr6OBb6jpcqs0XmOAG
suaVwIYFcc/3xkZX+v6I4DPQ1BpXYdzmrZUSPXqPdfPDkWUuGbZMTi1d1oL7L+dfkwaHrn1cpJG0
BWcGDSr/+aHsAGNodXJ/SDA9sUbaDy8NWkGK4WHwzPL/53v9LPZFur7n0ZeIbwG2rEKNPUXWpEH8
bALj16zXQn0DbTJBdcsrZoucJe9M/41YVUPhy3HWwAPORd0uVYClDEZ89qRT5NX2BVK8xhY2dWoj
w9cAv+5f83hO45jKZxcSf52dLIljw7hZdWNrQeCKlOHsdMkAYzniZK5U3XXSuRIh9TphBe8UmCrb
ZXNrWAZ2LWpKxoWA4tIjMxgC9tOqJSk5WAtvcjcab63I3Ld1ye03TgJT9eM8ti8Si8aOZJRRm0am
so2Z4llwilL5kme/bbfdKqy8wvEpkiUjCmMCAZ/fLwi3vhLOBMYmmAyTPpsd0UsQbfTViHgBWRaX
yP1rAU/BeO/zCNvsTU/+GxxIHSBWBl29wqzxvc2YM398Uehx93hSGwEpAVGGn5Wd/LeHqpozVXhY
pH/TO4vMhHoVLnmHOr2AdaJEAa8ul5xZm5Pp3e8QcSdx4z0SCT26IuSqXrBf+N+fqsr5a8SBgauL
jdgUNZYika65LhyIPr2dRlFmnXR+UdltvWAAnWKwIpX/x5FSGS0s2fW7HutKbcVwjC2DvvIsugsV
W4Eb8yk+g7WiWUsNprivRlJoQq8np9wLrbetQvgO3FYquR81kpekti6dPO24C/KEd4tp9XGmVAXM
0tir+B55XIzfrfFuL50BziQucpPr0y2TatY1Ha+QX/Spe0hdM0BLsRlzTwOZ47Yn2GzWYgpmZFrd
QNz3ZYFL7KoGT0L54sdhFFVlEWvErqWU60LJGnaDBq+/y5m6F5VqYhjEjoCeyE052FClNUbGfI2M
HqlcYzP35Mj9cRM2PrrV0o2GcPqnwdip/3kSQnBi+TLN0behtOcSd6/N0SSEr0uB0A6kw9ebuSFW
7xFUI0zIhvrztIpYnvig2NJh/FkCHrUTXbeE8jNYXAPt0RturbNp8MDZIXmA+CC3FSGA5iDaQRnx
ntxTNC2ZO2FfiWmuPuX7bTZ7iJ7Vcujd1BpPEpKg96E8ce8HDsge+yarr2wml8vErssuFvVDcBNY
E+DzWQWIAWV9dBW++J3NYnFC2gT2EOt58mENOusNzziRW/DneIR2hk6ydx+4UtF2KbJn+WXDL2yi
b/gqHHiqJqig7mQgAKsL9XY82b9QsE9nw11ttn1NY3CkRU+AXFpdYetqD2BBfUiD8i8qRFcQh88j
sjXvjdXOzRmiZ9LaugJxnBcdZL5vuOMluBB9CocznBO9kLUd7npZOqNPUNl1pOqsEcA9gS+qWmI5
+MjXANeIeC9P2N3cYw5pPephmLsxKS2Cc9Tz4I3ox7pyj5/yJbnJlizL+GoZwokBNHJsNJNsKRF5
AbwU7lroci7fV02nwBzI5qP2mXMp04oxUAhNDJZ6k8lW9yVSwvw85WkrWMCfkPQas+g26V2zo2qE
izZda7HxBoH6Q4ERXXLbbtKwINbTXe7OA3asBU5QjeilvLvjo2GrEr5JCxKQcvVbbCH21h1P6fMj
/+Amw6U/94DwgL8i+rBY+oqe/mRH60xocKrjMBIXj1dRiyAy7OE8fvPVXIqHyYoL6l6GHrSZXNj5
+lYjpKCTPJ785hax1n1pMWHameTEW4x6/iaQHOq0zyqAe4FqaWDZuAjcQChRyxvjH4zcf7U5Yqgp
bq5mGG30WDUdpi5PVLiTbUQo9KP4As1h2Ie3xw5lIl+DI+gpiMbSMZxCPacRd8C2E+5CQNrUMcms
4a80klBoI2NzIz9OKU1RYtUbtrh/8D6WSn8G+ug7hlQqeOCKQ3XL0ZH1UuWMrqjNiMomKyaLNkrI
+mqKn5fzEQwJBruMb0545kX9vA7KsTBtQBkd/ZgDbmZBduo9glXkWUal1vMyuD/biwoPM7e4K9bk
ISvFxnXUl4GC5xJ6icwWik7Ec0rB2P5DxjPS7LHNnhHL0dpbJa3X+gwwP1FP/US9UcbUwazi8DVT
gPsjABb7ZZ8ssFw3tVdMTxU/8TYODeQS6wWyeKxeLuJi6hv7IruDIc2ef4ER1NC9doMTUIdJX+Vu
Dt7Lwjb4Qw1Rs9f1ADBXo3MQUniJFbJNmFb8ViOMWoig6mWKLuhKrMZeTA1vqBmUdRCc4UMc012c
znYwGw/ZxkF/CWokwlw494rNd90Yb67gdKFRtB8w3wM/VINFZF8Oo5anzmAV7gJa7LJ+JUbmayyu
urXdPA6rMVLLIBLuroFrSyThJ9FnmwQvpKJJEsjM7xf4t92QuWDF4rKgg2pUT4ZNdMqh0nGB4lRk
JLdeEG1XhJyqjVQanR9lCpNGa+24bM5mQfh4lmNFG5jHqTYCuLrmzmxGmun2fuER5sx1R9ub9q2h
P/UqzRePa5/+Y1At45pow9boh5nY8nsa4SWESQ/BAuwV/p/qZn8ZevDDbu16KI1X44ThacgUIfz0
iMwXdN3BLUFshjUlpgMAGYMSzr4quKoUt7+IztALrHr+Vdxu8ytlY/LDObo9V3VM+d5OUNc2FvS7
MPgU+NQudQHtWewFcXH/iUk9FcvOeO/eTW3uFwS6FpVFic2LleoHjbx8RJiVaxUPbr9pRf5OouOa
afbFz72WOKtzVov28pOXD8GItUQ6VxK5ioOqkqfKsYZGrs90FNTvO4WqzcScqND3MT+9sc7gHpbe
0atMiDXImse1RY1fmp9Dw0d+IoeJNJP1JhzQIVuYojZqVHz2IaZwOWtdPztEjIDP/Vl7iM03F6gh
GxftIxVWmof0XgyDmcDtxP2Fie9864URVBxw62OiEAaMj52zzvAiDLiQlU2TwfXHVaR3TOP+z4la
zE8OZLqhVoASDoNR6ava5490efcWCD6Yges4tzs1DYoUlJeomjUuWPixiQdTmT3JQMUbvouGSOF/
PGuynzk8prYAklybiE39cEa+aZTaZsY8yiUCjM0I/BiXVh+oPECokCx76t5oajlymwzpczOi0+QA
/btAwlvhpwJxT3X2XEHINUkYW1AJ8xq2OaNSUcV/hBiM3MR40ph/mizFjdGsND+cfrzuW/gOWVg5
IKRmr5lTWRPPDTaTEjG0LBX1q3pdflJr5eSLw3OseHDQttj5L2WxUonDHaguiZHbM++0zNpC3glw
KWWIXkCOuHumiGil7Sy72WsOBT9jGYeIb2xcizDq/JdfAt1uZecd4rhvpiraUok6zAeTxtEkKDCB
+VHdM9f4l1hZrzSklmWRiVC7tbgUHiyedbIMKtpdv0Z+aVpwB9eYMQ+9GA7zpUtDUtslfhCOLdQi
Q7eU9mvOjzecoPJKwlT6/9fkPI5pdMUUG0SoDjpc2krXb4RIt60BON1wSBYxjUamcEDNlDNmJqpO
3/gzFKps6iqveJoZMRH7ATqKDFKlaeXueeaTIwbqehAPZyu0O9U15K4QJdPqx/6CDRLXyesXxjVO
T61ARnh2xSuVo+QrOWTDT3DfS6/d1vb8Qm3stTSidHlxI8+jdstTdSwQJdV9k/y4mmOe/GHaXkoR
ZMlu1RgB/5RrZg4wREKhnjACpAGStvl96IIpoDWi0p6/B/CRBCmJOxBvqnS16OQtZC4lC2ONoVjD
+kXtQqoj/t/uMLIFiRPLSMv5rO55NO0KAq02b27+4KJGjjJnahZkG6dBk3tpTBXBVTh/u++v7TCV
3om3kLETndPosHckFxhNB81LoJ6rw7f3vUNWtCfvB4t+bdSLL7thhR0vVSvSXoYkb0hRTPEIw1wF
aE3UhX9O+ohVuKRhzfu3qJJpYZwEc6b/dLv0emPtuBIteINdXzf375pZf7ZHAwCVYx0ST8ZvqJkc
Je2cM8Kw6puXHijIRNHZ8uaepeCmDDUFNVgc+G4w0EA89kmblDdrXWvsrv577CEhHKAUQ8w4ulPc
2PppQmxH/vt+QsKyGgCt3ngUcmHCKJ4FC1/VsjibMY6rUsgNa8FzCy+JfZI6XdyM/6eyoFEpbhUf
GiEcEen/mZ0PyOna+PHo0aCkdB1Y+YUu2JjvVXkgr/pMAXWQsrmiTwyK4O5viSaUVQuy3I3FOfeF
Zz5t1fFSocj9RNDIOLO9lSob2kUMEAl+E7sM5Bg1rlvJ2wqJQsBBOYxI/0rRYrk5Pnr8acyN4dKR
nyUg0xVI4jXd4yxpy/gcfgMimDsM75EhQpIp3VU9LEKczGeGVloXvB3rtzUQOoEHw7A5L1QGZRbn
39dB8IHklw48zw9hDzlT7I1pKHu4fcII7K02Ru0sTkAaElJx4G/CKG99bOMSM+0rOhY00hy/gUBV
frFw9h+Uxre2XeQgIjvifth6b5N1r0Y9oG6VplW2xFXr9xghwLg5OtcqICtqsSLqBiXvpJI7lVms
1V2nIVHbQmT2bKDAW7aL7gPLAYzPmu5rSpo2QVuXT64elhBlZkocJGtnHOLjXc4dFYPdgKjXAvs2
mGxXdZrHN9UKk4JX6XbVux8LDDPO2GjYxlXB8LiPla92PM+v3tj+jNp09iD6W57W8lhqCWZc+MwN
BJfl4jYLTsaoUKQktr6MRkCoT/sA8qu5fICtK4YKb/6oZBaYF0P1peN+wSv9zb+Ki8xM7dFLRoRl
GrJBznpI+Xa5eweZ6hEVeWVuKZCo93RC51L2LtWlar5obgMuTxdaE3d2bE8BIpy0YgQGdfn2T3N5
cw6CXsdgntjt5Mw5ufa0NETSeZ1Kg02c+nMt+5K7InwSOJAK0vaUTD8Gh4TLUlopk6m2d1hoGJKD
/rhgE2fMD7zpUZz+zryqlIICSQJSe8y5R4YZ8Z3SUyc/lY207Q2VQt+fABGIP1CBdC+xD3WLNvvW
NpqD2mP9LaBvovRKQHWtUY9PQ6DZ8JErVjcBGVWtZwU9bzqAHJS7sCYVxzvni5xRWorSYHhZLcx7
jnnueXR7uYi4YIW6DqzzXaiUYHptsQ+m7EJ+MukTs9Nr1YA3aaupnzY8lEabDNZRPsIonN9GkSt7
XMr5xFZ90zVV6IwvWIOT/w/BIMXFeQup/msS0Fa2xOuiW6ckhPBQNzdlAcgflMS5yMOTws7p1cK7
bY0RSOF8RPuR6xriRP5Y+8OTWh2KMLWLMSH9ZNO8L3NfTSnxC5MtNUijawS1J1fbNpZRb9hQlj4M
MMCvLK+DphFYloa1cgeNcse2HsU1jgQZO34B4rjgRglZRLxyDZr4DeRi7KAWxj4h5AIIxf9IPXgi
UQXcgQIHIbsmxCopGIkGKB17e//bgcLgMn48PMJPSmOWKAnxBAaCQ5u4/KN3n8I61Ssx+Dcx9Zcn
QJ05GiboiRIjOUgvnhGJ13QvPu+S+1S0+cXdHOhB+v5Byx8PLJHhFz7bvdT3bfvniL16btM1xwh6
zL4KnqolZH7Mh0+eO+D7iri3RgT8JGD4zo6wNcvXAsbKZOmjagwFCthP3/BNejnRIjhsphfThW99
uzh2o/X22IhMZtNfNTf+0AhekatgS4cj0eS8KB3EZAqVo9NvSNXB7Qv5YjpqZGoZiQ2SiWctQdI0
BUGCEGZ6i/JHTA7+ReZA+sUsjlt05QrSCZjEPHd0OZq2VO8f7eQvsCjjSayovkVSSeuNyypu+XCO
jo+aeouw9BznEGcR+czk4aKI430foHcnwtw/a5UF9g4GDCKV5N5UTYkiNQSJxAbnx2T+MkvaAQWy
jwC5tuq/JQh+5jv3MdwRLZMIHvnXw6QJObtWWv4pybPHJeTX/qf2zTuMUAsHmroWDnNHjBmNJsd7
sxcfzTO6/4WsZx6BEgkS++w05IczkeHQHD9uA6TNS4m2YamS7ayACkGfhDWsyzP3bvgrk/zzZLeJ
vgu6hu5ORy36BDBlTOBkp7X9IVM399ZNcUpDlXiWfHANjYV25P5XXacSZIWJL/eKOpuYn65DTV5u
nQJ0oAt5ndaQZbPs/LEXpuOCzcW8e8PfXcBWRbWumVKAxoScQsOF/DHT93Z+4zYGR2gJnuzuecSA
DjOngMh21/qakZ3UOfGls+oAE4bZYwV2WpItP6Bbf+s6MID2aV7f+h2Ndw1xZ+PlDMOeaBnLxYgl
eQrSY/kCm53mDt4IVLtgwQWP02N0zwspTSZMDRFhVlbirSZaYVSbLz6i7E1cgdtfKXQlC9WGIM4j
TU8jyLHqew8mllizEqph11AcDah+c6xaemVp0d3tUr/N909AtfhzwTjv0oAbxhUNMQvQI3b8+UTc
qEjcYqnq3vpjGOgFdvofOxGNjI9ag+1GkDbykzsxuDB/wqXOflQDUGYpmVm/WXzA8fvyPakYAdSl
HgKJn9CcaRpdosoeqvg9lEvCK+TtmrGb1HGKx1Voa9lGgGKTw3vxYadKeWgkBHd1VjMWHhV4etxw
sx3v+PuiDcKF3lSSexAhI1V3ztSpWE5jfAQbjPPivuiIeDO+eDFSfPLZIg14EENwsgk4KWfAUN+6
AEb+1BOiRE7DXb/KB3uMKlEzTMG9E6QC6XeKL1lGV1Ji0umvzlQyoaXRGOiwtTVG97mMxN5hEGcm
tL/6tlREn2C1bDA8AZCQikFvXn0lDhvWC4sRNzKaygGjqZxpoXTRVuPUQOoZiy/KdGz+QsuFrpJi
ZjEUEJpygJDH7mIis5sQ2Qcsuac1ghIAyl7WYI5vFVmNmgIfXmyghVDu9oKFAVf1XqERkLuwP5Qf
HtJeaPsq4Ty2og/9n0qFmKTfYc0jmxE6QOzkHlfgje2P5eDuDxhv/e07lffwm92rt/1qd2gB4CZQ
Y1Up3dwrYuq5Yhg4hDm9ZipSsh+NrpSKS6rAp3JWuDeYhunnJaESz1Acb6yXQx444Mb2PA88Xkkf
AYmDjQ9EV0wiOXEBpaVDRXYnWh1fz8jVNuwiRg68WezdJPcAAc6CmmQxX1BBCydZYOS+WJANXQcp
96U5ClGHh8/iBJkXWTBF7ZzC7/1APMtH/G5BkiL9ytxCoKhgHb6ofFGjHbRgbSwt2cUd832ZnJSh
DqGs+mwpqDwDRtiQq36OLfESu2tDaWmBS+Az8a9LZ18pyQ3k49HIlZMCxSnsoaBH5z3XMBSS6+jK
vAm/LeBrfAZVZYij3lxcXJL2CrZ1OGxd6qXl1734NGmUkFQYPIScflBcpw0Czy+OVXY/fyCsnxAD
LQhIfJOGkJM+o3C0NC9HZG7u9iRH8Ad2OFjjGbv7D1bOCCc9z0a4j97keBNJE9B8DFRa+xPDUHqa
I/C8xrcM/fAeFi0CIMRkbg437leOoKdZxAdMIfd0oWVbzZH6w/rj33WGDju/Y7Iv5UOJ0fVnnXjM
KWjDDqUa3vSfdqTB/NHsFEZM4gi6U0PONDuLQwp8BQajukkxv+ZwLV+K0hlE7/7jL3pqcVqLwwsJ
RRwXfYQ1HMC8SM6NkPSLSxXwwAwyPKnKdn3d/MOHLRPOw9aOtYNOOyP3/HiAB9DqdtmqfYUYS1+T
PCkgK3br19/yk0TaXDxn4tMyY1eAuPjcZlaheA7Dz20Y+7FCjarTTERj+gdELx+fFyQtcr4REP0D
2Ua/KyBvTIpDLgyA8sG8BXzFqR+AJZTwqAEG2FOPJOxSL81jXixWCUHQha0vebeSxkTmATHYiHHM
PIKifGF824h5rliLH+f+Lig0KnNunh+Z/g5iVpBTSWRjW2Dol3y1mTg6KvlddBRSm8jEnsmDyG1j
WF/lDIg7co3uxYbFX7hYctq4/pJWpP99pXP6QKOQk45MnS4Ust6I4ggRcfVyuMOA1NoIAK8gUfQF
/zalkpkJvoCb8tyYkizBz9aAqifSl1MF+58YFTNQbDMBKLfDDnlg+mDEiIV9PifpBjc4gFFFoVwI
0gt0OKK306RiCa/82Ve8+8VjadwmqyiXnXOgQ+RsC97ZNxt1LgyKlams1RWBBx/po/JE0oQVI+L9
2TfwKpoxobWTFLikfz9xbzpFqnc49hi1C5THxWrq3Wz0B5SIJNUFQko4jhCzILj4sAUjglgM/7DN
JStmV6fmJd3ul/qHOH+g0CwkBypZA90Q/D63Y+EwhjVhaPmWKnPiIjKtbOdDKOdCDMFAnW9YqGq9
ioA1y+X2THl6eMdpr8gqkTIS6SAa/iNQBKI/G1EEwxAanYtMTBgqur49njoQsXTSzxs+w+Rgl7Aj
lnUgfxVRvehzqb4McYgRrTvRpcfWDLPYNMByLeBhe+FR2U0ppyTiitN5D2lEoUhGxTivlR1WLMXZ
HqQM8t9G9hZY3SCZxMyR7G159A9QBNRpodnqHKnft6cZF2WxG4fYhQWaGWBI/UCYsQBoWueNy8qF
Je/YTKxaIjMHcYLHkbC5QDApuPJvHW57etmfWH+c1xDfnL8FUEYQeL5U4PBYqod9Qa+uz7pO3jod
JVpy77DHzMC6JaWo0B3gnBnf1NQfTGmEdX4pxujRO1YY8Z57mFItmWmiLTxtyszqQJQJVzuvON1d
DnMPAyHvKP+g3SEgDhwSw8EZsRFeB0vixVsK3i5BXZc0e09Us8HXj8+XNqtVRdzA6JKld5rIoWc1
OC2C7KwpUf3jLLmEUMK4RHjrdU240xX26Va1Cs0FZQ9fm51T4RU11g8tUGxDVMi/i4SAHI5C9DlV
WQkawbO8wfVCeUfnxxg0ACi/UdePUe3YyNgVm6w6gSxIGP+3q84ngKKsZrHZwRMyAJu0tPBiTGaB
YNkiGA58HO58IiXpCyxKOIyuW7qpnp1Or6fGvS5914wtIj7xubGpvLyo9c2lYKSHNRbqvM4VVQJR
jcoW5DX8CoVjSv2PC4CZWc2Lj3XuWvHkcgfJlXQtwBr3eLJMjoP+xgjrRw5cKpByO5h7ZF7v0E5K
sQphnN/gKdxiVTV1dFqzZneM3BgLj+sR7QtupAJPczOM5vGShp4zWzJKkHaok8TaBWAKcSwKSm7F
LzG0Ip8maNOy/qA6xh3lgO7Z76ETIdIPiyxCh2ENN5Due5JishFfQ7nhMFSUUymZHLJXBPCDNox0
GTu4g8X01Rmi+Onz7g8V4/ffhogj0YdNRewfmxiAsdbd6u5ARSqBmZXTFM3u4JjxCh1LpvPsFpUx
LD9t4JJaK/8kUY/4vKC3oIDqwsmiYFxS5PEWQDB5mHXi73tLBSdlwDJypBpyhtiaxqS3wHpHeJ4u
0s7sQb3bKFH80QMUFAmSy7sQDb0TOZRygJskUpfWP0IByPo24tKSUZVXFO3KkI7CL1DlFYk0dWiC
C62y/3RhkHNCQ2ksd2vLlh0X0n8tmg9ZSVO+9aqdPxz210KLGd9vzk/BjUL49fEAB1ivVfSN6rBD
H4N3YVlHPJJu0XFGMR5KFKgVc5BJIiBspUuuYNSMzUZBJqR0ALO/KSQIIpv26PbMCBon4KlDKPsT
fWD6P2Ztr5bxDEhiHnBGOzIJPYq7vIZFOGLnQSHvqCqSprVzrk+ZdvSstXmgc+RhrCEEqxsjAaK6
BdvZxOxkoN0X4ci+V5qSVE5SudoD62GpcXIzLXe8cyi0oFQ33rZVEtTe7Htm/W55RI3x2nOPS7ij
ixrwsMq+mMmDV8AYvh+NNuQWZLR6SVB0Na6RNMxLyeXzdXsqEzpbW+vxivXCJ8Mxh9XMprrxSGD1
NdVgKeslbHN8H9kj523e4jgBuI8sXxvDiRKJDAgQddecxP8gih13pee8+HtVtSH3/ZVpwy8u0z4f
wPTJuV8PpIe/9n9XPnrc85szL1U9mXRsa3hhEGLj9+vK+mWcfAOXx6L3APpijpcGErWZyPf1XQM5
UXMXp8zndV6eiz0FRSstgIF1PQ87V45aQ/e7PD7cbf/qwOBr0bpZR/JJ7DYLmvjbjBgDBUOf67y+
8nVL6WVLuy2E3W4zTeyOfRfTVvOnITQz3xtO36nknvPRYeu6IqChNAQCe5CmrDbDqjtgcWnCv6ss
b9R2G2Ud/YHR2uaP6apWumZC8dEGyVFqOo4llpeGRkygN3FbcuI4adtoO2QpA5v5CvZK68i393sB
b8GMSjvfJQx4uNq4BJF3PqgN5A7rY+D2dphmXQzK3QyHk7qqWCBpiixpmA4IifhaAsQpGoYaF0ox
omnIvJkvp2UXAkjy8ZP4fa3jugXjzIWguvadrCQrOY2s58WKPTL9gtwhToI9Py/FU4SW1vgVO5Qo
LjLMFWfU/CPVYcnNSjE4OKCjBo+zuNFjg7uMk0nzsqD1wNwt+ASlQkk9oUqEPkxRQc2XTQYKUork
ZF7MJmjNCp1P5MrHmD2xnIcnURcyUyGJh1He1AJNZymh6XbNhaLr8i3dTuwydJ6mPzI4GZwz8jKB
7AEXaY2xRPdLaBNZxETLJ8zEAUNxXyEdhEjqcWRxlQN5UX+We07yX5sS2tmdX2j+ekkfSMR96mr6
nKItJQmUmDRCvqOJ/J/adaSEziQsB84Zq10n3pDsG2l22TP9Of0b3JzRPGVs4mqPM4vE1/8Gpz89
KFGn8rN38KTtEB9jUm8qQ2LTZvSpmtSUDNrNuj32oUKJZI3pvVyf37vvaGx/LwPQZM35wH8GFQkV
jtJRt0xeMYJfPE/YdZOcbMcDb692VMXmeKPjEar1A117gnw4lth5HOpY+tkIIt1IWC1hey2Hvgqw
lBDLPKuzz/Fs1XSwTISU3NfyCV8nYbwj0Z3ohpRcfo2Yykns0gS0Dq1uK3RerovwLk4VeADacsB3
fRm5LACaV42C8Qrub6IyU8bTcvJH00GD1dwXB30DT4cArzf4gsoUVejt53vnAWKAX6T2Fg4ptCFd
h+opf1g1CUtSaql+9dbbR7yXvoExDso+m0vjQFNUC2gZdFV2bvFjnzGGokeQpnz8iSsuuz+FuXY9
fYSdqj8eWn6PHz7U5rpKCE/TM0olVjRfqZFOlWoqtCFftlc+SM6lCnZa1Bjl3R7n5hjZm8SlOoyo
c4FJMlML6ssT5BYA9R1+XAMwb24nQZu5bGss0YdQ2z096MHDRvmnjhxTITVtpFPON6XWt5uPyU1y
BB5nQERSiYhcAZ2JKlaQ8zEfyfilkTlJzsEYCiTkfM9946CGNHdit6JfyxKYlDZYR8gN649RYDBY
C8fl62ubgW1ZQUTC8Z19p7pizlK9mhBQtBf1YNNRZoCAwSWDvDLUhzmILUvR4X4aTfzG7zgJzCpW
O02XMakxJ35PXfSvBR1L1KkCG5p5pPiZr7U8vJlVHfICxbbbrtKOWsllSSj3+fCw9kZZ9cE5yM2x
hPXSzPY49YhcEkZWErw+waQZsmLOc9XMcMoWJeUNAeot1+66vfzRiKKQ7jxE3pk6JknGDkpwmGLa
fal+D0KE3fxAb2gBhITlkX3JdCKWRImrekQIXE9rh9RTRFtbxpNilzA3JHdNYZZ6B6/qoksWgZi0
+xIhXVZrT5FH270V3I6Bx7bt7dX11+RA9UVuKtFxjc0cF4N7M8qWMO2ugB56gLTk/qq8EwDhPN/o
BAjTnfIjzW3I2OAvdVHSb+8BpXboeLmiOIQ0NyglkkDpua2opCDOqL+GZCMIBkCrV5Ngwr2yx6yI
BTCLW+QE8Xf6taYwSEqHZKYFwgt70pI8rftOfpFuoXWhOUmpynMnV5bqGs9QyIfZHAgg7/JlZJKD
BDHZoym4FvMUga7nuew9VIppAeT14sFSVlSDASwIH2ie/xCoz4FiJPQa85lqSIFcrUKjvLIk7GTk
Zdu0jNZRPAkdxQzP38aqRa4Z59u5QpVRirYJyhyNNJ2MjpV6/ABx1zVIbjDIjS7ZIFJf+kUqwQff
g2l5tu+KAZM9kxPSYiL2pfODPTQvhsY/my190KniAmBudNvdGTgrbzDzZaafneuh0amG61yOI6cZ
shcA4aJLmW2Cy5Gs1rQVczKMm1CzizIoIL9vigz+sUerqvMBbd6nazQ0EbVrPlFnyNPw//Nm5gog
Q6IepElS3sXvKP9AbhGl6w7AdPBOj1ZQK2MW1+ZmRBtvvg8jUHyI9kNKirkBCR69IWERz45XZIvv
atDKGDVqWL08VQ4yyiTOPQ/LLasCqHn1SPkoaSChR73rC37Gv+bKAKM2DkV3MFklelhZtQmKiMb1
7xvWiHFJClMV55PLrd1aVlqT66xsKCXFs56rlgPcuEnHit3vaN4U2o1ad0hmxz2p82FyiuU4fWbO
13JgMqMOc/USMxQo13A2YvYGrwa1n5NOIgcPRI5nIy0Pwb5K856gJwl0WYBaBqNRSPM4UBrLQHSi
+ykqDkVBS8czpm1ecr9jbOF3uOQlE0tNrblKYdYF9pvb9IQKLy7M4KEYOykb2iOarQ2XkqNb5Ep8
hPUTxcwLkwDVxxDsxZ16CTZjsM1Vou8fi0PqzItVAc9Dm8mLPZDybImqRPVlRchMYDDoDJMgtXBF
6b4LA1/hkmxa+36qETaa8cIqP/oL6MfQGyeofxxVHkcnZFDXc3oKkbb+R8fNiurVlhYt4rIMErdr
cpjAPYVcvCVrIYWd7TOHkOaqBzldn7TGX4FKtg+MV5o+QFt0cN1YJgDIgPeoHzZRCDMnYM/Xv4oJ
aVpjE5w3cUeh9zYoKY7o1Tra11o8nkz8SXcQen14/ceKLFL1Qnmb+tHbBN2Ir6pll3U4+OMuwfaZ
S0B5wM+CRV0EjGf5fKs3+k7Th/A30DDopBQ4IOY/qmQ0IL82oUg9VJNA+3U+fWvMYi1lqnb1LmKE
xgy+FXTWyPtucvxP2QXWrja0LiF6cDqvRjY60tcoWyTedIfbDqdS5N8I4JjahQlKTi5oTPu+DRdx
PDZkSRIFcFCgW88SWPz/5m1ata/Teyhq82zRc8O+xefYWSmuM6juETLhGAoqeR9q/YunX5bCS+Np
uH5yae1Rn16c6FEyikTSTXiUwPwk80KfBDp/VWuO9lzFQcDkVmNOtYok6p7MXIhyUiRX2p3AAnZ3
/nk6KNL6AZ6enQVkkIydLGTv1lmGxWi86/snAMBGOkEghNxXLF/zd/GIEbB8PHP8YZAHrX1/ur8V
4zfqMAa92Jpp/pYn/c5n6UnnEcRJ0BrYbILTNl4MzXNtDsABlVppizLTuuB98nMA5LqpXyKFpJls
mWm6vZUHGEaCMrACoGWH/4H7Xj8WPGpHY6L5BIeDYMXIDB8bhGjCkhvIviEzyJLZQDZCQAS0eAw2
PIk+Y6fnkmadXNw77Uv6GapVs48TBb7MqqLudnJIh/SsoPSMtHmZo20qs8McUrz8jUUSXWZzsU7S
4XlchTjvDxYn0LzXR0xo2eK5owt4plkgAZJZgUuh5vAU5O6MGrD7FiIhX7LT3ncteNp0oTkj6iB0
m/yQeRklB3nNqVigxVYsE0qsTg/TlVUSZr06eDZBSAhtB0sMhLIfDgQXWqZZtfG0PnXftH7Y2uQ5
7I2mKGi1gF6heixdR3Y/TNnOqJH79X6sKEFcYLNTroYrwKMaqRPxnJxg1nfnbYEc7xe8gMHwSWeF
lmAl1JAuzL22nKhHvy71R/6X2mBw/SjrzwMo/0QomGioiCm8/en3+cIYzYVbuHn1bhyH94vl0Oll
TO11CIW8I2E1TaYbmNpvXpEn5zEhjjBDOhYs52eH8mspROos+9Rz3/LGxViTiMrcGIlQYAK4IypZ
rEcpZE1/4nPJcRZHZIsXcTbDuJ+x9sxbQEtehPCSmvE3Vn5Vb8wghrSsP+W1gFvbVmkkLyaBK/hH
Gz6Suib5WM8UvAsU+trzG116+PGK2+u5knjSNJlf4TOXSo5tiv+4Qx2FC4KhgW9XXXvIkynlx1Dp
N55YhoCoA1el6SRUIEPz6rn4/G4+iSGYm/SIHKszRZ7KWvbXiQf7TD4yjaZpPoxgAw62NuvETBSS
qMY/RGzp+ipowU4CC6uSnQ9IGwaJPAO338hkWUIGDGQ/szjt+hR3K2+2TQyv74yjBS7ILLExF9+9
tK1gWnxU1eRx/bOYfO/f+AxZvq65rTGhO1URaIRghkmVaMDaDGo5JFQeoCEmlHhMev4DYag4tbLn
OGXVK+DBdlefwQ9GvyDxqusiaYaeqdymMlzjbG1a3uR7c6Eot/mt7gLcItxVUi9XP4gU62XEylbz
wI2Hzuf+t29YqPf5EFSmWX5JOfB8wd1bHJTLk3zEfBG1fpxI6Cz3QIAbP7dQ1FQ+FxZCACDMiemR
Y2CzP+atCSy2jpEfRTMrpC5sBeii9P3nNsKEGac9LblajVPlivcU5Qdk461edZxpsU8eYgQdG8Nd
1bBwNAuDDZWoIZs/wvAE2H//5lP6yrl3cRyPFOgAD3Habq3OzoJRnlo8ug4ZNBqjGehLS+CPCT8z
7yATR26wPUEIuseA/Y0sDjH3dqiBigPfQVQ+WcoNUcSzkbfmaorSX6FyjM4IjcJsW7xDwQghXuWQ
rhZ/a0fdcNQiCf6gUYAc2c+A+neWUWqBF/SbNw3YEwNHEOg5gQ+xj3FlO8uF0hsIS/jG6MEZA/RB
QV1fm63evRidB/X/DGC50oCb/9ezzhMATxoqp5U5a8UhjHAmkOCENMJ0buCEal+598qH5HOrw0w8
yE7tpQ9MXl0C3qJwE0wIr3dTZ5A9ubxej0mQybnaBfJr0Rgv7wJ0WbOo7kbSh57+9m3zoiaNyIV6
XfERmjM9b/DHAUE3cJZyW1nmI8l94eumuCyD6z5bWQCztZNYTfOgzz2Gj2qtEspFOL4vH31Igfx2
ySeic90mWi2N315pw3tuklnrHr9e6GXg8dpfqo8sICMjIURkUlyyM5pM8bLJqJiytuh1q9T2f/E3
lcpgKSUdT27h/UJlEKyWfVcqsXAnJuZbTMbrlD0pgULhPmSnKfrpT668K+KSyyr7Lh8hoXb14Z0s
nl4Zeh29vCotYu+ii6RWu/B89mIB94nZngh1H2nZGv4BTW9jf/XKi//gTRdggwTVwkbOwuZvJ0pc
4eaPYjbzssF7aQ/pL5BtxDwlW8vHYnrVDbFtkPAwdH2Yx1Diz9Gsk/4tdkXKOgRat2YwMjsLOl8b
Bv17VBfOeYxzkE3AoHl7SPjNZswHmz7X1a8mFzftc2peAMmbcQ9qAD1vqE0bQGdsP6i1YZXxM4Jl
hrD2wTCc3sYADII7bL8G0n0CsOket3PvGaiCcMXIBHh21vcBZQXgZdTqZfVSeuX8O7LuGFIgnf0x
xKH/HwmTpc9ofuzUEEohE3thV7bBRMIhK+2yHwJlitRxPrKoAlpy5gWAMINJ6qdWYtvScK0hUxok
nxCKxildFmuUWij5X4giu9+EKdf8cStABF3z3rmPv6HvQhXXJOSifZ1ZXR500UsnM1n7lk7ah+Jb
j1C1/A0CZpRHVCA4yded1ykbRp15BL6TB90SqMrHmX/FoLnhWlb7YkSljW5DQ564gjU1c44+WOtK
+g8ddN3RVp3roAtkABMquRPve7ms5ZlGTyVBS4l8tGuLSaktU1WIspiKQol6QUHJUc4SktggAs+o
sVf4cg2WMDr90bAWJQn5O1S6ogShiKTXoBrKx/F+Rs2zeWUqogOYYbUNFwh1uZdNQPgGJFM7M/XS
gQ9IUN7Px2PXuHco+1DYBCLH0ZktZuKlHrJrkAOxx19e+WfJ8cw88z0YzuJI1j8mHoNjKLGoe1SR
mfp4y67Cw3oYRJkFQdr+bowkh2Wo0I5EeL6jEs2+jPPwoOPDdK40hSg9oEaNVC8rOFamHasnewoe
cbSqcVgXGmGUziyuNnAmTsLq10y5tJ4fcigGtqlUJxhuGvhMj1hgQOFCF1H4j2w9j4yAzd42mjXO
hel/wTy2eCgT/IHn3B7AUbfYrYQQS9cgczGjJxd5/pPhJQaMY5zLCjmG2Uxd53dl8d1+dIU6wl5s
DTxeCqk/ZGfhnbRwkTk7s57IzQSWaertnzcm1a2/Tv8dLWFnKzbL6gZLKHKmO2LslnbBcoKvH9rP
qFtJ90VbxVYkkwJCO6JHOvuDMix8qmjrhKYAY7y1a+9BcohRnPtgGyBN5xjWTIRvl+d3U1gWUcVE
1IfIbh4wrNxMnGXIqh6xuKfOPkqlE/qCUtTaTNYbhY/CHWb1FdVExoIIcWNxqNCN3TIppPt8n9Sw
TKUn2Vu74uZQqCtTjHzBlQ8lbP7M7yHE5TdFpAsR4AWygKcz6C5bpKaXmzoPgiV6PIX2huD8vLke
dYtEkPuUypueUvgZFFn8oPrb2aQyrG4etUK2LmFBNc8wz9ZdCye7KmWNdK8Bo1Wp87F+qSh+kKzb
sWaQGylz+NDEZhOLUUlEL2YWABJEWMh81FZ0cTbi40JxHQAqtfbpizWoVm8YzQY3E4j3mQ2N8YkZ
mFKPbjU2FWbPYA6KKlmcFA7sDAeLCYDjxZJBXuiz2rUrEDQVKBkAjW5i0Rjnxq+ROnwkmfewwqhs
RTfb4XnX3+2bE+O9OXWBt8k3PvzxkskctRuu81nFv4I/g6KJtDZa0tV7ULMw4vyoMPdZFu5S3F/i
9VMCy9xtVXDgUiyad8j6qYVDCWh+YEAJC4x7JMeqXWuUzf9lwbP9LtJfwgrm4FRVu/9Kb792fY/Z
GImEACSCcfqtbZ8ZWJ4uwgvM86wCS3XlX4kJV1LyzR4p+ETK5C6lB2zpZZOtmujYP1gsgV+Uw557
0TI2JONhnAcZOzB2IWWC5hHLoITc5bGochIi5EL9uC6U8bTNNUQyfxkcJp6Ukk7XXEsGdVa+RwH3
ET+TpMGaVIA+TarMoj1MTT9fCLE2pzCaaT25fI9tSwACdjcpYAvnkWIEv5eHZH/M/z6ttcfsgIOz
+PvMkZrC3G/UmfsBdQNmHHDixSl7czmrz8mOULLj6R/P2Z129ODy1nke3j4uEB72ltBvCCYgOx/2
qDK10NKc4Bav7EW9WRHRFnEIo4mDRcZcAoQoxiYGzA5EAsRBQeAhgdst1ff640fqEMrJzVrHV9Rf
mHW3xpuHY/gJkVhUrgbhrk9lSjid47c71t8myUrypvznhIkrdY+KchiGZnadeKaTK2I3DMiXiDfF
Ec3A6fZhREUxYXdPtaJO3avBX3m9/+aEANN5Zrtpti+3vR2Ic8aqH72oS1+234Civ1vH3zAzeLPh
6tNKlpYqSVkANS9+2zzXFxyHz3hZNg3eeRjt2tl1gx8GZzAQ9TNtlYIxNzGcgHhkqm2hNI9uf5jr
PJJiiWsSPjBQCJgTKIke/dNpExqJv4XSj7qrmQYPKQiI6Bin7alrvK6FJMoFoZiHURWlbEDlfnEa
hK12GQQYCC0W+SSPasasp2y/nzE4AP7uRsneKYbB+kAoa2az5j0FMn3hjjfXL0ZvcdTPjk6thukA
+tGrqTerh0DC2MHAKRxOzphMekDrlkWwUO/5/cGCgA3a7Op2LRoTs/+rJYmUhErjUhv12UE6tcKp
9rbaRXfAuVyI03kzKZsB2KBmylQzgqpBlgF339yrfAi7I+TOcevsBr1Sl00Jf5PGyh4Lp+Fzu+BQ
mRT+Rc7k74lkaGXGqm6Gkx01zPwR6g5hg75pVFpr5vIoevPsjUvozht6xShwYhYbij5CgevULxaG
sr4Cwt/b67Uyz5VtL1eOO8Xk/Vp61ONRf0eadIY/6u1YnTmNR6cAij6x6Z4Ka3o5i4J/yOmNxaOS
9+BchZSxdLEply87u5Mo6PpV7rbTpDW9aeBgopeYC2mZx1QMDNuQi3klyrMWKMGskD2H9WEMBxSr
teGE5XWtxY66Bw/oL4OGkjxu67qKwb40e3s6DLLXqTk6E1EZGSxOnfCSBOVLqtU84qxOR5CG092+
DEsmxH5cGMN6quFBF4tHRNH3PQQ3WNtcUvct0/r+f+R6zsL3rT3PcoBIdMLfq9DHq1/w8nBx0sha
jEjHeo7S8z4GKevx8cw9DcbKF9z+y/jbF5Z6S6IY4JB+FyWwlWVX2k+1QRpu33XFfHbcBxLhv5v4
uUbmRd3YvmJkK/xPzCXIWE3Xz/CQO9ACeXuoZbsNyWq375GnBjty/WTjzJaYx4qHcUObxGWApzxI
G6BXGS452ijUT0SsUWr788hmTFZFEAJvPFd/rBBKi0jmR2Vz5gCnHJImsFoC3ln02U0nLAkP4cD/
g7MRREHtX4u8M5L2YYCAHzb68+28xoCS/uJl8B4fCQXH1+313M3ahK82gZcJrsbQEPGY4DYtIeuL
RWz0uGvDO0+BGlCVlqq4iBBnR3POZcYh7C5X4eHt1aCjehKhb4nCx1u7o9XewbzD47AJm2WhjMRh
i5PnlYcZkR0uFXUFQDho54selvRdg8qLpkQd77baN3/edOxCXLAutUStlJA/Pgiqx90Vstlz3NeI
6ntBWO3yEnjv3E+1hIP0pI4FdtyJ6E4EuolfXoD6c2u+BbQEcbPgZGzkL8Ca2Aah+Tt5s4pAuiCM
rkA7JbEWthXGl6/Ib0KKdByu0k5oa7jbr78m2txx+MOqYwzQE5OQhgIFxlh6xplYwbNZ8vILGlNH
h22o2xwGqy7cPfGvXO6ZV/O1ZGxjy2vwIp9osc/7epIbWBpBwcM8figFY59oITzhk+bqN/4yTYFL
XDCuXkV6c6wHBxqy2APr5g+aCBKorDd41VU9jLg4iTUFSDekc/MYKKX0GmuUCev3LwLokSODX7FR
28khkPZ0Mxx50GzuNpd1wozE20p0xejH513qHGeX00Ogx1fjel+/A6gYSXxjlqgX0SSX5jPTrgRY
IXgynLQqGjX1goYX+dErWZrfbvsXlvxk8yEtu2V1B/zEFQiWTpJ3a1vsj96JybhlzNODEHbnVE2r
7YB2PoQ9OMKO9qVZOuvbWoYa/D30xpkn+rYcGjuzlqPGXR5SZ7X0g6dx0igRAa+fBwlqOl9c+GoZ
p8Psjb8dALhlDp+gwklOj8pEXJoFypJGdtsii5xq/PkFlC+Omfhgya+E38pHAfPJQL46RjBGhCPB
qMavCr3WUZMNMZbCB41IwjuPqbtgP8qHm2MR4NAb6VzCNqUlomhF0tek+lKFx7lWYNRM9+rzPKIj
d5i1izRl7mFN8oe5gy0kPFGglOPikiQvXK/nBAxSnFK+IMoZXZYAgd7k2xi6bWz5IvPPyyB+aukn
x7GHugNUYIG8beb4N27wrTO9oZAb9+KFHbtfXE6WtXg09ui25KVKhY0T3FMMPgrOXPBjpw6mDFtR
zoEbPXknwo8ohKwCp4H4UNstu/NsW2yTGhuxExrh/rGdhU0acAmwhFivqAzjp1urlmymC6rh85hd
EsDIC1BqzY/lwohsSqmA1HWVPMFw/4j5Hm6reb33fUv2F/N2Pqg42Ful/NoOOGqcNsi6jXb1xJmM
N1ISlBtsfdpU6vop0EPqst+TsgAw5PbB9yfQ2RuZ0PjN8NLHYUY+cDzd04RCwIuTvZTmLDo8S+Za
C66AFH+EQY/RLisUfSHEEJL7GJjOtQyK3ewtDMwBxyVjo9822FGjQsgsnO2JjVAjvsOE7kYqHDm+
C9ZSC1/KUKhLa/x/f0cqfhjwxqxDS2WzbpB6B5TfExwmGfMzdOdSs5q7lPlcWvoFuEiUZhYlLQzm
TTBjGFbeOlPFr+p/s7EQkkxYdsOklWEp2XNSVeIAVEtyD9uR5ZxwI1W8kLrVUggAGqRhUn1YUsQ2
Ec/0mAAKIt4KD9aUjqtJKAYPD4Ruancx+Jl+t1sY8TeXeRoFovHxi0JvNB2lsu+7VRCAn1QXEWRj
vCd3RfycHcmW3e1wnoKzAR2/nmbdNNsrKLlcMYVMuM9NWrjYSa+eIUEQf3yv1rfGiN3WUx9/0FL5
DBvsBVG8v2qtBajXXD+1QUJ78ea5dixjs03KxaThZO5kVDk/CVerY3Cen0N1o3OGL/4xq1nzg9rH
Nbn96GOj3UMT/zf5EX0EOkwylHeP55EShIyFb71BJdm92HUyfu+sBHpBJgrZoVsdFZTtTrLxiIg3
niUterQvuNOViuLDduvihDJXtgZzPmsaslYPaFwVYqs11Oo3zLDr6/ik10x01z3aogOqM64+rcb+
eEjLNa1VzJU41uspE8TcAXVNpuqj0yn9ZMAD5Qu6YvT1BMDj79M7PenWaEKNoak7IlaS4BQn51qe
v1PdPPnH9rY9wWPcmNzIiCwC/onfrnmgXNJQol/rGQlJkIxE4Gi+rzu3t6PMYBbAHyaNu6Cpkoct
MAQv11jDA0gCY4Vph1Qz4WolTTtnu+cw5579BrcY/jXDIFT1IFO1ZTy9XU7vUMBbfVMADlpNnewC
uox74xIPhenjF7g4Ok1Vfib3LgdsigOkffl9dhUun1WeI/arhLSgalpIrZm3suNl2MXY4Vqxwsbx
S2txPsFFoAjJoGaWnHI1OT4eFIjZ3Q2j4nGi7nGf9jLJF4PZiL8cT6UxMqik/p1LMoAnzk4HxR61
wMVV6qGQLoILAyuRhpqNlsZRqmbbpeQLG0rrBeyueeuY9Nebw0nF8MqoQl9unVFcudN7A603rqo7
uxJJVb2/V9rjYR1XAnCDGRakQYTHtVQbvAwP8nCMiE2hEKvfpUtb4CHH1CE83pDTJunpNRY/tKCT
lTb/NHMrvGB9c+0xR3DzIYmuFze/8imt03v4WGPlaXXBRGMyZDEqmpqG4sUZ9wYZOO/xilYqsV18
3MMI4eLfzLbkMFCXb4A+vtOnPs8QCBLY4IuN8UAbmxwxvQ2R23y31XHS4+Z2uI8GM6d+uEJQ8onO
LWVAQiVP77IS+p9EubEdw/narkeT26TMfwSxuQaDiQfXMDEBBp02o8uxyAtR9g1w/zBJEoApIEvB
ZmkYVfpdQT0hXVSmhmG8QygzW2GmRMC+juYdme4q7HswJ+d7zvobXdJJjMw4Fqy4Khuipu3p+TIH
fQlc/yqKClSZoxJIFA6o9kFu12sM7bnIHFEjuCQJHuq/bDN17OrT9kqVP4RQLa9iqIvf3BsjS7rr
xbUpk59C4tqL8erig22Buu8ymT7rFH4Y4I5/vf1wYBX9MZ1AG8OyKxHOwHAikpUUlEe39Th1oCr3
W0/M8D885V6Q4JIGp+FXVhEzQEwJpLEzUOUiOq6GTzSPqTehKEn+lb0CdeJA/9T1CCpdK6bG5409
nFQ8kU9BBg8bCBP4kXl73tmdMesJv7tY89DHGeDIMl5x8hYduTVWiazExNre0iTmd5Lq7W2N7hUT
EXSHwmbzhu1xeomCOs+7if6iVvHj0RO2P6dK9yMi2XPDcnPoMTamzPAdH7lEqNTIl2mSAAs/FYvJ
K8LJxvzTatRDVaFZJapsH9JxlJsUnyuTUFYVzTc7O0SubkBXZToEFMrIs/vMX1oXPPTGet5ognMS
G5bC03XBcB1KU/+yd/a7nysDPyCEO6YnFXtNU7hYJOj0PGe4aqJOl8RN/ZZ8HPthSq0M8SjKPUUB
1W8nWEjlqoeJIah5eIZHud51tHAdL3gP9wiE/N7LLZl0bvMnDg3lKJBsZZdPDshyOLa09HbiRSJe
2r8pg3fRa3nR8PkbWLsWInzcLyYNBWvHZnxmYkeML2H8FAgxZG3HQPjwy436fpEXIJw+9szOaaqG
/lfE9lGGcyS6nY7eAgy1Kba+/VyIOXGyVZajjAVI3AIL/6MCsjQxAM0P2I9Gd0RCDNIohof3pm3O
8LQWyVGBzdeegvy6bXSR+/IrwBek678PHQgfstKAcgucDx1OMOkbof28zg4HurWTH2CwlL/rQGIP
2o8a7/BrCO6WK+vmJPSuKfJdMz0s0dyAOQF9OF4kKy7cyJ/0lvvG2JCN4eqWr6HeIpCwS+tinGak
iHaaItP99KY2bZ2ACk2ywsNKcQXWWvw/XRF1JnN98ruM5rbFyqwm9nCBiAUIAnvh2sPMC5rlJvj/
Ubira0Yj86dx5zlzy2UgwVLwPVDX8JsVaLQbinFdUxbyy2Be9OYx8iOMbn5YnQTrKhqcRCZvOa1l
n5SfD/U5TknDlnj6vXfRMlcW06FHoEeBuIWLZBF0ecLhFsTgJ5cxGGoGJv68xKdWhEj8rl8KIp7T
xGUw3qdMcoEmpa+/HwuKr+JUoQlNHLMnX9lfxqSlSQLoqzNjsFAC9bS87X2K+uulzAlQyHhWHykr
aqEY/ulkN4aJh0z1xLP3+EciMff0N8mXAqj75401sj4EJ2SlBEchl/Epr6cGTar/MG059lvCc2pB
k49nSn4zSFYgRWRi2VqZyMp/lPIm7XyV9crCw27qpX6aWBHCer0pH+8g315QXjMsrMVj9MqeByJT
ULTY5k1HaYA5TDNWhKM8V0RgWtsPgQBsjYgoP7Rz4UxQBdBvlIXBiTewQpLoOK2elx5O/z6RpNVN
evMiR/NWkJFF+GilS3sbrReHV9b3cYAuhdPf3ythl4ZggkNJLC/kVYVT95cNQKKKWs8+laLCF7z3
FnTHtPIyo6EZlpZXxuAwhBqDLu64aL2E633tW4PF9/Ap2dfwM6/AmW6TwTN0d9G/zKwf1klTHvqA
QKDjlFjke52dhxnwB64oimBL1K9XxxHbUBf32eawfYaiHrALAokdWJH8qRGZG+gb7NIu+v9OagFe
ebm9fcdbCFcEgWjaIcCKnzbL1mjrDD41ofIAhANmKuyfXxV8I7pmxdYv4nSJPJW/krBaviupLIzP
oU7b3JYeVNQS2Sf45y2UOFkQcoFyDc+qrnQyWXp5v/YLwxnd3SrZ+KbC8KuMneScMLuSwMlVUZMR
/7zzqxyeQhOuBrS+59d1y11h4CZ2NWHS5QsThLF9/yj508+6T4iusxNQb4F2sLpGCSKnc0KUmDGj
NeUZuZwSmu+ssG7TI0V1m2BdVlBCL6vYMqwvCDAR5bgNEi369nSOAa0tCyDeIbRV4rmPGcXxSGXU
3OIxDccFhffZPilNM28wvwhMmYfyGZee04+1qm3oJO5eL/S6dOc/CwAcqCSrX2TajRGxOZqBRrCE
sVYAYRx4RKer3lto8xGeRNvSCYwInaqYRgDoavKyz1U5qZZEkRpVGLmaFOPCsdBUOlNEr7kvjsgf
KexkocS3L5juMRTObgglxh/1Ut2feFVAgGR7ywhjoAGlApqN4WDDz1us/CL4zWFKd5ty+WEpLLhx
Yn/1u/iQxwnzPTYFqpnlMLttZuwTUAWxXCEzyFEg6XKzCXSwqf0yh2mEW2qpr0Ca3dHds4Fi/7+V
RHcRR29Klxo4/A6STtSt7hlLw1hXPSF4/TqBdm/6mNMAkad0h5wvdKC1E+TdYc8ZwWtrNAUzmXvP
hE8OtRZIhmj5wvvYbDV0wYoaEhLpAw+UcmJHdd/nX2Sm1+TSygQwFy6nzNRxio4LcQFVYKUv9uPy
wLQdysTdNWr7vJQMgpAipOHmoVbi6KbfQKpbyK79v47/bLqEzDjutQ+eX7aA9VwJrrYNSwHL1AjG
Y0n8sVboatG/Wq1a94ave2iuzX/77mBfQRxeNT0Ogk1MUrDZt50CXwkvF1vPy7K709jmioJwRKUc
5pWxh4hqJ6jXpxXWcicUloPAeJYo1n1lADBjUW6/QbniKD2YQ3TZPZYEU3lZqcBeayoTCjm0lMXy
8PU6vh3+2pOlKe2EcLGUgU3gEAnIpqfpckwtxT4yN4uQ6SDjVVQoeT3kTAAgAln0W2dBEm3FQcgt
xmG+c+FwAZFypBZmL0X/7XbUTQSVVzickbS96G0Br1Rm2ENAeOdUOFmxFz9VN3qcT2JFxds52K14
epVHpt9Ph+xCxGvcm1fHRhz26PKbVOGx9R0Aw+uKUO4uxyd9p90NmqwCFYcUtx5kKcsVp/tZvUC6
nGCU+ZlYGWVvtqLkQrzzaAfLzO88Z4JI35zCA7YuBP/Q0Ng9xYk/lDrMLUjPxQ8TtgosfoNGaMRP
xtl2pPbC4UmxTRbUNnn3sL1jl/40NCGcWQ1VzJSoCxpADHyEH2vHa7uZyAy4XPn5E8wtC9zlZok2
dJCkwV9HaL7fNU5u9BTk5V/rtpS6OTileFviuShL8sGtSlwNKBmT5TWXehw0DWXi8/hYZ3395ckj
jryHuoBLq3aBac5hgYUpVAWg7tmS0mM8poO0vcwIjWvjFYuVRcSBg7upj8FOwwD5qqRhiSYRtpop
PCQ2UnkvrsSA3hxeMh+cm4hgB+0I21tA9Eg2Ypt/8DitBLEIU0mnv9HAMJOy3mZAoh2UrqaA/vlj
mioK0PxbiBRgtD77t1prb7/TdA62czo3sdjLqT/PVxI5jetXWW1gB8eJbxHpq0/p7Rs+SY5MLWuq
HNHXVkDNCySKU6GP3qs8X2kzAVmtUmVoEl6SFzrYCdISpZBMCx0qT/rxFh5xsZ6Y7pDDzSKcYtDU
HDDfO9u4lcEyJcKsX+dGhiXu3s+ebicU1dhwKK0EfVwjvsJ8TmUVCOvq1ZBVuoW1VlDhMbfj1Ocp
ACwuqJhmr8jrJ2WelgoOnty0uloabXrSjjDWwkXleKZXP2nLFS/b7yQnaCv6JHnkslwFqh6+SHnf
p0ubS3qGT1vUnA59grYtSzgnRX4jiMSbyG7CKTewnNX+CUYMZygXl5p5ASSZRCiJTCs8MIeTfBsH
X2of2py7m5HzDZ1IQy44SungjQsWNs/JYI8R+BTfgby53Xli2ZVjd6a06eODndLGFOzm1jTSW4qg
pxDY2vlJCHJGq7bR4UoaIppoDp8DdHpmZWgR3ffsjCsn1b7PVacqXWtoyq7S0hA8npZeZQxqv7i8
BKqGYOek4L9Y4WePJ0K78Iy4q8+TIWWcqRxTvvVf3aCo3qYdp++Rqt+XyqiOBuGEsLCw2wUnXAub
FkkAMDBiQfB10t8PFKK7DgLiTqh0kV9LKdGc1mwIU49TA6o9W6lN2JHoIq0jAVofTLxCW/nO++71
GNPc2OCkwDuNTv/mOdYTos0KrG89saVB5v8p3VsDwd6Af8Dt23t351F39/fqTTMgxucVAASHLL4w
niG5RRHBQj514/GGsikHFBTHC4dNBy+Pl3UKpHLQI/FO+TEC2hKoDVvP0r0BWVX26UxJ/Zxa5X6i
hWzNvw66vECKaOZKLTwS9TxmKZ2m80RMGJqYCLsbcVZzEYr9h0nBuD4Jx4eMm0M7q5m12I8rugKV
UnqLLECRIH2wTLr+1Ay4bP6IgCIEeTwkpt5w//EPTVVZZbzEFk2j0E9e4FkT9W44mArCRR19VizQ
PKbHfCt4VHA48kLkpHmKqIbhwWHIbM0F/7pZRZ4ouZYLW64ifdYiQmWA6LmAlMjCJ3VlAuB8Wq2G
mNdBm2gXzQ3imiaPBp9YhRHV/ivxQFGjTtH+yW4L2PdvnTK5Ko0jw4OxUTGDi5IfBMOnRMfxlYFb
3kVjAULPllvOV1oDuCCfNmy/pRmE3HUWwzTYdcVkXeE2gpjIt4TL8g12rfDbIgZR8PSPS3eslaQp
FaYT+5TYtcjsZ8zxzLMWPE/+RxMJMj1zdZzzSHIyOtJWcpnG0jEo/2Z85NEZYFp5ccuY+zsS8bpE
gZomYRhXurEQ8a3u4W152OOaasG7VwLBJ8gSXglai+aubY7IK3mBdCzKR7VXpn6rh3FqjlUg9MJ7
lsphmnVBUN/QteouPCjcDqs0D15VK5RKEtlzZxUn+BwIsEDbQ92gYrI4XYvK6hc/6VYcKzNUN8rR
uhnvzssHdW4IaJjdp/onMEQCLpKxVlIXr3GmD0t1JLS1sDw3aY1qOxF35TBbu4T4WdlFi3jvdTP3
iqzeyeW81GWKWIW11TTW2myis6xauSZ0pOgFQ/CzQyQZiRlxk9vVyQCDtUiPvG4CAgkeIWtd0JGP
LtIRTZNB7cjfVGKsKN40cUiq/ZCeKNIRemhPLVBDaMj+r41+V/301hVRyOC/0n3oxmBlrbANZDLZ
rOCzYYl45l1GajDj4W+i8gmk1NpXQ5+hzQcNwGlRYfnH2mGLf1GRq19eRBZEUQKoRwY231K0lmJg
t9o1v7rMRyj6KOpmpSrlHQmI0dMtJdeCmq4LOhPvsKPRCjkkzoQ8kgljCbOOnKXtCDXNLAdbf+eY
oCvOxYq/qWNEdg3b+ILk82HQPkgdEgZbR/0xYnYdc8ULlsSnJhGUPwkwD7WMd62tW3IcPNhBJVgT
Eo9IXd1owXo+5o0zwEusX1wk4RbgbhdfpC/8ea8pGvqHljbr41QH2oEYN7m2bQAHsyuAD7bk7zCF
apSgyTgSeNr4zXFG2XaSE0w2f+KRrPuGQWicz0ljTVJm3aGh+Rib0JziS2NjT+HeEF1kSlx/kDPJ
dXWzfTDTWgQn8x9NGtnAOWy1UEBBrePFdbG74cBOWbIim4swiwGHvNxlWXPz4TriYkr25F2qfVMU
tyjOgRJpd6v0F+TK9j1rEGWvFN2xAuCLL+/NJ1f9Mob2Ks4IUKwNIsP9wdjCiXbGn454nSa8z+eb
9ZiP4vheRkKF9baHWL+aQ5iPSetRnscnIvwnVes4yQVPnPtOq0tggvCzYSLwElHQJkzDWdijdxO4
IZFktzHg/SO1fySEE2oyTQidYZsE61BpxFYoxdcdDaw9N4z9fD66meFk+hUiDWvM+uv68OPgK3nm
aWp0VmeNIBDIuq5yQqclNqAQjXAOFrYi9FcaYvd9Rbgt5oYDKzx2mGEqPN3QoToVcfz2V8JLDeOx
othe63iEbRr8/9jiN5MOF5tX9EpRIi8miV1BrFXF0+9T/8tmw47oCj9bFERC00TJi2hKc0fk7xGr
LYKQAh/N8I7BGC6ifKzXGbtsXWd8CzJkslCiR6ACuYHZI2yzXyOWnczERw1E6Naj53NZkzp+9N7o
4FBQsUyqy685SQb73ssisXuvQ9FsT83aDR6KSyLb9+E8A4oLZ9BKf+QV2OlXPEA71cX9ED+BW+Pi
9Niuxc6X4DTGFZ5/+2hAQCWhPFMH4nX14UR4qZc/ZUC08vXHWowkPEeEYVIjRDPCfXbKbUbk9ALQ
58/j9l0aQrAmSgydrfQ9JbaNJxMeyyrgVxNO+Uim1sZ5ySm63tT39SEfW2GWhgj4iFgVeYrBF8On
8vCqnWyLqNL5kM+ZtC+qPKfjvlOn2iHOAiPAdub75cOVGLzrx9Nr4U/uVBFYfBeu4PwwmkOnR7wd
wwXyo+xpSl+M1npdtj9QBppqGNExntFgyr1g+0ywcHZM92UpVtkrg9PefIxYeODgmFlKqNR+beXv
wY1IHxeiLUXTGU+EMzRGfrhe7SDXJkibprNA6mKvCifDlCItRLuxx6jQU5R/i1BHa8lh4BzCrj7w
NhTV/B2OXIAPDkg1ltJoTM/nJF/pT6vxj9UsKHdRHyJyQiPIjPl3DR4Zy9kzgwjzcoqES60PbHS5
xxXHop6MpHyPwDVIMzacxaEB5KdrDYf/mgc3WeAu1GgVTFLNbW2x/KtjUKj9jr8cLHXsKb7wpdTa
o5pXPDevLU4KytvoAmqvCZfY3olYnPSJqHq6eCE5DOZKpps5xRlKOiwEhkxcRxz6T++RaqmFLR/s
dzSxEO49iTJ6qLi7KDbn3XVZlcWisQc6DPkyGxQdJTI3F9dooTdKqqKN/yYak1I4UJO+yPxk4elV
/PFQ4inwTCPhSepd/Lv2S1j2V0warwdn2F6PE92ZHSCzrtSMePCIfAe0XwIEY2uD6oJr7YBLlaDu
XyAUChfGwo+iyAjipaLJVYfaENwC3v4DcLMqCq2srIOFVHAidUhXWke4JkFFGHLwrwsTPkIVWwXh
mEb2gGX3XCr4TAqxgvY+NZY1+kmFgbX4d02i8O+FCWjMDPWjGu0DHxkcr5/f4oUjwxQ7sOx13Ujt
nLIIq1o7lagPRqxf2Ki2pbWtcEUGheFIbAEai2VDyR0JQcuV+9fCV5jjlQrWR2r8REQIaczaORhu
bQpPaadfdtrjN5ebuSHLYMOY0WVxxnPnK2YcKw8jVIAA6eXDNLSrqWTG75qAt/grRHEwm763SAXI
wNzOqNxjis1A0TdLBriEuwg8NbdtUcdtxxUZoB0UsSvaGuwDqL7Cv0FwjtnimKIb2qiQ6GxuKnCC
0/Nx9sWRAfH6vT8NkQUT7Uh8xOydejOX21C7UuibgD0Zuh//pIUznPD3wrowqnAljL6awftUlbUp
Hho6UtsjPrtZfwql6XG7NKYRhUH9XLUiqdrZo9I5FGKyB6COMNuz5RtZ+zh/VaJVOsrOcPFmyMsb
7Cd8mXRZczH5kBMfZjUDi9M2C+3MGc//Ov/mJxOLP7IMgrXLuYOTrK++c+vBUIHrRvesUoXZtfdJ
9Z+xe+lZYbIj75aKK8RWlS/D+qcyYPzfaABup3R0m1pVhZZ/xUU5QPAfSP8LWgEa8pOGh/Whcfy4
xunSBqXSEsVofKn/vHRoe6SijblhBHTD+T5vC4kpOs2JZ7ef5XUKwO0Oq1bJy1Pm4D/h4VdZeq5N
MAJHIL7SdHddKNo3KJDZ15FHvfQ3ttkHLiJa5pbL4VPxpkvuRWNv3KV8bxAk1Mop4vg4qesq8aKQ
+jjMw0zUiZ2wDMzNB4j6dmEEiWU/qgDtmftdW8bEfXBhzcIkXnVYgUcnEB/QfnZ/mt6uO+qvvY2o
T4K+698CjtM9Ax2hzyPovv4LoMFzdJy2sp9kCasTEitsURkIbWOopD9H+PvWydyZoo2s095H/ZxX
QEQwa1RPLR5D9f5a3V+Ennhk2DE7SmmHNLL0obkX2ztss/+A4S6tFgUjvFvXQjQ0A3zf7GwIv9ku
4CcuivEn1YqOFXZIiLCpPkPPSzQL4JYya1TAH2mNiKstVmvPnsy9fwQDk2FhhLqqIiulruSNZFoU
02R5soyOK0cFlFI2O60D04wnJ2uD4MVzNUR8ZRORbZgCr6Iy/0GESMYiE5o+e5IdvG0k61YkIf9X
nkvo76NhlzV6sSTtkDTvMfdNNzi6rMozBz+d8Ko4L44srw/Azm3wRCBd+IDCIH4yituJ07KalPRu
dYACDoDvAAnW43ptJ5upPN4mPDBGSPheXkKUAKHZfIjTzI1tu6hM8tWSMiI4hlqbl089iCbWMAGH
b+Te7bbLib79rHB1rYvF51Myp2pywYEGnCMpE+qP7vfZoBout6f71e75QlRQX16ww/GdoCfncSTC
EPmfz92kw7yRtpCdti5O592/cl2EP0H36I1iJOZJTpuB8y8xtFuszF3mSh5PKRxOJ46G9YcgxdjM
plNGus0PtiT+YIs+BLR2blqfQ8LFWW8p4VeZLaGSvcCmvlZ3/Zhr5dY4R7gyelCaN4SD6B8M1N1E
mxCmzI8diJJIEPyhTTYjZvevU4D7uY9GjIkQlNIdKQl9n/jjvA79G4xb0abZl6RxHFA0tJxN1Po9
cpKkrco7+bRGiXJTe/048v22dxhVk2FmQdgE0uBaAzFK9rfzjhx7i1V/uskmP1h1rir3+2jFYT36
c3svgauXCuBH3V2t22jKcqrZDmVzOYucHI8j8Ks40EgU1Aeug2yirYUfzgDU8lKruR80nTA74n++
RFHrEXWXmdTIn5z/Py5RgkEWeuwZUoG306YU1lgH7jx3SNGErsfqvl1VjCEI0YfX15+nJm8xXL3m
iqO9dXLfId7cd3D0uQPAa4grGAnCD8gQ8qGlXY9iQZzLZZxlHeV3cfZKqvGILWLLXNr0+NhmFUzC
2xrJkaYG8i5Ky9OsrNjs4apIig+cnPOWy+HElvAbVgLFnyE3MeZoOUOuf8j3mON1sAZvTqly/oZy
00zejlIQMhg4yTAY5GilmncAqqcLiTWPliu8CqVRZn6eztPLz4s5D7hiCMSMIniaxBoMgqUMqjNF
md7q8T2rssQj0gCEbDH3eteiWST8Mm33nSQYcfSeHwst2P3haJnjKa6sKi6PvA03qn3/RfkO978l
2b+6jOf4NpvOMcHQ+06PX05/4THm4+NHe/CdoBoSwRr2Drs/2sNjOjUIiF2AbcVrKhcsV+fgnOln
uAG4UTJ3rsbKkOjmrOVl2Dsb0P3CK33eIiG2d+/MsvtHSfXrGDxMz8GtkCytLeM1r+K4SP1MHwjO
//dFEtHHq/zycYbKA8VtDRKs1zL1x7+WptCZpulItf9PxRzPYuQ8nR5qq7yYahQjaJ/M8/xlJ4mb
cnK8jDnajkY3d0kEx91qNteRC8bxk9HYd/y89iyuvJIOibH4JhX15q4QJjnW+rKz6Wu2/9FCHCuS
qIhlhFMRzruGpRQqUSPQB500I0QjNqMVGM0CiJdG4KuCS3MKz3wyYJFQ7sl+L91wAbUyeoSxxEe7
i+KtgIQUMz264F+zBUpbf/7Htp0iyH74xEhCH9Z4nap0wz4errFOgAXlddyHOxP+dsug1nhq9ofs
adbdmUif6UpVk7vJDRSWZa321QCilznX5dbK+zIvFmEV621DPWOz2Jej6FjEnxUP0XwyQSAFiKKE
KnnlgZgUcwbYEKyqStHbQAkkKy1jLZmnbna2Z/IWAKKgHkB2nxshVfLq+e+QjUhIad9ZsCP5HyAM
KgwSp6Rrb5cDSqyTPAfq5iZCyDRDSoAoVNVRY9ovUxt46XkaM5kbQnSaBgKk12YdAV/SEX9Se/Bc
g9nW9XKbfEaasKdA+qNS4RtpdS4HUfsSTKUY6TWDdtrRfoiyTLmlbF0mF2CUzpEIJ+D7g5LoVBWw
txaDiJrvexW4/AWyUPFVPaxWRsTF3U3G9mqJmWlnsywuOuGatgS1SHNi3LUnXs/fo25NLfuoGvDU
yVi0pQBaZWbHONShq2kK9vqkBEb7tIXaZkFSeLVoHPxLeOgMoEeZEriYhiOYLz1oKmO53FeV7BCI
RE87VJCvDDNO5xx0IrZOBQr+NXBEJn49ta7v737lDew1U5RNTLfHDzI4/YcyR4oo8RsEGDs0AViv
dP5BK1aPmmATdfBPWwVqkkiAZ5YpURxJJw8Lmsd+PA56UxRNeRAJ0okDJX1FBNhGLSD1f9xsI/XO
/yEAZTHqBftz2pDz5cVJIxnbKQt82rWhItmKCa560p5s29mISelKK6X/rEAclLU0Yl2R0DGHVMFh
AKzXJJX/xMBZfIyu7xnAD084q50SVksnT3GWpUXMIIEvB10JGMmU7EyXChnT51xiOlrJnz1uAY3Y
k2NxNi1oJx7RW1lUej9/d8QDnrveEuKPeH2J5HTtKP4FGlvZcYtp+IXaslhUon/dU2maNBPpNtnF
UUtEsO0Ro5BIxvUl9MbtIKOxMPrBtBo01qH9yur2lGtxMUujp7XzUvlHnDCZErY9ZEAfX6txQoZ/
tJ6u6U5s0AywgmbaaTuwUlBa/ain+ahzyMLHJ7wqWiHFVUmlhUlgSyUzljTQ3mdYpeleFvvg9JhW
zoCuUOpuTylbUgXkKmz+bYGSCYvTSFLfiSeZ0SiKjZrODTzjEYVyGIUcADiG17Rj6ub6WCK9r6VI
DgMqnCSijG3SMt/g3zs8Jul/18wer8A/WFyJ2nI5vQ8F5IN3K1QLc93uPYtSdoYjvSL9gRxu71bp
zGv2ByWtB8alCMrUqhgJgsNCPqNpDAnUB+tF2ZzJLiIDiIjKaekZxWrqLKT4oocSP6UBd4BtGpwa
eEgF801zkj/H14KJD6lKO5CvUNvSqVkz4jGQ2+FXV6vIVU6ERcUqLyjiJfaO1TZ96LMlqjsI3Zsd
cOqb+7LPEab73kW87S0AzqnVai3hzbbYKE/kLahb617Y6yEAh8+kjm8Tl0vEssnSCrREqKFHa2Es
flcYSccmf6cLSe8x1olaoGTog751qeh5vlrNpmzT6pw/zPvYEZ8uUvS0AXAEr0pbERCeZ1jczE5z
eRReXu/HSU63onsvTL8otboZVihzg7R/ZNcfsr/x0hbvSK+yGgLZruYQCWUVvHRUhPLYOScav/6Q
/sJip5F1kZwvbLVI7SBFsXsWbYmMBd2TdOpoeuN2uUCJODrmD8dRkS6I4aLAR7AZ27gHvHqG4Kh1
75diQLkFu2senkcP89RUfruhamai2x3FT5B8vTHHX2u/G/72yyUrQiEmoCyY+DX2idAC+tEoUIEy
VF22ILbenNgc27lC9+Bf6TDR8WlX9wyVZkmsrTGSHN+5WyD2IbzfbpIHdk1L8D7RriZtCWDSj8uy
4cgXkCya4D03/Hr2vz4c0D/sIHLXMcY+05mBmGWQQuJ4luB6NSH7JC2kvm3yuCBQuJ7ozTVXTxDu
oibZUQEW4Z2D9nsqHUqlxrio4C/THCE5jdqivf1JT5VCP7Z6Bxbbi8YD8zaE/TA1gGhAZuacE/X9
7EQMUAek3Rr3CV3i0W0Qf6zUPRgINjfHGlvCm8M8JLiTjMK4Mai6Z1oLIlwoSbH1uISR3X9Y/2A2
NveKZw8VAMmVORDpLGGuh5mrzi7eFzavtJ1izMTAF+pBeDGFeasgCtAtkR3taJK95dwjtBubZ9/Z
SuMm+eewY1rJ20HjVIzbeezmO+VgYbR7cJgU8wPuC2+QBZ1P2ZQzQIohCGKWVbpSaKW7MrPmKjR9
07NSThoJR/aEtZZk4vrKNdAbfuW/YvAOHOQwFYJ+xalA0uxz2qbCYrdSKVRe4w5xvdJtBfdXQIR8
DbxF9l7xqrev0xUMLYZDpHDbzd50ohU6R0p15NK5r57nbRSDTbSkiZzecwwHk5F63YN6Ur8/7ZlE
Sz6XoCDwoWHffvhB1DNJVC9b7r/TZ9ggfLc7JFAX3fYP+My6QSaVXt2OFzWwpzSa1DesWJ+bzFck
Bsxl9XnMdhfWgqLCo1zPwiOMeIQFgc9D9qnkwJGcedcBw2nfiKACsChUkSvXJiBkZqKD6XB4kqUO
H9kQGVlal65aaH3nF+R9krIbnEUakm9XYNEWA2g3zZGin+fu5McdDLi8YgcghR0iN4elxraJWpLd
GgMgaNo3OVsAE5Trk6IBC33GauHIOYOzKYoFJIGYZKAfKGWhHW6ItaW12eEwh0p13C0sBnFl77EP
VHanPhjrDeIvxQeYInSwY5bs5nAVfEBeJUslrGZyQzzv0dtfcfGdikIrVbFvuElHm6M4xxbSO8nY
9LbVUpmsmLNGQSs0q5BPJn5uYMl6zuFWEL5cp3kta93A6aE3Os8iC+MeQbemtZWOu7/0V1YjYQsH
oRKCtUuaaimdeUDM1OdDKfayvK88lLq2YTYbURwaDBezxGy60p5OJYlmJwLtl7P9vk35vwYOcrGo
+fIDvMxVEH34mumME8JABdYkWL0LVxx5Cpl5HVMOCUUjp2awsLO+s83Ks3iYPfRiaYErrYMpUAUs
LRa4L1ls/nmPVvBrzWcgJsZ0huwwS00t9Xr8j8vh6vcpV1+ww8QfVdjxxnt+xAvJiw8FGqmL4Mkm
EPIwa/IwGTOqrkjuCW5JNwc0imnDnj0/kwkHziBGuY28Slbgk898CqhcuRYp68HkIm0jzuDvdq2j
oAJZLzgiv/m2vIYyLWWNE0sDbUg2Ki6rgy5UCL24aGdoQ7eYPvH7etPBkPnhTq6XsXpDxG2B6JAv
ljgl28pgn++SBLjmLEOGgieXIO+FchZwDtdsb0wKQaE00kJwMx1V5+Imsp3pW7gKGst2b9vY4N3n
NHx1I9GAi+osK4Dm5d+jkLOLW/vgZF6n/eydzqFcecndlCs/f2exXH/2XLXLMdN/cvtvxFKPZ7gs
dKCtXoLA5tIqGvUcRuy6pNf5oFDahmJs94ao5Ockra5O3z0cC1KaNxmGTq3cPvzEUJZP/XXujMeX
pdxLa5q4q2T68gGz2XAJiDRPwO2/vgmMuYaF/ICKyqGbja8Kkza6bir9660PHrfNUtMLVgoCnIi3
S0LFtZ/+aQ9nQAhcL7iysUCRXAhppvpjoqLbgoJzUaO/bt5P2aC2t3YpmZAiV/nE/e7Oo45IGC1d
bYdYKaO/D311VEINqnUVuqdXrEw7ENatjGkJLObIjYweGlSHamysnRobBb9W/176c4g3b9tSyqdB
IEk9tWeCJKG+YlELEg5q9BVRm+6a0VphjnGyAH3FjnLjvmlf/bXC9YqWOO5lD+Q+CF9M+qJtJuNp
vgh/eoqUVwywGU3iEb8aSKHROsAZLc8p8HNBqKWD1xYFh6NC90WK0vzaBYueyjk04mYlO8U2rvaB
Uc2+nyyH+EnsmLgVLkaR/avp13pfstb041sPWHd7rjsUeQXrARwpAyfBdZW7JMoLihn1dt4vJtKr
ZHPrQk4wXjjXuATjLq3b1SA3uFeI0IZ937zyE+wV4X5InXuM/oPNRJoVe9cpRuQvlQCHq31AH6Du
ZTTT25HNAB12txHd8vRXPCjeWQ58oY3shtD1/9F/E1y4am7ORLdmjeemOBPVlXllWDycwJKB7LUR
X64nd/1hXseQjZoGKQT2B4ml9MYtBxutJOB8E6Ypb41yGfWNo0Mfm93w8i/OhBYR4ns1LJIUDQzi
yStdn+24wUA+syuFmMvMJzgHBcjZSpjc91b/t3bPZYTfefm7WKh7qAgW8QHaSUfUMrz44u1oW5Jy
6/vqNA/qNGsE3C81Ip3LJXW10HbveVp4j6vl7Ah7moYD09OyXfReeCOBKIyt8PIrUZyFdPZMBiH1
Grm0GToG9cdVOSuuzwFy89Imgzzd+6raffh0ju7skDJwLLc3LHqwW8bDNBF7mlVWAapRlwQQzlOC
F+wgWizT4hYqURSl7T7/Qp7Iw4a/iNNQgD232UOFY7y9+Z9acUSDfHsOmWf2Kq5+6AcTSBCW7Drr
HTIhZ3WQQqxjiJ09jMZ42/X4suYpxC0e5LTnGRmQ4Vr1Rv7nnq+GUx43D8f1JPcKWQNaUhTn9VVe
b8aZHDlGNKPn9JHE8vO10WyixEfUqg6jh+I4dT5bQ/6/8iY+j28VrEcJhi5xNLLn0CNSFF0Zlu7l
GYYVFsn22OGF0ckn+xSYlp/fUX0CPYnfq/V1qUMWDUqlC7ElFF7DlR+eoS1tNB6uW3KvegVNUkCd
tFR2txgIhzoJ/ii0LBYEpGF210/a0UITlvNTQrRLbIAvke2BSLaKdOT5yKXMdLb6zFIbYK3JOjbr
jXHa+xLbgL3g5o1OMGMnHI5rhqeJcH/wXtXcoN+c/gNI4fYgQu72ngzgTYPeDwInApfTQ09aQ939
JpxAbJpYcBk1OUqSzhIyPMsyKijKNsyVJVLRkOnd21no8VQ2JwvJYEUPP1VjOqKeoJxSrAF5MJ9g
qSbmkiRQSc5SU7lkI9+ImXgCmi/e1YZeLz8JJA60feHUOqnpoATVKiZuW/Vtp5zHP+vw3A3VvefP
fmOK0e+0GorLviE0lrHVzZnA+czWyuhSJ5p4wONFNgmD+qd/mOQMHxXQO/hvNW+d8EH0nfHg0lnt
SbpVF5FlO7DY76RHmP1jqYZO+dsD5E/qjDfXzEcFOvvjvAhxrcG44jEyXjNJgBKwmmTSO4hkzW9w
OGohheBDKQpwVrlhmdHB1zJGENUnjsajs8Ya9OcCd848Lg8yiDKOMMYOiThI81cRnx2xV4KHB3qD
z/nCYI2j8mzI3oaV5r17TFCUDB72egHn0Y0Eqr5qY16GRbXybKXXYA+GKLRhZiMVfrYMMwGWurVj
cfXV/ALTk7u747xoM5GCA9HtVWObRYEbX8C6uFUG/aMBuZxtZJqzr15grKZROnDDT8qKEsE969dq
Qf9M9BJZ7aZlWaQ3UmSs7AG4nUzzTQyaFucs4EwzjXNqF++akX+rOeLZY2vbes49vHnjFBNM1wj1
0lfXGhfjZv3bVnf8e0n5KqxhikPuEiMpkSdhhiUb1OD884Mj40yWT0cqUOjOjvAJGpsMdtB4H0l7
k3KDypbNdyGrp7YeVFSs59TiQ+uU8zUoeSnh9TJDv8L/iEqDxbqJfV0IaI0728wihOijm8CPqi5b
eRublhhQXYp75ypTFtFd6GlDuRfoTpbN6iCGEFi1fVg6Y/31ieyDCNshWtCx5aFHLpXg2QXQmkCC
HdKkIbzQai4yVKXTy8Y5N5mNjAx2cclLbs363EZRZSopzfxah+OPlGztYmYePVCzLaw3FusZP+Iz
FeVUX9SYCMgWtowfSTxEWRnK37bm3alk3mygCSYW/X9uyPsgUIYDpz3NUs2pWN6m6L0e0UjZFafI
V+Fh/F4XRA3rscQqZKaOnxPNZfig93nchFCMUmV4l/1evB6KNf7jqFPdyS00G8192cZCHxXx0mcX
lBYkFo+eBvF8pZvR10IyDH08O/8F3irfkUjGQBHNHsVD4C0jXv694YD5HVyEXRBhJnBTWCTSytOw
V/1cDsI=
`protect end_protected
