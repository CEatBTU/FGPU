`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eQ6nhT7GLP5MtXb+fBlbtE9CmT+npnamn5AXBYnTqfyjeOq6DAIwn6lQgTicnJ/7b8vS/pIqFxJ5
z65AlaBqqQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ePvgcUCXHdPAno8UEDNV9Pww4PHTFcoymZ491nBzb8ykBBL6o6NnFLuEgwxxviKgq0H7FWPEEF5y
7ZLIJXzda1ao2w72+vmvWH2EZiuCaN2z3rPNz+DrfsXwAzGb1OH4/Iehy3XvXtGI+zucH7hSsj6a
Sc9vBvA8dBIKfwHll8M=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dQdlOZYXt9reqa5XybzLiaJAnC7PUoDuampMZ06ce/L/c63q0Q1KHkbmXMSMS6lB0N1ReSUcbWpj
LRlGAf54lf/vI0hCDUKC9qOMkfB3es/YMzriqQ5y3aqWB2iF40eOUGfvVNgW3SNszF46OzwxnUyy
6s7ae4HTuu6Oqwopmts=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ulzmoAatkfiB21vOKwcHgYwoa7BgjojqhgHDogYEawtrOHEVucioVeg/09JBXSV1+1CMAQE+o+xo
TYQoBFTxNbgb/B+5EnCgrZE1BiPORtAC5hOAj+HPBOOVm2mKA+QWDGunM6eHx7nJAgBSZg9T1kSP
eDygE/deOV+bjrO3rpg4lYTj1uDBc/gqNdTHFpKqxuyoxNx8OcaKnKuxzrW35ZhUKqACkp5kC+kG
KelDgsp53UW2XScy3KdDdEl006PI5yNCmgbk4S5iqeSNRQ7MMmIg6hix2Vt3lFOSl5HmwiP8A5BE
3f1x2AvKprXs7WCGiBI+NJqQkbQovB3T0ml7CA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OGtogh+d5rJyPeZ2theFRbW3DATHEGeseww+Pf16AFQWeesc5Ps2gR6yhoEW66CSwrYkGfxk/+bn
0YrsH/HdQo70gaMKCUlaK5kI+6BRzwRPhe6gK2gUTfsBGgUKmCYt5HOyc6kfC3EA07RqlEl+KnDn
Z+Vweg+pNPisU/C5h2GCwOrJBgyua2qstCNZXCViH/oG68/+0B6OVtP6FsYMQ6Ffyj9IhOPe+Qzi
ntX+aTvvTuNEKh9H7VaMej/Av88br6g8iPHrBXcroKOfuGf4CpdRfQGJ4hrUodXcFZY69Z0DvEuI
tAtNz/BCE9leHmEs8edC31wz/asz8IjBnNwWrw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YN7C0KuBvDQtiCpi8qP6cS4kuAQsZBZ/QATwixLjifIRlVF4p+2Wq+vgTTFt5C76A6zV5MlkSu1P
De/LheUyN0bIlepSnrBXYk5bHJ/wtCKf2eL52S5bBQV4hSrTHSUf/DuCmWsO6nYRhOobBBh+wc+B
hQWuxi63uOR3qpe2uUP0VjroyoJ8au72wQAUSpLYpOGiUdHScchVkm4TZ481JZSNyPMnPorDUQZL
jGs3VLfQblegSlnSPlyLBb+vrttOFNzLspmj1i1Jv+DKfUhvr3MLnUyGGg4iqNgBY0huFW8bIOHG
f/mM6bayCz0lG2m/RFEyhjemIQSpglaRAHB99w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 67920)
`protect data_block
hatu1u1ZcAW+FJ1F1qIzVd8M+jrmpd23JO0sQ8zKAqrAfC0aTwA8JxGlgNuDtl4dBtHwl4mPL3Ei
ukxGIC35Vheg5Tv8KRq3KVpRUJ0D+I07Zfu5iZSP73RgPlR5umqeXbcapJ10PYPrVHlAE4Gnshyz
+CebUS4gcBdkkpfJYIfEckmylDrwGt+FQeJdkNsFAWBLQszh9Inb6+tpsiHQrlG17OrmPQZnzvVy
UuSiuxJTj5TEorqFfTxjR63TpGOqBkqOX8Yo2cp0WVFWnDbTd/tuhUbgGinebdLp2RbY3cQfWtfo
pbfom9sGNKFME7KjcYn8afh99AGrEcQm9Wox/VDBiSl6W+C96ur0fJB6AedAyIclLQzOshQP9/PW
va7N3n7eY6P+TIyUTpZWWvofhx5hURk3b7PAlBtYfmApp5v2pu/qSrDenvFNOOmaEvmIkNgqHw2U
g+va71Eqc0spz5PAS9cTC5ipVbf0fCLhRyIwhr9QpmRJkqDzwD6W9+Nr6Rm+FNlhMZm/hmpUoFhV
w19PVNGraBy28H0eqHcuf8NGhAje/CrfD5XQAyCkD1mlbmwddwhHCDkXwmsj65p7yT2gNLy7bAGV
CMga9uCAoP7M+YP/kSaAFYEZN0REjug7BCN09kn71DzL+idq+l7oNkBa1Tp0ZeCVDOpdqGj2kNNw
XzM0Q+tu4U63XuK5fPLGEFyJy/BHYSsl4j/ox6UzimytSMkvF10/nacuK83L2DGZTj6ZOessuNQY
GNw3F+kBSZCJcIUcKm462c+XifZXUm9LTHO3iDBTodK2pz4a0pT5KNBHTw72mbc7+MfPkZPtz+Aw
km3UzPP6cX/I+s8RIGQiJhZy2wXyU+FOsYt+4cu4G8sMOAMlNyX1OUJrjRN1V3Ip7olYSZ2ZWZNJ
582gpngwHypkR1Q3q/RAmpH4mvSSp9gT7dE5Pe2fSZw2Bjo5UhhpzTFVNqFHyCsOH4EIwau9d1fa
3yj3F5Dyk36moL2VpEqBC81ZYAOICrjqlVmAjVkD9Rg4IRDK+BgfZpJgUFP+i+TdADgoTt4ngU5W
89Rsi6onDiRhWUQSMCbdc8dzvYd/U1Beqk6YcA5oUvd2KgjTj8ruQq+uOwA5rohHYRqpfEojxEpF
eiIkrgao20ZwsmxBGuKb11K1Ps76GlsFmljHMx5Lfgljd21/lAKFa4/4XXqAeIwXRlLlGoSTtXgQ
fU+c56ltPrOgQURlVR4eVVtYaYdocq69zy2rpK5NTvs1Wh/Du5y6BO6FcUTFJyGqqxr1ljyGhlAM
pzZi691jEY8Ck0ogk5GRRvrUOipqBWwzqbzm9p1t+e5Qua+LVouFUc+SSV372zw4Jk7XVPCxUA+H
B3ZWK2LfalyvlHDtOBheXAL9mysRu5jB0H9MM2CPPzlX4OXZyjhMdxRzcphHUZV0QIhxdZ1pN+hX
oB36w9/9ib0cmslRx6Ot60t3ivfqTKzmrsY32d2/EXTthgbVhBX2/rXNTuLLAQGJMuGrQLgVul1v
EwrIwJBE8HE9/S8TBmddP0lHLrzWk7Lj8nZFb0VURWoqwz+oHFwH9i4J2yJap/2MpH+Wpq0duTDS
/UYqt1BfSI7yxciu0S9tsi6BmvYpQ92Nm1OOZ086cEbV9vPOJzg7Pd+oB1UppyVY7zdxGXNpc6+b
M++F6Qc/iFM4brEKeJUVMM75Im9XzmiH8UMoB1k8p8Q3pu1YO6YV5JtOFHREVHnXEsuWxkwUfz6D
kd7R0w2z57kUmhBCl8UQ2Gl8jyPKwJN13p682wf6o3Ah900UBPThNMySiu091hNByVz0lrFoIoxd
wNYu6veB5qX7IFAF+HQJiFkvC7RfI3rjYh/TwurNBfXQDGEy/GQvdVCi5BC/KyAG4fVuEnmpp80i
SBBKz8w8Vu1zyiYRN3rf7LCvalLZDR33HUgjoHiztEKEeNGy1tdgXSJEGFKT+U9fgu6vf7vDOp2K
D5dbqaDzWmXsmPW/5Isyl7G73gtu5zyxqhWVUUmzxCilvpIEm6WnHRR04KldrvRVWf+2xUH5NAyO
KROR7YGAVRIwU8FNfTM9WQWIo9QQiAWcfdC2WAcJ287ycgYj07RyYfzhohZ/Bvl5pFTKpB5bwFTF
6HcSPuVDL7ade4G0jD4dUSQCc20kVBPq7eoiJl6zKXHrYsPosz7L7MHSWhvHfmGr0WNPxiBvfNTP
VZXikghW6lrAx7+Z3iCtEq6RTk/Rh2l7zuR4TQsjoV9yl7DTB10Qtl5nx9/vJXF2CIcoV0RdTZtO
9eoCvxV8d0soMR6I1oe2kYr6UyLbtyQYgrZsAqtjTGOkbFfLqWxQnI9ooHyidT5G6vM2KTN6FwJn
vXesayVB6hGMdB9lladRLqcIIXoJFNHbxLzlO+ZB3hbc7wtoEw45wrN5tXMktBD5Jtn6OrWWbqT2
WZvwtxzWikruLG0a6m0XSQVya6DHNT0oRzcD6MxzkmVgKg8YQEfwVjH4v23AWWBd4mcl3GsMADlq
iDK7tdS3TIpacVsWhjZOXw4xmBqWbGV/ystel528hquS8Ny9ZG/vBDi3AQuqbF1RaqwTE7Aplewd
9vNIGsrvsgX/NQ4UIsEgoWFd+sF1gIQag8dke7h/fQt9wWLhZD9m3UnTdsqWWD2hurg8C9wCxYb+
9HnyLdRNEbbC8OnJp/dIrGTd0Z99kEspEFfBTDf77praWc1UIsMCvUjn1rlOWNfV8Kv5krAYK6sA
oEuFlIznWUcn98u71kvUAdQ3Gwx7pdmHy2IsbjhuxhJi9thqbeIbTZMlB47onhPYWN0PONc8aAcf
NEUTaUL1JVYFQsUQw+aS2NeitXBVAoUiue61nMeeda2nAa88OFNDzYnCCKsgnwyG5eNGxgYS0UtF
XVgsNqAT7tnNYiCUq2c0fauJPDT/5by2r4Sa0LcJhivXcBekEe0BMGME3uzG5Iqd6LT6Hf+A6ijf
Gt9abIA8UzA8y66AV84zbmeRWupsSUhqVvhcD4uiIHvO9f3Z2RRJag7d5GQRzvC/1n2rn12XGvyG
90NGI+FjAS2s5BH7qR3n0g6S+9mowMsWWQ9HaG7ULBgzuBo73m8B8IsT/3Dg+sM3WQS7NI88cbTk
gGFEB6E4/OWSbz2azeTdJ1NVcNXdrArqSoezPAjco9W9+psc5AR3nEI/MESAbejCIkpeApRc7oQP
do2pbUM46436OYAvJH8tA5K0ZdTyyE75tgusL8kkgju9wd9IhhNCfPxYnWd3JjsBmXfa8W1AzeNt
T5yUJbsLcLJn9W7oM6NKlgZW9poqodkdzdbjeB5Qwh8RFowX6oke4Cjs6S4hzG3Z2A2JyBqhoXYV
0wOa6DdGl12P8UGNrYAy6gnKkSMgbQ9WFbm4Ju0v+mjLDO0DCCWBZKgf3ENHk5oGwcunf01DrsZK
dsKyqITLuGxwNum64KSk45ptl4XErbNRcMMLKNk6F1iSd44FqgHcaq3+V7nHawyGGl/UicwXGqf9
TYUHaSyBARN6oZuUkeZsOr6BBqCpWUwMWBLJZkNON35iykZdR1Xb4sf2IZ4PgXvlndCiMeGcVsfN
3YBlHxac9930Gk/Lw+svfMzta8JO138q8ROBmnmYRsOyIPhQ6o9gt5cO3bOs2PCp5FEd2hG1Iwg2
C2wWAGknXbIv4LNbybLRzRNpDMx8sxjFO6DN3xagbCnmMkQt4NLyiRlZWdt0/0joNx/inEIIATQv
hNMUytRM2SQ/B1/Z+5buu87rjaCOxk7VgZRgrsui6UpMr6Qc68T8FwzDhXwR6V/wVfrNyAeQ9g6M
ogB6JZrAo7WWwc3LkAGOxVKOsi5LrmYpQ/VFzQ93tEcCAyxLXinkSpaBzTc1vTnA4fBljLUnvrbg
kf8JdUSFzHOxWMeGci94C6e+R9GHb8zk9CIFw81TEiVTA+aY+9DvbLATYNHbTCZSfubSnBABxNBO
dArHPCDw1w4UycA6N9rHsr/fxw2HC2s3rsfm0dV4eYHyEChW3JdJ5RTDvPWykPxpcIz0yZHdQQuj
48ThWjT7mitpX7NHjsgJ7+sQCmMJ7suWJpzr37SIKWQO+KLKQiRHcCfcSzepZpfqfH+ZFUf5yK4Z
zBJATxksdWMakwkJMoDasC0WlrtM3/P6p44FQGbpngbBOtaFYEKBcMw2EVIFWSnzN1L2nzySL6HD
fBjNFLuVEKkh3IgoCVVa5aWSAHPx7dexgRnra6pzQh9Mw9XVoFJB7lUUdER1w/a5KDLsQEw6gWxS
MQG6c6/T3xB7d58sfbeR7Nxqg17SpbLnJiuaRAwSnWHcJavpr8CEtBD3ONQbJd2I4gzfTcVr63QM
w+Nkxmi5dJGqulzS+v2Jbnf7KFO3XbEzX3PX6B6EurnXiz/L2PBPG4s0tXMFfez3KJDydBJ3nVGx
Rwjt2sYHIDnoye1bNYhdfrT2tgS1COiraWN6l8Bw1YKG4isNq7KQG52vx+KfmreL/DEidrkO41Li
d8osaFTPjT2o9OyXLQf5n2V3/+yPDfFMpxjEEcenUCMeMC1kZaAXPddaJInbfUdKJ3cgFPsMNL/I
uqy6RLAEZCit63iZbIGn14kKnzwpeUrS0fL5F3OvpCmqvveCdzJscx0x/eqyEk3gWPEbHBUHqelp
7ZUGoQU4dkUIbfsXvN1OVtiLWJPDSf3w3oXwmo6dYOeDemVo4v4b/kNwbI3/MrbKzDE5jMLHQ5Mc
6lBdixtTwUuyppwb9U7w2Rp5qxPRGTtqXs9FQzwDRmBxCbIsmueHYysjuCtwMERioWpH7QxHdc0B
5p6TaSRlRCDF9jbeSftZPTTmWOaB82orBXz9JnIdXwnP4Sg511vXeT0vRz+cn1p2qoP9U1eyxec3
o9LQgWtVGN7oabOZltNNVeSlmdyo00I+ICc65VQeUYJZkMoKwBJEksl1ZfEan9IBaeLjC9zVz2vP
Z08V+/vG8jusojakwnCWJFznrmYQGjSiqlRAwPxhA22rf419sbn8BJATXjZNG8LpD8KzAVm8wEjg
XWW3k6HVPDVc9p7aVaBFDtjag91uPxB7rHcWBrb8aw99sGmAM/bA3sHK943cWTejGEY5Sd50toUc
dyjGus90zUeiyzDTeTHYcIzuTiOKByvoVC4KnWadWdcD5m88UI7H6dfCHWmds9WVLe0Usr1lDCJ1
ySiZviePoN6i4ftctju+FnuBXUd3fgUt3ve0C6iPaj0FodbiCeFmjvF3d3R8W2UYElONuy+7bpS+
cRfnWaF5Efw9q6+Py8PRN5NDwpdHYuJY7/9oHY8/We4tVTiitQ9r8N0gkDmDq+qK3v2fAMFVhL0o
UpN+Fkyw0qg65ph8cohQvsUeHInzFq1UFv5LLVd8OHZ5UR5JGxFd1nQS3S1K6UWtSDdJjBnKzfeB
oO+2cjjvY+FLZ2rLC8q9gCwKnJ6Qh6qRubhZDFJujqOcBrAxWhQuBtVle1+7I15n0pX5V1dDBSCS
7OPZxOBINNeqC5yHNw502K327L6ZyIL1YbE9u9Qn+nbutBfMenzC5/dzz+hF1esBzsvHwnCPKCbx
+pboxmfjuuG3tuBcFWtCVofAH4OrNpfURN2pi2V3VCVZYmN5oq8jiIE7KK1fKObHnVzbZpiCUSGf
T2HCDExtUNOqAmA2584Nr7d8o3P3XwfhECLP0p0BSpDdGlXxMOpOXqWkceEgpyntJtebJWX4icEi
ne0KMGgMQj1Ouc4AfJ4uAXRWj75iulpGZW0++cYozzI7VOxs4w8oPYHVfvk7zdB6+DAnkRGYKxi1
o72sgnUsnmm3wekKep7xZZQ5EYukIJ4v9OraSVBjBt8N/4DcDaVCN0QKSRc2wvnkOzFXATXY5P0A
y2b7yhDU2Oa9Fy2rNEdMlW0e4tNGLdY0jOZj5ot9ZgxzWxQ0Fty/SMAsb9reBHY6pjPGUdRVUbE7
c8/jqNcAwaxQTzIPcFfdRaRVFVUJqvUMJOJ00HNW58A7xH//OS7JqAv6vc7hAJkzEwnU7k/sreUf
UP9R5UzXwGxWtjDQEYsW7M6fOom2Y0RjbOim8+z7j79sSeH5G4j1k4H300FjPQnZ+n4ReRCyzGpG
9IXFt5CST1BPSElRhQxTIpmHFyPNbWjxTdGZNeq5u7MeRNNF6b4pMnLTqwZ2KINiDry7VLZi7QWU
eaOCKF/WheX//W/QKNsp1u71e13tR6FbOmY5jLrgqT2QgUu6k7dRJdv5hgwWGkpE/8pjk/m5T7Zs
MFf4I/Yvt1btPk6K+XbSIZHXE4zZmT7qNgm7EWzAqB3C7WFgIZbXWR+yoF1Nd0s+x1DckcMcCD/0
PQIdw9dpyoxrtddn73YneQkcxlDoUQKi7Z0EiLmtV3NLyECGTf0AubBr0H2Uicb7UAGvNML/Rn2t
AQpS0aHs3rpQkxVOUXKwARnJQpI8t7Rszj7IjdOaNUuHSgxEhDXl7eRGTpMKNrD1zmTMJDcaOZ7T
jDsgfpts5wmm96hCOY/8Gr/JMg3jE0ELzov8O9RHnvR/bds8NVI6k8/XUPN3uTyemAybD2+Tx4M6
XsUMWBJpTQM2dD2u8hbSbCnoS0GR1mlari3W/D1ue9gRoFrl+dZgK3Lzau5DERRaFZI3VeqZVjkA
KCWppDWSmEiw9FSf55es2CrL5uJ0olKRBIc2m3WIKK8U+8hcgIU1RMJEDWH6vLCcIED7NtcUsM4s
Sc4axZXBEOpiQC5+5L5aCyy6Di0ZN8xmfbVM2PjvmSDGocmkdrhyjZYaytwyH0Cutn/JovJA8OrJ
jJqVFdILOqq1bctrFfI3YLH1PRZVvuNOx/HPBrn8/SRIk2MJdQnENquF2APwvIgJ8H5dYTKvSYOM
A+CFkMcFUkhSPYjjhsEs2VMQKk3Osb+i4f3wbso5LnnyWyDPiVMpahVg2mSQWuCW0W/mgdT7GiIz
3z3jX7qboZiJxIaV+OqfjNbGk5S5G0X4qKqqyauX8dhzLVFw/oWwqxtJXVI//KFqQzeZa25UyAfL
mdn7wbWXgSeniJ8wY/WPczLquy25bVkQzy8DCiuFSoG8YSJGnvQ1MOGwSNkF5kfXCOdLNGjA/LQj
sReoMelZzzbIL2FYaZyywb4xRIL4eww6+N1+QbKukx7I5iD1W1HxPfvJhTAVzSNIDHlBOi8GEVWy
Ke8vjfj8DrgvOouYfj3oNPuPjF3Sw6w598xPeD+Gjx4U+muFHIYVoZdB+bFK8KKXaVRhdqtMq+7O
TrYYp2KQIaZBCkehLRIWe0VrZk4E/hvG1joc6/4WikUqPLcG65YDNoDqU79IBIBlA6hm5oSU1nQI
o/0bnC1/AXsgJLuTdvEhgtvYPQq20M3DZz5Fsp7n+9TV1G75z8EkFtF6ekPjIfR18M5x9SkpKj7q
hxrISgdlaxj517ncJT51BhMNlZBeKtGgFIV4T+56EcaRlDCk/5XKDgKegHRGDD2gY1E4uTCtzW+Y
rarTQ0oSW8R03Qg+5QMttDB5WGFdDZSAwAgNJ+MbnwLx6Id0h4WJczmn/kEain3bWjjvHLOBEtDi
3tSEFMJrGtFngYwO7hhsfs3UecwAtsSEk3H170mUd3oQ2vLl0a0CI26rXbPmgrzBhVCnfuNiudyR
glbn82eemq5U3BqcdUGHKGyML79w8rFOm6U6L0hoBxL1nq4Smx4biZ4owpP/EL2ybVxMetIYDO9j
nd1PHmjY29lrCEtDweQC7wxRd8qMU8KE3ePt5T5nNkEnlW/RBIIl6ae+Qq952Fvm2s1p5dmigVro
5Ma1WHisnZjwP2OuK4zzsWwvTNnbUUyAF0IY/6zJUIrl70vHh1upjLH0098pgh+6h0vJo1It7Usd
aziE3cLYkQ5Rg+22PkqnJ+qyZzywmvzN+LvdaxenQIQsfgkfaqQzym0qYhR98q+rNzSG0k7iU/bT
MCppUB/X6OlND/65I+RSxgLHjF8gt7gcNXNi8od4dVwYhxte0Jdtjvd49rvOP8w7iXfclIMFsmKZ
mf/cCqwK9+P8bZidvOeuJC8fiDqc+wgAy7gOhC+63r8+tb8HLVXBnNn4NL+8ub7XTuhkFOBdbfUD
z4tFxBWkqaFBjC6agRtbkgnSRAhx2l2OukgWMO67aG3oMPH2MGEKuZsXk4FF0v1Gxu1FvlGneYrS
sY1qiRWX5BuLglkjZtyxJv49vLa8TvishzZV9ygWqmoJ+jw78lIrTXORIDI1xwy6hUlar6aKJIiU
FlHvjlBh8myPV+pkG/b6CSlNSNErZr29KabXQUiOaYkAJTXqT8ot5XRoyAAjlgJaXl1MM44zXsiE
ii7TfXweDBcBdDUtboMqJClN8eO7zfsYN/OcN7Awc8lqhLZjL1sDYeviqpflwfHAK47WVVySGz1u
ahRgVqkXzYja3uU9N+FDhtyJB6CCylX0FYw1eBEW90gfHEnxZYTNYq0osQVtGNMt1DSrauhEibE3
XLMwucKHDOLLAr2kNDTU1L9h+U/BNe+588xD5re+azXDEFLrtahp69n50gxTfIcxy5Dq1i5eTVAk
K6+PZfbC1qjwpVLnazPdAhkKzNtvnMnsUGTPg4S/ehVnoqDNfvrYjFLy44uMkbbeEMKHxyfPpsfc
TuUlu4C3160m5CPUuSE4QSwhsia4Yw4Dzdvruaz45YW0i42RPYF8PHS7RU+y7WU9klyhQKl6CkVU
NDqgu+EzsgxKDtFUaRmapjePNVtyd7HdJDdUfbx0N6BBJ9NgmM7XSOUlX9WVNRzKnksnnhogYHzn
P3wkyWuqlbnSVovKHrx4/ECC2EhuBwAh4GzojwzvOsVtm4x6Ua2J6/DiQsVO/GZ36pl8vGIzB1eh
AmnMOrQo3RMLzJVMDn6uZCWONZEweasDi1CCvSN5F1sAFsvimnSHDrcVE54u5o931B6CvB7wcgXU
r1+hVkMfm2wC86eV6AopplPL988uS1TUZtXmbHpZnzF+s422VszwYag5FkjkeUzCz9KraVPRlk2c
9WqmVRcELTEpEzIACtlH8cNPvlNyq6Idbq3Z2E4FZCNHI+Sxf8h5i/yP6cHHs+fcC6NIAg+0enGu
W02N9u1zOqXIy4bWQOTeSOtaIFN5AenMKEQz34FD+8cTTVvNvtvLyXGVKXZl614mxPh6OcExBmST
51b6x4QQwnc+rpwPc/+CCEn07AH1urp+Bdn5kFzKw4uOqUkc1ZmjwKw1HK/ln8abL0coddLovcDc
F/reGzGYazDVS0QNBx8PE6uDRhSvndmTcsJKMk4L7akeQppNpVPpayPeEb3nVTz0GyaPPIW0gXYg
w4AKNfhcD5uy7oPJu/VSYENrfyud58dFD1UhK14DHReNZDohrFS89hU6DWm722gFNewy8iwYjuY0
fQZJYV18Qta2baXL6WBOlAIck1elIOl/lQQ2ek9pMCQ9iTJ4MmMW4Ff9EOLa2APo1OvkrkI1oGAW
od947drlNdHGG/3MF4xcNcvoHNWpg/1I+FWvi98SoKNXTP8IkyygCrEKFdwNKcxkMqMOPHl6zkxv
ayPUNQnA+szsc7G1oNsd2htFJZNHrvO4R7FKcc2j8YsfxUuUV2K6k8mVQaoPxBR81UnCaghRsEe8
smnKUM1oBlIdy/ZYVznvO+g7kyDqkNEFLw2b1+KkI8dxNrkk4Y3XjZhHFTZr+6w595/irVKvvq0N
N3OIvuALhYKT+ALqXbOYchT0Xmq7znRGN/IMAJNgaHRfYmoFJ5RoV4x6ZjwzQ6gXmzRT+2IFoK0G
nlPmR90HaU11ToDdceLTkyPS1arbRE3VwfYnecQ4HldwySQLJJKWGdvG/Bpv4G2oycG+M4gVpDo8
RYP2YJxJNFzOtpr7W4A1524QZ2aLOBsVGg12An8A1SPhEZX/OqkxC5FwfBnxhKkAhCLzths4r8ri
k9ivlO6Iq8dfM/xGDaRxXlQeYRskzaNRmXl0rsbGuXtoOneJKr19oq12XIv469/q5nn/nP4TeLvM
paM2uBvNlnPLn1Ft78xq6izjbHj6yrOveSDGNX7zvbxYE/DiW/4mwAYmnodeFwirTHWdLTT++LYs
0F+bcASYi7J8aR1Quzsc75TP5YKC1x6VmU2S/l22/hjeSFrzbN3X8NBg+Da4de5auA4tkZYANbDo
2J3YUpif6KFftjRzv2jFBtJA3T9zub9jkQThIUoVcm7z+OVyQp20molcV80VXhv8NnmMt2NGR8K0
i5uRFTqmAdgYGFdhzv2dnuXRGD6zx3+sluQ8jXIMNyURdb+hBWrqBDsLyy/5mXQuTbW1Dl6UH6Sm
YZHrZvNiQ45fk43spbZToTBBJ0Y8iZtVaAgFozkxcQ0vNv1h0fD2+xi8c7KZUikbrzZlceRN6ITY
ry4u9c5zxo6pVx+0NXxNGVb7vKC4+MpIxCPynhcUKx2Zc8cfWC/T8/HyMpPa7L75Jipph7l2fSLp
3OuqDGe8mypF+DLDGnfeOi+ijvg0vp8eUWIS3gVeWQgwUIkCT3SpD9A75eGRhbmXiLRmCSeHJE67
SJ1cN2q3ve17nBPOmxHrGS2A/DaXH2rsQdtq4uaQtsrMsOLETpCfyhQ1l5JX9QmZS7vYNEbCWL2P
PmkrR7+J9Cj9Uk7T3Az3rH1HvTn/HToFABDaUsQ5F3uAeQHVHoRc6HxI2Aat8yoA2ruSlQwt245M
G62ru9jAdGBmcYUDNSnimsOgRE36TEiyI/OP8T5UHIU2C9h6hizpa8LuZ+yg+RCZ5VBhSwdWM2cV
d+C3YTeLBP3oUIm0InxYBxF2t2hKtjIvWawNducYQ53JWK+CkEFaS9b15uci7jUij8pgmeUy12Ft
g7WyDq8YeMxhVF6fWSK+53kkY8h3GXGKBFb8zHx3rVgbdZZCONKN44gDUGqrPVLKfT0aaR+HGNU9
ESUMHAGgtgU0E4Siow3N4lOa69B7npu/7ogFens3o+uSzfMNFDYWq8vd69+LTzwOZPGURfT/KIIY
Gt7UPek+ovfsKmNR2IbVzZO5WiFDcnmA5wWzRRya/OBe97jk6uwdmuwUCjjtbhVsayrzkl4PYC7A
L2zGesmKTRX7KqHQZMC98ivw13rqJJGydQqw/785T2Es/d5qTHUwr/Vbdml2wb3dLWNkLPJDAGTi
vtb4Ys7MQinTRSmcdhEOpOw4GYRa+fO20DmmPj2pv5psxMCtmXO61K80EuR+kVIPr9KD3OFB/hi8
dPlniXaDKWBPy8Cs4khmreMOZY50LndcQxzQnvUMe2PMcOJQ6LhKa6H1OsSKDzqIFSVJV4Sds0ir
emogBKgC8lDnrSuoCsrS/qdtSswlHvMlNgt42jn0T/7Jz84opVqk9jp6bNRh+UTZ30GLKYEpCXMh
YZjqKC+cOFETH0HvIP5vjS7DEdfE2F0dYVir9ZeJ2SeffB8Vcw7SQ0NWc/gQ40y5mfSW0sLFirfN
fbhAlBDVTtP7fxKwt8DfVU9B8DZA1RKZePZQLbEXcjG2bwJtwsVtGF7//9YG6lqN5pM6lGrym8ge
qxxQsdlRCH6TK/ct/g7cKWCB7noMOQewBIjKmfxOCEncZWapCyEXvRPEHE4en/zuM3L/MieIPW6C
005ADVbCteWe+CqEIj8zmoZsTxZpmmR/E/TdH16UnhlaJusa2BZORlKfCw48DchLNQV+RsMDeU/u
gzP6UhQfe7moPdczvGbOZsJzx+Z36p2DbmCZE3cmBJuu8iEq4sQEV8YOhOOFJDTDeFvJJw0mQhkx
zSQRooBErKa+HqAfo4+wnw0aleUKtbrc/BCqD+A0aqAxsVdoTsNvzhY9cnlskZ7KE+GI3dNREVp5
M3Fak68iZ88OffL2u/D2IouSUToqudIzv7H1HBzIik42HQcgI6szE5DO/EuCBxlGlwCJBv/CesNw
EgtPtglYx3S2VqqBT2td292ysqxi+wQ1e8yJZhNLi9aPjOtGESlkhJX9Xv4CqHnQFGREcOzM1Az/
28F+xGAmRKvXb3ajcnfNKbvAyGkYL9yxnGhJ69f712zXyvQB4Uk3Fc3r6G4LNhAvg7XIEEzcSc2T
JyDCu14Dosj1/dTj1raTDRqexi3aurIl2cvFw4sDkNAbLHe4tJXDwb/Ie2Mboj7Y4Vdiv1nWhwO3
TAzFxcInSF5PvulfmI7Wu23JaeEV5B3sl0nNokbe1bPZLoGm3WkgR8weNyL+J9JBtr23sXbQLsvl
K0xlIQmbVhy9onx1f0uNVSFKmUxTpTFYa9KKmy8kwHxOWb6za9eGm73ghmZfoJRtIdQXf5QUqcJ0
9q4/4ATa+PPQOHetzO9zHVw5xE+7QcXIEOCrNLgCfQ9Icsymta7vyEnlfVHuANiT+s8XG2Bs4CDI
aj/S+72rMRQTZNiQauGJAEfCrCvupE2mPdG198F7Gfp/jw+JRjjjboTpIxQzWTcsLJXkmrp1DidN
hZObCXTcg86cePZu/rvZ7icGCn9R7ToxizTyRkxCxI9naUU4RPixfnNKWQEqwGenJlIk5d8/AeZy
L2OO6ry2aGKmpIEtetkYjI5gI/VFTSODrbyQ5zuJO1Hooi07GwsxciYp2HG31vjfbvxWlVy7vw7q
FknblNM2BYREPXDI7ZQPrNeyS6FF7rXz4W1S7QR2RkFURVhK0dSKpH7Eo8I1ePEjXyfE4msaL1wn
oy7Vw8d303+JvtOQL6pXnrThZ9GHGBRwC7Eu3FLQKvU0a3JerJ6BxlUKeKOSLnZJC+yuCE0ygd1S
MG7x0BNiiln313URLUzREmC5VTFfkV2DzejCg9xHoZfE92E95SnvAb9t8ujn1KgRWOwZDKexZRAv
rXqR0/9fiXTcvRhCk9Rz2BleIWU23DEpKQrAc3HGt+eoPbihDgc+PwGqvzDdSOAE9BpDNEs/UQC+
0qNQXBMmjSgP+4YTn+7sBkPOTKfgWX3CUFJDGyES7vT+pBl6q+NmtVOPGk2nBcGNMEpKZqfvGfT9
N4LZt+10vZj/TV3d6RSibTQKEXfpKwACMcen1Dmm84pHNJ7Deq0st3TgRRMBGaWb9WWaW+8tLmLZ
W/fRANUYRHjGnJgMkWYYOBHrt9qbYe7Hx/h4Mq/9r4Kp7n9kBcnDgaVXByLgUxzOt8EhqcYi1TCr
7B82S1b1qECELuSwv2SLds9/I8f2gwrBlben8Nx2DSffzgs40bABAwtF6q6LZg/nnpXMTSoXSHSZ
SK4ftMzTyGtnQeewvUdyxV3PZrhbBU2grMsY1JtIZ1q9TYB9P3gm3NGTcMEm6WWxHNMdMtPDPnUT
+OF9+3s2EHi6Hiy1gGcpB9Hk2O235751acG272iLtDNmBYRYmZ5aAfWo4B3YZtW4Mopd8iBYStgm
T3VOLaYy+LJ59gRSCW9JfApZPwVF6xK7BNRphS6DY2/PrSgav2PntCFi7Mvx0ClGE4uwkfJNMAD+
Pe5RjqYQQpr1ThgggVByn3YhiEup1GRWySxNULA/+yiUHDYr9STqQQoSavnqBZ1iZhaJjfCYli9y
ow4o07v86rPOO4vXOv/ohkaI4+SE9rq0vgkSTRiQ+EWIA6BcXzA/QfvtzFgLSIv5kc2Ic7emRLBF
OumCpuGZFYV61VPdAPSMoZ44cwh/qNB1zmObPAWBlwVxa966Jh0BNTPOQN2UGQEUBGU7j7f0o/2t
+ASM9yhK3QeahVWSpKqEW88A1baPvKgTWqHvwedkM6p7TgOTY9A2ql2Hg+uGKFdlkzsQSG4wUiRJ
TtVDXVGa9xTfR7lsVWGlaRbQVZyGHuYxngU77RHp1ummSH5/oigOiDJS2sDS1hDNF0Aa9z10jLX0
j85YNnRmNNe3TKfJC1rTCnwaLs6jj7VQwRhNdykIQrcCCcnAAYxrrdevs/eKKoEFJ+WLZ6uUZpak
BZQ5r7iGlk0QpsyeM3YJLjrxpmFrHjXtZpeo9+cP28se7zpyF6LbzXxhvuO9NtAOz7hohi8M9N3Q
jYlw70JEiULzFuFOj6/wHwhGBBthLWdcyLY/0i/vCRmquMDvOYfJhHO7gWeZE1e1xoIR2JwQ8da2
LhnVk+hp1rqgvF/RfeY2KpdNl+dwj/AV+Dq9O/2b2fFSzKYmJkCJ5fBLXRFUyX9qPt4oIcQSt+qb
iKoDPsqkpAXesGBQZYLTVXF9QgkxNwNNhzkslzydzjYCmzslQ8HUuphgpYwhb7r49RzkAY1Q+eva
dueB50ABCJTg8ALnJy0IlUibVNmyzI9eb+jx8bUBjtYDoP2OnyBbfaNfz9MMNgTsqXvtHquMzxCT
KKwDQN4QJnUnyk290gH+kjD3pDMvxsDCzdzfmGL7zkf4SkOd8Jkf+tjwX160JBvCGLZC4X+y2KTS
KBH0HUs3vTpWo7KcTZALv49kc02tSzEKYu+hrp69pn6iEa9A2sybCCR9SNsihuz1rAf1gx3PPLUb
VMvXcqicg4hPJ0jxKpT9utfa7rAobKrGufx97qJauBEXEaNITLB/qwG2ehDDLgnaSV3l41+rNS4j
rudPSH5z6IVLC2P3w/nftv4Zvz3dVma93fjnKjyRvoCTCgokdUvC4EBMXJURG2TAuWnrOUIDiBS0
mvdNr1Hi7hf7/h/pG6hdUJZaSMT8GVaMEKi9utogM0Kyssv0jTfMal+5j2AfGwvUAHG33xkLEheA
bnI/qgw7t99/ukbzs/Z5UEdIHFf5tDuDv4zbYFwLD8SZ+yLF1/S5ALbeSO1BgnO+7SBhTdNh0ZaN
CAuGvry29lE9jWAM3XgnKEEJbIbwJj7EIDYiJudrA66nmGpSx3lNdwBpLTPCASB8eYzvhLeJoT87
fOgNbIJ4p8KmrHHiBv6XKIB6PhFGVB12NsYrtcv0OECi4j/etW4DGkEfbbv3SCUi6nNuk9lf3Ono
IHCoEjOU83aNGFXYbu5ouNOPX3nqP71IJnG/weWfXusLm6NJuBYCeKPd6yE3bWhcv+dkajvJ1KCb
44Cl31f9Ivn1mGOK91dM+awAW3ncodUulwqSulV/B+Xo4jykSaIdIjsreZz0e2GPxxPKXENvcdx2
HWKStJaYjLDNMvW0ywdw3jCCwLBMSBg92rNHwRwn+SvpyH9osY3Q+aG3tvybO4T4mgGvGI0zwDCA
l/lMq5TX/pqA0gPlakPnRHc+UJYLj23/ulJHSq4bAYlYNuVzY23vaKlL5q7ANd/bQgJQOOZPxymO
1AJzkwbdATO46eOxK0wVi4UioVB8OpqhpC1M5ItSoudLU3BVmtfK24S4Pe/QLCaAASzy9bjuu0xw
ENE3W0B1Da8qTiHh5xYYoGQ4Tgqaf1H8VE7Adxbf0zEa7YghrR1LFvuFbZBgxbd0dhqL7OAbY2EA
nWyA+bsyh2S51x3b5SSiWVCqX9IEw0YK9A24VRkgjkpw+hBcURyEZot6Y65ST+oMHbOImf7+UIIp
H1D8Brx1nW+36x5cc699nxrxpV6xjFsMe6kCfu5h2NCEtGpquNyFLcvc7RxmbaNf6kexMQZhcqDw
Bes2HJqt/Q32kdZnjIFj7dCNcFKk34g9n3BRS9TFXeYG7mLRxntEoih+dOSfNnRi22Rpdqey25Gm
ZgHrSGp3nlsvwMUx2k5N79QLfHy6oQmZKzXyI1KFKlHIkqMkqQxHxUIFHv3NE42ZfIEgMBL18OGu
cLI9OjM4CQ2DS1RHqaWbvZ3dEawNsjpNS1zezwlWYlZN6u1MH3EigSh7bM03X+ZsvcPxElSJkJ5z
CZoWf2/cokV01cfvrIX6uxdoP7nVLZ3goLU4IJKldf/fMiFAn+TINTzGUj35KhSCbb9FTTWuoXGe
YIRUuznHLMnJiN7gK3KbxfqJBPJ9Zy2yzKdiO95IxIllg1DpvkE0ZiHYXOqANoDfY72aYQGPigY6
rxU4P4m+BUTqqqLijoPOOD5ozMEo0gmkqKMnitJrES+7FsxykcssDhHqU6yuUk1XT/IJgmike53E
+jrquTRHrjnApoqa2jD1ZgGNWQqdaOho3mR8od3HurptPAbF72XEQQL0f3YNRh77uusNH9HfGUKH
D+nuPINJMS5cUZEk5rHxwXBfk1O0gl4YmrBLvFAiFZO//f3dSTaAsp0fV49JbMN73UoXS33fg0YC
CHwFf3fvErhbGTfKIdN4aF999sRJnw/De4p4ziE1YQjfM1Ox3IDWbrpemgseJhXnbV9eUhzBTanF
4SCkLNE5aqwli3qX4fzkhvi6QtYUsdr1V+38e3PmAgoaOymBt5gxWOylEnkhROFIMmj0uQZ8gL0b
F3/SqOBYc8hDDyM/5PAUlBGwzsGVJq4FCI5ksMfnp/Y3deipPT4+41Vg3G7JSnhqMM6hdcWsjNHQ
/IdUeQ42P57AADMrfZYpseRfn4Vd6JyAZIUllQUjVD8kAVxbkU9vwIqPDfr2mdW73BcYgw+loK2r
g4TJTS1MG8+pRVtqYICpSnmlsoMe5YSTJHx/MPQeDLXpI1K3/ACMX0nb0D2wZLhP1ZvGNRu0cZBL
jSHVBOIh1WOlhkOPbewUH2N196mognXplz23hMrJyeq6sZTpTBX5fR64WTouEoqHma5GwW7KktQ4
6GUmopNJOFKM/qQUnDUKgwmIXQ9pJCt6zSsNhgRLwPNWFXtb0jhNgF774kusKxBacMQ6SIDMA1Vj
UP00qUG6vMd9H3wKEspyKstmoIhPSIatrwtBqxrj9e6UxMc5Tp+Y7db5++bpnPZrEzr56jr3QiWm
KC6X5Krszj7mWmuyZjz2nGYiQVavoPeNt3FSK1b3/4LXsq6plnjjSIlQ2wkWfHuMy8JcmzPoxQI1
/M8Xgy84ch5voWOZRXe9e6KJf7Yq3+H1ymd6tb0CZs8FYmL3WaFAoTCbFMZRIMllUdgPANhrO7kO
/hsz6O5Sf5pezNH2XsL789mu6BSteD92k1CpgY4sLWreXFrkzLle18YLbUJH9NjnawOPv8Stu36F
OE+2IFoQMl41IGrg7H7iveYMOLhAmrpnnTVnNlTok9l6H9MD4EzFAf9Q5iyjxBCPXhShwOd2DvjT
bZcr96Cl6+DChRotWuxkysx7q/keWYfg76EgF3cCengtGXCmHz0fFX44i0EZPQJcBPYghVybycd3
VE0VHYmcqh7aZ6ITRwbp3FWt+PlysAa19VCiEtvyioc7r0LEg3N5nTkaDMbIYk21E9/2bQkfzYSS
U80W/1cRsdxaVmmOeT78/1AAtI6B4rwsbb6ALOM4Z0haT0ulzDDXSzhT5tZWUqDkLHHbqBzyHPWP
D9ww+qeRjhhFYcAv3bZyStPEnvKx52Af+9+Jth5OcOcZkyezYDRopHMzQwidBqL+Mq3MGnYLTkgv
hk5CnSqL78ifcXcmTS+qVgx4WtMZ3bMe3+FGsz8bu47c5A079UW1VC33ToiYOJ4bR3mjNVKyNw+E
jJCduRBPMVHDdAWgMGD2sOOeFXXW4q+YD7qoCoSmYP2XjgEbW5Maf3X0DVv1NEyCpoBm7vwUhaX5
DIdF0hrprjipTFeVwqAXDU8LgdXTDFsMX5BxNB/BXfl2Pw10QAfrZhYdnopwu5IVa50bc7fFdxzp
TnO2PWky4QMDdpjg4sSWwdrA1sEO2ziAKM6Zn7LHs28NdSkgAqZwSQ37B+mFJ661rp71aTyyJmOl
zi0+MmfDUy7puezINaapgPbcpmFKOWTq4QFQJipQR5Lmu72nmYujMgOVUnoZmO+Npd/+MFpshsgm
eFpSG7z45PqRbZicrGOiT+VUqlHtwF8bueIOzErb6hMZcOitdpVQep2XgFGYWwX8dS9e79v6jCCS
bbc07cacBPZ+x7VUd1l7P8qbCQMZ/t3nEUQ2hXtzLQkEbgj80ETD7Mevotvug6gqVCQ0SYkofN6G
MwD0UthpUpD++olI6jJWBg2V/ovQH/JN3ZIjlXJgSuDCtFDyIbH7IRd3q2Cp7QiZbhnku97EmxA/
qR+U7b7+V+Ep6ERtRPFhxPbeJ4GfddK0zhpquwgou+O5FymJ8eIlm13YX0EeezP5unlL9SNSBcyn
K3VzBTwN8ibMDa6y6y8UNj8UXIVXJXlmqu7T8uJAfJtvWBRF4LilSXKFqOEoJc4DpQOxmQkoy42b
872texpp359AWNhH09AZT0AnlmcpXBIk/cIhFQFsFiOMq2P6EHmlgqVINAyoYdXc/rYVoSEH3PU5
Z1b/XxHBCEFvopnGh7W5qiexaZzZ3Rjc6MrzJIH5H5gFP2BBHSdMBku01c+wLh8+jd7DqaxLcRmR
Qd7/fKd9g4mY7DcEWo0hXNQDTzDpVatIfeYgHhYXYO9oLvV5GkiO1zLreXIQezyUHsLB9r1syvgv
jY/jJzFv8RTl3+ncOvlRl4ONd2OePxBEecaCTXwK3BdQoTnVnC0K7vahx/lsm1xvlPvNrtVh9qmZ
gElwiz6a6J55c1LoLQrUlqVBGgBs3KxoqiSdTR4nkISP8KHHZzAZ22i0mpK/ajDoPWk2OLsIpXeq
6jGi8j5OWhGLlUQOuoO6e5S7GK6W7mC7H8JPWXyiW/V0EdEExmXlHS1stNaexTJYUDHrrBa6LI08
bamb2cgj8/b3kUz5+iQloG09Dhv33edA6nXCV0EgbvOw3jHj7/GukSRwLjPq2aM2W5Asa0w/al22
+eGIDK2n6+o8xKFnby/HxWUxWon1ob9l7ubOJtz8k3N/2fcW4yAzNm9iYB/7LwOBav8R28Q9t+bk
Fg17bm5VcE5Ss8iyzalheK3dujdAQnOydNHuWZ8RXB0mFDVXO4ug5sJQxeHZbCBGhxLCZ7jIygbT
010c9rY5Eh5idS58C1XNJpEMm0Qu0niZMzgW1O1iw+Z0b2WSu57SvGQNET0jAPmC0+nJj+s1sWVR
fQySCbXtRdfxderxCqixBs5N/VRI40EoLG/JsdvppEyQuaV2DZy/FTBF6Dq13R8ZTPpFRedE/YMA
wbM3w2umNhwkxu14xlmgp0ZmgddG2nAAqWZqrDsXWHNSK4SnAcJ+GuDkz/729v5/bI/JJmGu49kT
wWF5C0SxNyUa/Il90Jyja4/a74Fp7c+n3L8QQLHTTSIBz0InKUnK1z2kSLLWb/w5EEhg5VdP8LkF
5v602ns/gqkTaF7um/4VBh9OvOP5CF+qPyVUXVS5zJj9NtarmKPEHJVwA7xBQPUBCwNoJFXSEyvs
eOiPjD7UvZ2hTkyTp36J3kH1SlPS0tKYFprv9YZu5uhOBS+GGZVj3QDrP30YJzDxm9M8Tm0xblMJ
TnGATeTScqKtrFCiOD8QgSAkSN4B1PqYIzNZtifCrRXQhRn4cRHxy6gPTGoPCzjaJXXan6q79Q+b
c2A0XkdKfccTs53h9Dm2/MYs8z1cMuzCpZWvdm+ujdcEiohHHMmYPay6qgqlGdwlen3Qs3/CoZ/4
SrUmCUlUavuh503j562msuRjkpaXOQ/nkmq4L1iYW6PPjva8kshJ+jVOShxlLAZThe3fcl+Pf5Vp
kXFlSr/P16l/HuhDIZIdK8LMrDxWBm9l3svNeQ8gCPwPnEV4UnY2q9lS3t/zSiZmUUxLqj78Vkcy
ddjl0mQI5hlD4o6ZQBXD3RJIH3HAquYSsnq4ZYKuX+y5Cv6DWuWkMfZBCAttp9VeB0D+rMaFrGyF
MHHE+2mcEDyjI35ZXjsNo42X80FLCdmIQbrjbWSUU82fNTmABofVBuJ6JlVY2noWNbfDK/VETgxp
gx9cZ+JNPUHj8LJK61b/8xz/Qx69wckrJXBsx6rYZpzQg11zJs3fiaFhhPLMXN+sgaMz+e0QcZLm
K2XM/leCJ5xzD3vnK3EAsEH3AWoS3t/DeYX7iGZY4+gh7nklOZR7C2qUb90Tj41MC35cKFyJGb7k
Zt0flxrPR177xxBMo64tjcenXBE0NmSoJ59DrXXI0LTGBd+2p9+8e27wXk5c3dhwBfwfmfEAKeGc
1Q4x9bjPbSazS3haGHgDLLuHaJPlMsZKCXzHRR8SuM+yNGEBsgML5gBR0tHSTCm2cbLm+ivuFVuR
ncSBY9q0I+iCgS6K6lAqZ+IUpeYlPh1V5/6ElsSsFul+EvKqNt5Itgd+0OokhJp7MNM8QZOOME43
6qdgAjJ78h665ST6YsVW7px17R2x/IMFjqYLB9V0svTuipRmmRknHdaZN+X0qm3Qtd3D16iZNyuE
FR/3GclgFXLEIqLGf6rj0iGH53Y4pUK9aRH0Wx4oYCcavl5EiQUR0oUrCorlY8QulUUCzRiX3LsI
b5lLSC2UT1OInp0YTBSFY06+EdiT/zguuN+6sk9W62hOXPwieFUSgBr8VWD6vYfAo1r0B+rJ5GGJ
ivcOl/OFNLZp9srKEdVlWpADHj2nld9eFxztj216pWZ/zl+Fgx3Aw/ii6JnACMPjdqRyDkeoOjA2
Y3Slu2AB/tukScn/Fz8ByNI8NSFuBOxd1NqBPVj4JhMGUJzluZoQU9d18yud18H/Uz9tYAw4yqV5
pwTOll+YEOJ408SBHK9tQzjZSpZyiALLYXrJiPJhg6ibnog+CZbXNjaFsEc6v0kt7EC0N5p5ZDOL
XPyYxl57DBxH9c4UfvVWYg7uxrEkQdJFKBeLFCtsTs44U9H1azu/k3bZZvGMSI2BoJ5FswkUnQSy
VlTWiEaSrCEMQSWZIRLQmZF/Lfh6Bgy3SpTWSbAXdRk7UvQM0EQgvje+LaaeBRo6JPeW2Pti9/rA
atnsq6URNNA0UG1fX7grPxCB/nAifF6v26aZvmkxnxWArHRTaKMuQrxQM3a5NI5WOeN5pMxxXVAe
IvEp4DsKI8hBCv91eN8juWMRuAWJIz3AqA96msBlfiBH9IY944okTEIcTqWerAqm+FWe9hj4jCqr
NE30lGMzj6nxmWJkqTaDbsCn0l0h/o5H9TCE2Ba86I/nFeL3tsSZERmy8Vs+cD4lW866YgpRAEda
o8mL6o1p4UhV8HqL+WhLoOeJFIpzYc8kmS7qSQQQmews6LLvpEmYVfKpAGsfUgqsYvrAUhMdRsgd
8CkJZgguaaQdYNqqycPT/znOBZgofDI45VCwi/X89rWbpt/duPU4BGfpzQMNYWC48rmpICHXlBG7
t2LVznhQW/XhP3BefAM83R3bfBW2JspuWvmhuy9OECK5dmt32aSmq3G3DrPiqy4+m67ux7lmArVm
3XQczzwenCHDGasIkQVnKFP0j+wKyQREq3LdEmHrD4stFext42q1xpN9U7m1lYJNL3RpSFchEMJk
a6+/3aZ6v2LY3zPikwBZNfi6/R/plBc9FJVcL7GWTu4Y4fzDqwj65WMTa/HUQiw9MYXboaQTHGyy
zOgBnBu8oCtKTrKSR3/BDGFbIADgkczL/EhQyQyxZJyRPrJScMBTA9ofs7dQFzrLZbbwUjEC0DfW
+6LiZK2HoG50UV3F8IvSmjZy6T8+Q0t3jECNoVkT+U80vhfKYuu+jwG7pe5e/DQ01moajr0+4Vmn
W7j5KXAnAv0yNgVUgQUvL+g8n+Ct9Patmms1XUrqXGgCGSEm0Z+8auU7Qq9pyhMl3s3HZPuWq33X
k92J+TxEWfG3JUIByItFRn8hMPajXEWP2pa0SZNObYRMUAglKK0sHqwl22m1qzJRHoTOMrl5qVzj
pRXFIdDPnZeZq92mABASCvI2tNS1A3Zs9HsAFoy00NR0c/58BEF6+Md+yMmNG7VXDxsNuVUaOfJ2
bhd8z3cISzSotmKxfEu1241TqlydhYZpAqFR0cWOSleqYjArZ3Z7pQGF5cIbeL79a/O8ytpKf0bc
QED1PudzyTc37zNDE+ciq0/KEMT7MepInllPAQ/7PvPFbq9hnb+77vk2dt1xiuTOrWIR+9wfj3Hr
RlukoaZItzboDR8NAMnh6IJLrs4OcDJ7kzjqlX1/AiiSra7yJlYoxlBN3EghqTFmB9EzeH6uzrkK
WXWumV2FZMzDQKBoSziEwQpQ8YytS3U/bEMt8/5HkaHSk8KYKSOTuqBEJ1sFsLNGkZTCbc5VQ64B
A6az8BjrZuoHIoUcCNKl3AwOfiXGbHXTdPYHQn1hpLQvIpxV9nBVo/W1aMsPq74ORH/hiQFPmVct
kDrCuKC+JowyOJJKs90YHVNFJ3eKbYzWre8CUpuRLeX8z0BfedDw5PHcjzWu6h5gMcQ0/sJnsz4N
tnVwqIoSWEN3cpobgK2lC3n+FiDGED5rXs//wyGaU5eEoSKYk+Ha7BDVCl0MNGy1/JOK6eFhEOeu
rw7MJuMbQ86Bgd3eHZqhfj8tIVI/O+oDYnWa/w1Mn6rO7R/SVLu4AMKa+h3StM67UWXSOf+cNodj
zlzwEsEQ0AjorL2yDe0slgm8fEBk/VfszNW3eYosz08n6L5njMXexbL47vN1FI5xMR8DfsdLMZf1
bfGni4R99jarBv6t84k4gxRIPba9jBi6I69V3BIPjdeNWAb/hoc7c0ldyRxo5HFIuFn3auvGD4z5
seBjxPo180nWk+imu7QshoAYwQb9p0QxiR/sLxVHZERqJI0Xf9SngWvmRngE+65W7AK+ezDjgwWp
f40IvTx2kROk6dUfLjrd7hFTmjFU4vYbW3HHnoxCZ1udG9A4LTDxCMnBHbFq2Wufqh3etygYXP24
cFS2ccra9wD0O9BWku+V3YzDaNslF7KRj5vwnDCXDnszO15SQHGJk8uS8XW8TghPnFkG4RADIW8s
gGCj+HyZ9U4o9Q9ncHMIAhPY0LxnMytVPDG7QdDPpMsHLuKH9LJpYO4742OQocnl8EHFw/1tm/El
+kwLZM9LtKr/8WqLqyvPK6igBDgMMEPNfZD7r/A+etwGUZsaxtyzWnvyxpyiGdkekAwCYqHPULF7
8D9Gy/4SzGaoKF/OHslRPraytT+VQheJJd+sZVXXoGZ4/JdqhdTEYaE13/RmplEw1Oz01m0h6HR7
RTnWy6ezVhVhvhpYT/TBCBxQ1SH2ms30OcuTGyAaP5ipBO43akkIoJQR/iwbz382+ho3YrZe/QiN
SL6i8a2oBGoFxGhnLgGTYev1JI2nnz2LF/F8q9uglaM+wzMJaG905fHP1cScIFpOJcmnXFDlVw/e
J3sbUtMjhucIpByfHR2wlvC+0MOR/9HPpjw5vnmiTXaKDSilF0k991XFpPuwNQxZYhw4LCVklCeX
mn/fdE2NbFcX0Kqej+jCIbvimFJmHL4JzcrFiRo3nwtwfssRo0GBC0E0GRfVbx2NxkCe/Outkjc4
3QXcLLtMaxafX6fMLHSLLbSiVjVNqdu7PL+ALx9/Ak8MgY+YtZiS11D5B9U55vaVzCpb1rIqUtDU
U2aC6vctQyd1aAy3IgttcSJRJGJrmcniaewDcrVnwfOEVBonbmLK+RXuQGShvNlljOIibGM+QF1q
R5d+8/1Um568Xei4Xrlb1rI6obOfrVwgARDtHl7jhQtCnIkEL90/M4swCtIWqAik9GAHBBpozVR3
SWKRcpLXMd6+KWaiEjm5QnwyRbMgwtn/HKFr139wqRNKnMe7gxVSJTkdQeaKwcwVT+C3zZRDr25o
uzOVhQHFFzHk0TkoF7lsJlb9XaXC/LflrjnJF1tMcaldR+Pir5ehSC6KmKrHodDc+2QfwjOccvPH
Mc7Xt695k+fO3LOyJ0ncOHoDHgzEVVL8swesHi0In53mSHhQZSUlOo4CFtdzI2p7Nz35VCEkVogp
IU0T0BDadwJySy075XSWtUmBnlPe8TErOI4dR5Jmk3GYjU6CbjOK1LOLUwESn84AP3vifHzYkeUL
TFUc7OqQIVWVuVf+YLmeQI1VyswyfuyQhmSRYI27Ke9kKNDTopU1oSex2jWYG4yc/BWsLXYYP/te
tc47RXMSeMKAYdhfYbocCs0Szgq8hZmwp7dkZgOhdZMOyyhkKOLVc6wpE2xrdjFvLog6VJVWCHub
CEOboYiaQG8kJA+OTFlCj1CeDtbyjzPbCS16m9uOYvHTIQ6VH1VWr8V2gruU+aaIXIafSTOMmjJb
gTDHE4klKG7eHB8nBU7YHDeHrbZ/5TGONjefesuv7CFLysyPfv00ttpLzCQw07I8ndAzeiiLGwO2
gmJBSeAUQ0Ui2CX04OepRlZKdlxcE8qZAprtOmbXbKL9++FhzIN1aTqiCXWIVFEBgvUxwea+lY+I
O+nvRvGT5iN3oNQkBohES236S4amttAj+PB4ptIBtZbKFw1PA4pzxPSRbAeSFjpUlIhev37JRNq1
TQ64yv4fw2Gy3EYW2nw9LDqRfl+lQSV36lSrPOJlpsDR4Cac1SuwXYeVvt2885N+bnWC0Q04MKin
PxVG7WEhfquK16Dmreryae9l2R9RsQmrWq33tf6UNpeYEKzRuNJU3lqpOwXnDyBPQYrPcI7K4sef
WSfxjtTq3oDDz70QhkNCiS97oTvwPIUEsHOHR+ptNi/xX4rOmSLvNH6hMXi83dioDZ/DyRz4Id7K
+A7oQPdxh7MZT82bFmn+mTrCnSE68tkX1K+6rKp42dLMTCmDfZjOwkfYRS9+Y10cE7lFYbHpGOfT
+0JnJ0CKDGD2vSB0TJcnJtDXmNcLZMayzQxG/yHpwGeS8GouKdXqhentVw9Q3L8TBnmIkLSiq82L
40a7PaLjdzO98rLq+2Y6bqCr88TO/75eDrAVJJyLlEhHhdumx/dqNEe1NuHpAya2/XKoLWhDB5m3
95HIojplh91gFcYC1qnrqJa1JI3NtfsOzj4KCTTIy6poW7bi9BJQL7rfolBn97VzpRZO/kiei9qa
dyAjI+MD4mwjEw2TKOKRUu1qN/9Wd1A1Zy9V9sqDnY38cz3EVV0UE/sb7sP79RWmW7d2W8hx+n2B
1d1SjRb1IQObbdl60R2RBF8xmogSMQ2eCiBBLWvtSSgrCrJue55oPmJ8uk0Er6oQ1wJKt9ABh2Pn
9AnorRwTo2Wrp7Z72pI/xHowKprpRvAR3c1GaxevhfernUYt4159aQRTUfqjQoem6rHL0pf03rPO
p/U/g+VUus5IXLIcSyL4xyeFoe+ujodtE+GjnhkxjB+T4ptvfIQWNkbf442b/1hEyTcGAY+GDfe+
nCuW+gJBmu2yrm22VRzQaeC9wEdo+E7kqlt12cers0drJ7apiakn59YvpYrQaZmyGzXaCibrQol6
m82CVpHzZ88yY+bbHLy1N81PxGjmqMLvVHnLPkMFACQZcLplUHReuiPyFwDG+4V4nS7HX4VyHYHE
Nzkn3SJX/1WAYWvwXw00ue6ZubU2Nuy6Ax5vKMsDGxjGHHMv+KJ8YpYnwH1D5ZwF1zvdo+NIiaHZ
8zArw5Nw2Yel1RqmAG4zqS3+wTm/ejHgd0JwZap7GCIX/S0hBU6hFpsaIFFC5/ejedhTEUeS2Y/Y
r43VaTmA8f5AxZpNgBBbICVmlDhV6tIPmN5pfimDOcQI4w0LnTQkpIMNnWY/iwridgov7vH9IhmV
BRftQ3EfP3tcJ7wQWM80sGs2jTEM1o8aa7OFkn5opofDbWB32gg2f6Bz53RemWd+axtGOMIYCFSz
Mf1TrwKY1mbQV/GrwnS3+TsVY9jAGwC/+2OtEM4PMJdnTlG3ygvGYDnVUENQ9MmhVhJ4micnpBFl
5aw8mWkCjTZXYhGJU+N6jxlqA9O2jq/8uUarYd/KfEi4DxU8ceAhbgDpknStkNaCejvlDuOmg3BJ
GYkQ3cGXouQ2+/pk/9HenrumR2jEU8ydNSqlmeVOm2Dnab1+83dLdWjU1EVWqD7WHWEl74Dg2yo4
EwHo3buhduZXc8SlKEydyfgx1aTEvnDJCB77JTqWuoaSz5x67Kr+Soywyk1w9bzLskZgAJhPfXzS
HdnJ/Ip5mDEO+L65iRHYTzZ/lcMUuQ9Gga90oL5N2xSRY1j5BqdiuQjaEAu+xVYyalwkJXDT9Pyv
/qBGlzyZO3ma41BhkRIHyp1T6uGGvCIDIB9NFBsD4tu5JYD82LNDXGQvnsxkY9QX/WiWDVi57xVR
ApfDPgmlGlvKL+H6nHJTaZjUyk96Ihp5NNU59f/i1dlyxmU9oL+WE2sRs6xBNdqK9G7YtGh1FlOp
wECfQR5iGVnlQkjZ9qrwtyGku6yhQ72uuOOtBELPJDrh3TrQO+P9eh0wNlaZSsEKXmerEPheFDN6
4bXkHUunR08D//3fFrbTm6jE4fjZYgUT/4MaeSLbh9c9GzWecjjWSVPhCf7jZpPHoIOfq7vtFPU9
rTga4DxecRb9FLPTbIb6o8/Jeq5t1ESVklOz178KDV2LGfRigy9BxU/JlJPOT9T8PkjA6oJZmlCp
jf21OiCRtoHtpmBcvWh1jCXThUxIcAoWpg1d26Q7nDu7LNDGNmjMdtCu7x4fJysVR1qKxSdSBasS
FvMr9cW2qom1FCUEhV6SMPpswmaI6/KLOCUh9FnC0srZSA3ifa16tx/PS/bUUOqmaaA+x5jHcg7f
2L5zifmJZXz4uksUL6ufk1vK1gpSQHSEV/XNklFUYEw+Gh5tQ3xSboBC6b2g35OtJNEclVriW4g6
gkQlfFNZm8VfaWXiN8oZ6yPrbVU+ADUaSKyMD2cI95g6hu6HUhC+PAtONrEmqOUnwSLGPVCN+v50
kFJQV3k9kJ6AfKx5uolbD4Ni1m8KBXocij79Ix0516T5Ly+sZooZhUuZZzJnMyojSeowQJKY2TvE
+JsNwMxGvI0zskZ3d3BaxUmnyyp+KLVauYJF6bOggycZP3+m5NosQzkOKOhZt5QMkMlq1v5mLow8
Ci5MKpoZ5XAukQM9T6iR+onv6NY1eotb39i9UDD20yYs4PoMom7bFESzvYGsiStcFma1XN83j7GD
hO4rKMvsyIOc+UBvqUQpoyscTF4Binvjl2rWIK9xPI3NB/2xs7RXxJ1gZA+X5ZNc9dlQR39E7qI0
FPJU7b43XGqMZX55bSnAvwW3hCQbC7hsE+Hta9QfrtzF+7LkYHpeNstzZLx1VjvUTQxtDV5YDKGJ
vlEtpptL3rTiDQOXvZBVZrpNE0i+dERhtsxshUY3ckLaVPP4uCjBds3Cxh2QnGhF335+pfAoLy3p
Q2SL+rnED8nY/YOmSnG4zoEpJctOjjx5ZVhPfMV0b4YogaYZHz3Xf9Csv/RBXq55Uf2ImdTdmCJ8
M0nqYxCJm9OPJLgHZgAhRZNyHwJ0+DfXEaPQHcLdxKNOY67kiOlV3ofZM3ICP7cQs2M6jRoqYzsW
swEZlwZbqXzsFzNfVhkLi8n63JLqOfJhKndzFyCiHPxQ/3XAiP2JPxJyFfB6NpTw+IJfgsI0NbEi
fjWFdhMuHf1Lj2QUAccfFgLy+SJWtfs2A7K6L3paciE506rCLD9NNX8XUwjeMXoheBUk0nSK1bqX
eqp5k/kd+e5n1nFX+WUg0cN0XQlTyYSnX3Qzl0NA2SEcckaUrSjF64BkuABJm4+bJ4+9QQaR5DgT
GO5kGPOcymmIrp3EBnJEl6RbQJMPot7miqXN83IVZ3j1sGUjMEZDeTf7ke0q185qjoIGcwTr6pAS
R66kSbHt+QhdOKkt5JC8wSVQ1Uz3y8JN5+xguJHJ0iNuQzRwo8qpFgOtuvB4ny/ac8nygBbEKwlS
5frjlDnVEHnRy7CzXXuy6DQ8BWYeV9qFfw3t+FYIpP13P0vgpZ7fuVS5J2PprHOVoarbcc7nkI3T
QEjiJ9k9Ss6EHQSs9n1QxiiFM9PZgwl4QKEb1r95Qits1LJzvyKQL67Gv0N7QTbh+GoJcOjdfZl8
vSyKJ1IGZTRiO9/MM/ElR5mztwNRKaQvrTuP9/dEn9rrLFCUheaeJz5C3QU57lMKirxy0orPooyo
SPL5sjAGNEaludFkN7/BW/tYZZgj0VYFiWZVBKr+G/fEpky7sjJ5qN2meiTHVLFNeOMo+xqj1o21
dahhCBf4Oko78d1u19/fgxwucEvrmAm88Wc4qzCSvwi8hj3cM/NkaXBlBzwNWxh8NgKokNeNJC4d
ARi3NXtT1mrTZOakbv5sAGx5ioBh3+9h3qbTaE/nzNR3vFo6pmzrpygs+5YiBcIQdcgt316O6fUe
+oaUCKyXM0sXDHMCtIAk1YdValPs2dY4HJo3R1fCgaO+dC5Vm3vYhuyReP0DbEdJD1ZXDT10ina6
fwq/yHkuBojQtwYTqW6OMu7lTXtwSk+GrrJEIDa4mgPq6ilFP3qDH2Ru+MaR1jOrQyCOZV1wa3g1
zqWG04ZXeIf8/eLBSTWyl97ul07cEN3vOtYFBzZd+jpM3xH3Y4ogsTfk4/wZz9YXH+obdUXiuuEa
Iw3q1Z3XZzZ5PkA0mFNfHK+YjA1Mh6PGjNpZ6KU2/9MftUCLHXjRZGGdx4uniUQGMX+6kRj23yj2
SrSgZWM+DQGLuDaEz3lMShPn2qediDzUNFRY+fcw4H3NIuFxLPQhhQwwcacZgyhZadj/8EAya8lY
rwF2QnA2d4+8vZ2CCLBglFqGG7J3Z22CIukBerXu06DrcEWnBSumS/bRuMur3J3hl2kN1E1Q7SWw
vBrCTLIrqEaoNTKDaLytO9VGUwWa7RCmbM+zrcb5kccjRv6MNXILvCQ3qLPoIsR9Q2nt+bmdecvb
7Muni+CpRT1AXt6pbm8fKGfJ4e4xiPQk6jZWdORz7Nr63zwMKOf4bAKpUtUaYQhL5gyyEleYY/0c
mYWf2Vv8O/xu8qDWwr5qB3RznPOKC31pQpRd278pKIzbUzjTu8RxIICpt5d3w30EKwiNcEC7WcVn
m5xLUnZAJPhSwpXMihJoPocFt8oOBvVWPwqiwUIyfTJmWn7EnmbPlf7MkMGVJknnp1ooEvgu/aXb
JaWon+JANK9iOccKe4G2ovlf2bjlYy+W65r4Lq26ywkarfykNKUyMqR5XFJChsw65T5xSaFoTuYA
PtweKLawYKbLoQ4kWOWSAFXLjmy22wJ0/lHoHno/1Tl/zCn4Z4ghDdEJSdujGjFv77vULAfguMHI
BpGWIUKT5LwN5uWkmksJ1/s8be8KM9y2hEixNWLeX47OQjVm7ZfKkZ1ClBGKWYOudishxy0++0Bn
N2D0AWCXLkRKLmEEL4uZlNMg4ikpH4UBFik8/v3ZLJjdURKMvUZ4s1zGXQ4vIHh32ERYED7b8vCi
JIgKr/63Wj3cN1M4ZOeIEHDpsJXeUwurI1MPrymzEN6gCXDwj7IOJcshma+klq3uUiHjyz2PSp/k
wI1YrKVjzOUQHdq706syT1/tjJk8FjhphTs1t7QzjCMNLKMrsrhxi+FOaHUohun7B1yK1l3dEeZu
o+N2SgFkEc0PWlzG2vaEfa87CFDFXvI+iJMnQt0cUEXDbokSLnss2TV366ukNZt7pKKjLcergU/t
aGtkc/NdzvSDo6dVJEjgYZ+qAcVnHw45Sdrxd04y82DjHNc063gMmZkgDIaCH8o0T4mheH4k+dXe
G3bgp5g4L1NORUmVXk3ZMJsrEl+uJmIMgom43FCHMFesMK+tJU5ZQtAJbm35FuaRag/7rE32jMG3
Be/uOoQfg7bMqPUBNyoLg0isKTjHYArylCQOAVtDZS5QJCsnXS1w+4NI5C15+ZyYKYou+orBGVRc
ZHhsVUKz9+P8cCJ4QrbYOhr8VAM9CMZIhntgbUR4P7vRm3rHho/ky9tSY6reRDPwgOgXcu8bSxAC
tVxp0n30uDFu3/w5a6K3qKuwAJ+vARuGa8lMSjhpgQ2Tmp6Q0BefM5UHSGFocSnZR0g+nHoBCvRW
s9A1iwKOt13L9QOy7E9yuXPEdfR1fHdyW2PqxRXe7Ow2awY+e2qt/2tsfd5S2LUJiytZqpjZpe7E
RI+qS7Qcg/PnXlbee6c0n+KdiSHH3heusstYVM1HWQ5/dWKI2dI9GPlRXMal6dDYrA7bnCb0Ospu
O9ysGfgdfdqOYVnfujNA4/R5mr7wlaN9t05rUmNfZLwTXH1NvOh0X4rOcYTve3hPSL8VizaeorV4
YBRfHb4g+thip3K2eBL0jBfEoBTgrY7EVnY/vOWOOgFtqi6eDBSIZv5deRVmsqX9zyX7qi44gZre
mgDqc5PWpFv4t5RQ9o/g5R//GqQZDSPI1oYTDKqaK3wQ/aMKmVp9kwAvPgJ3dnlbUPKGK8is8Tb9
H/yqkUBr11aJ2HV0lU94Abvf2h2XniJgS3JMVsXcJ+K6g1m/JMXYjwpTHgnIEJ1kQjhIzD9o+CEa
Fclsub/4MNI63MDUvdsPj6Q5I0tYt6B1M9PNqlvHDI6IwisU+SevOW2k//UstusVoE4l9p8sJHKQ
EVPnveuyxFtFuf8BL6LZWr3tY0cASPGvtCRDSr3vhQ56L6TzELbwzts6tf76uKL735euzPqYdB8T
63+gbVmUtLTdtNlTKIlM1HMpv8C1NpajKX3kiAsQum5nqkyZd6P9LU3241Ev2VyUQ4VfcEx0WDiD
XMO5QzFnW1aJXFE1WQZPLA+6s6n078SahmnTiLOmxUuEEvWxDzyRPBmh0s/izlwH51xhl/2EI+PF
XPs+aJIAAtxL55HefUdc7z+sNpuzBhVLrd0gH/3wyZeLfIeLQjbwJzTYC2yRFQwvVgF3rF6PUNEH
gVk81+3MaU1vyXbPW7DdCvOTIvtSdG+31D2wE1oyYvVDxuAb+PmZEO2exl3YtpSPrL+eSeAHscU5
gGyC7EgMKPt6+m1vz5qmwIYma/8+vGs1opbQHRiG3CCnyLZ+dUsPkjnQKQIRMCwjD3kJogDVUd0I
dWLtDBuDfM0KAKlaRN4W7NH/p3DJNuzFoGjHNJmyjiwczZSzXj+POvvzX/I8Kxs06oDfEYKXQQl3
e4CIk14q2oXD4zywhViK4HWp9mI1diOWDKCwGCkL8a96bG5sWLmpn6VrgwtpcY3DLQd4ZH0bImLe
HtIPq+pHceuLd41VeIkSF/mehHqLPahjVf0eFzMbD8zOCV8JCIywtAucjoDJc0xbFhOzA0PhyBAY
W4VRefmUXMUBrK0ChaImfoq55/za7a8nebXCJ7Pfjvw6U7LYoE7GQBs2fLxrbMG9ySREoBtRDzkd
yUfAohAh7wBExtaM8m1V9EYv098umDtrjnXCyFbiFaP8Fq13y/3X07kWnWpbFM+VwJs9uolTck5g
fLjIeGZ9JQbH5KkNz/ltaxv5Ktbh3o98CktrCCqFJsdtMobXPwz766FFUIGOQljNV67JJYGiRf4c
5EVei6H+z7Kb71Z2xq0ALqIdti5UKbHZdVdQ/AUAKfDyL7yMleln2YVo4Iek5LCm8AcJUEmyca+0
ePAhbVAlPVgb5yVBQ4zeeF1l7AZW7lXWfytHJwVvX7e8lXZH/Ty16bugBv+H1hriUqDiMBf6glST
dEhSh9ziTbA0TDBFAVZQxB54vOp5ELJuXJKPB8Ba/EW6iO1UuSrhxN2gWW/JDRlKoradEAPopjyC
uBjkzrCsAiWHaHw27yj4/7OaEla7Fb0sd7aSD4NQ12PHedonGFGz3lCL/espRe5HN7fRAbjtuhgm
aGNA7l3oNHqoBpt2jgUVuUE4xf5J3OXHP5h82EabuVweRi7KmBZeVzNvkGx4HYpCgyf/Nx8CUbyA
V93jZIKYjczmbXucF21oXrLnpNLh9qI21KDenmClpFvPSCgr1e2w4plW6cxLO2sv4BzDzYKqdOAr
AygyiVAzrZL7eaTGBuf++zrcrfznqpXp+pcXm0Jp+8d37HJ5JT9AIXBzailrp17u3fInPh3TtbmL
ICltdsJzCIlVAGeazbMM5lRlaLD+D7Cttv/S//mFsXtERPs7A2Jf8b5FjEKX9ccw4xWChxEsytld
EnkWktIRN9S0N5rIX2X/Z0MaDxhZ2d4Ym06exJ1HOX2JauRsuEpdKUPd62/qUBKk5SasJZh4Ce2N
4dQVSnVaWtxUtKYMMmUDabTu3p9za0XzJiPgJu0h3dHcbjhrAgBjz1AEtbHYEJHIPdJNejZqmQpq
h07RychOpo6ObFycYTl17z3cVxXDRKRoG2svaw02Z7qDHiGS5Y80Mkv3M66VfAVMTMUVBHzaUkNH
0X3u4EhB2Odx/wgNji5coHhvnw57YhJMhUspIfqqcX1UjHUYiLeWEwsq9elC5AWqK38iuOicHsaV
EIzsVriDErdx/LQKsbAPydsrQI1SLRR87NwcDYnPuCZT6Qx+FcJS8rm13Pw6XvgH30804ILRU8uv
96LUUYOw43hEXdhmiMCr+kpZcWaH6J5Hpb2UVBbbzmqb8StqffPnZc9LMP30K9dAmQexd9oaw1q6
GPrHaWUCjA21FwbVnQyMpjUTcDWGSY1xXWc3xynRqSjdegljt0Hslq1P9CsnBhfCZ30ONyFuQ7i/
eupXRwbUx7P34vuw7uJQvvMNeKcfi+b3+U/LQwEE1woog0i2XxGdG1N/tI3YHpFCXy+BybErRWI1
uFowlzgaM/GrwKjiGqGBspwEIjOlzFXPESpdgykC3ZOs0smsfDKTd4ifVeEquEOGKi1LrlboAeKn
o7fsgMiAgO2HXclpunaetFOvSygT2Sx48vFlruF0GLDiJixft35+eTzPkaB2In79xxcV6YfPhyrC
NCFZiukvSUaRaKotSySYbnfxEs+jFdQmPdBCncXgQGeObW7L1vN7uVxwFtazASmbqLHayFd/rjvx
P+nKmVVpqVuHRq59dffYfZpYwyC+xk6VRj+9L+NdFheDSA/5fh3VrZ8PNrqF0VtuNV9P+asydNVt
6mEPcODB3IA54s8LsuoxjVYhC0mre8P1efYstY3w9T7F+OGb7KTsL4UuAIKMYPHAWDHOf5qhNR7r
MgTP7k5JH9TuK3drskEscUYqAMlD/J7yvfG9lM9HrrM5ES/43i9u4YMLew5kCpurC+FvJKBqE+bW
KumszayP0ImQC35Fxsm6xQ2FsJi43A+JJvz79sUovZ8Bav2tM2awEPF/qtiKZ8djxDVrWIIE9vmL
K68ArqHrU5HpLoFsepacl34ixeKEuyFRYWYBgg0hGYmxmuxi7i3hSd931V9uKC3KH/cXFj9tpx8m
htbR/A2NjluJrWWYqW4N+IXNOovNDHGTp2Kn8yN2JZUITqboaUO3QZzXvqMcwTcFXBNlUGlUELX7
2PJfKNdyjfMxNX6Y9ROHXAZk0k0jIeethqb1f0ivrF4pZmbb0Ua7U3u6kxLH/MYFYmhadKQmzI9A
ieHtvaYroNihV7wXDp3LGDzITyy7dX6MeVP2f10vHDiEB1ByZ3xVkWXMxk08E/306BD3DR/dhnN3
t3ktz/HUN1cVVvt01lPh3WSBFp+coImss9yuUx5vFma6DvIRUfhdALPL5jZ6L++xlrhlgjkYTY2y
MWKzE8wy/HolHlLS09UZD29cYIMo2YQ9jLP1+17U56RC6wYZcuGd8l8oK4TNXqRWhOPBWDeMMt6X
QuiTl/ZgZOKxvDEUzsrxjg7yj/WnLH1r0hU/ecFk/6cB8pvoe3maTgySB9XVoUiwYgHRigrwEMt8
dDBVJe3e36yuQMp7lbx8sgIlrQtk+SgPaCdcudjq9ta+nAbv/vZdXTwODLU2Z1/zrT0qeky/24Ld
oafRNYWAtI8O1NZn6N6mO6wi29wJy8kMcNm1QebN5/5yEIrs8QeL8iuMzm0dUFqjxsRrSTOwCQwn
YCEAhMKkMf1R4RjYjOt9q/GCBspxCMtCZG5Y/5F+eNXp29OBtfVWESOl1HUIdDQ/pITZo/R3+il/
/tDryr5Uw1c7iKFHlQt2juaZXyMNQmH8zxGj5oPIowgR5d1dzSuAjiR436taU7dMA7Gy7nlSnXzz
umhq+XGtSJYld2t5h5VwlXnjGJmnla1i2cUKlqeAObqBht2nThq4fUYzpwVrPOUDjKowBr+hnWtg
xiIhbU9DpaWmzAFfeOJON5N9Sc+PgdS1gnyZSJSJqE5FlVLpntqAsEHp2DWzNgQM+auooM0/f0ky
HXSnXl3t6gkIzp0BA/wFLDoMOnOG8oqpvSCc3ts5Z4i/13eLb+7qhFtdZF/dTxc6aeqZ8dwb5fdq
7MwU7D2CLGEzynXpHJHn2corwoQ/7Dcj8SNRZ3P3V+GInmOVQGIfPzZh81KIrHB39j06kTnLiIDy
0AYC3QCHNKfm8L0lrc/+5rmpvOzCSQLiW2H/JTVZJpX1LbDS9VW6tZH1eByQPGA2DqLYuIgRtqPY
lFR4ueX2/klVG5H9F7WwkURYOQEtRETA+qm1xgXDhiYL1r8/kHEansQfXcNchXCdMNfJGSJCnI1P
i1nUdM2XVQBIPEEjbfMy8cTZoV8mDYES3vZ4gYZLiQTIms0Oc4P502uR9m1hO3F/ldetSnkUlhlE
Mi0KKwM2Wi1ScQZcDiZJfnWJs4DkQZzTib87wF8Zfamkm6YOpXWnCo9WkyqbOFXrwSYOZ9KsnFpU
vQfiloOMQ8B/DsiZ2ejy5bUXZMYcY3ct6AlQZ3FBb6+25dWAPSI5H1jbYvVfZyVLOAi2R8JkWo+I
QXXtS7zvfgaSBbaJSgPBe5VaudhAkcvo8Yrine992kyo5bgT2pUg050dhhs5N8ywD2VULwfRv8EB
K2m/38wcs4lJhjwcMo3sJ8elNILd19HHY/C/ngi51HMGKD9STD+f+e1Kncptbk2SAzuNulyOXJM0
qmjUtzEb4yjb6aK+49N56SWTUQ0NtO29dPbKJ4gIEy9UTYIlASvBVqzlyOf+cAPGFNWo2UT8YCkR
o3TnlZ3513yzgANHOP493HyHaWv/gskIcycYOMfXJGVI8GPy0/GKOftLjxgzA6jJD9qVGQUAsBca
eHn0iVUZ3mqdMxdP08k6gRNYwshkGveaqF+CgUarTmXLMsqaUdImJehqrgfi0fYI7yIjNexjVVO2
MCJzOdiA1Cco5KvTuJtLRC8FYotzoTQU3d4//65Kxqmwi2KQJNteDPzl2AzB6K0/u2XLwkOwRkU9
b9Y32oTzbS3x/8H9yNb4rDWmuPJQs2/dqXh6kHiaMo5MQXZBX1xt2Yj0xCIPsvuBOoEysL//TPyF
BfU+e4rEkhecKvqPjAm0qxVNgT1DOjY9C5BbUNw35VfFsqLQFlPrEgA0sT8866NQaW1msWpi5Sak
7pUye0+pB8bNg/oW3jGhTyBj/dipYrOY2i5wDLq5eBcPZUhtm/yIEFnOlh+SN6tLYEukX5YRu208
gKj8pQq5ex81VLh109u7YuKBcT/ttz0jDaYdbGofT6nR2iAPNt5Ryn/REB+0dYAULDd2qHmIdc/c
thNBsqfPj1EnxDfyiGSaSpQWpQoRlJr3DMDYUkcPgNa0Me1HtvIdcanFUmsH0R25A7aLWSi31oX1
h92cuifmzgB1nA/ItyBYiwXo+2yUTLzmz4q2RYv0M0Q0OLwsYfS0brWJVQ/mjdoF5KW/6uJiQ4td
Ty6Iro6bqTk9Thexs5Spqtw/ck5KDVjJQrS2/dLLToklNSddnMLP3kuUVqRK2xC1cJMLj4UoRLz1
ABYzWR2Lmk9MVV8KK6mmbMJzCeMPQ1DpucGOy0NtWyjZRghxgKacQCVECMu0ce8jahdYlPrv+Vzx
Y8B+AvmZIlsveu/giSRmVBVDKhDvvHr1ZOB5ioGxbp0gLHguyTJuCGs+gfeItigq/A48jhQ5v9bZ
f1qXN6xXxEtTCi7VaVpdO3an9Rda0Pxs0Gg03WhzQpCxukdoxfaI4egtOn8dL8YveFX7hLwrqWF3
8NGIjS3tSjCK1uHvv6KMv3I2GNv4Br0tdcfMPKMgEtJarm90uanCNCVZbnQigP3w9Bh+nh4zcO3o
ugSR2vit+WezMoOLnehllj/6woMEL7LRSGZz4O4EEx3qrZOkuqdEdc3YBK1TSnbpSCbezVh4h0k+
artske4esVk/7mrO7dABABQfeFFNSgrugnR6EYn3to+e7ugv2PFnURbGLl46VKIq+fMgvUdan0Ph
f8h9V6vzjyAMmdH7AASB/Xa/wDEmwSxG7rn0RwnScaGG/LYXOrz19buv9pHA1/5xPWA5elYVmViK
OO/PaW5Mn9rg6FDrMNlA39vMpnn1OvZidjbs+dgPqrPDErlrcxt98Hg1tUAPQOpQI2SlofYL92GY
MVGfYQDl+KI66M8WzDKL3yl/R3VkRmmwXJudbyjtCu3RCyItQhkdbMUGazp+QD3VBBPjJtAVI1b0
M7zj/g5EEooZyS8OlvzqJl3JL1Hb4BEg9uuJkByC/ArVYL0k9SkovXum//Adqh0jTw4CZwxA3CWT
vawfTFBnxhKTEkFkfxlk2lMoUgvtHwKbt7O9T1Pek6hQpOEBjB8zPAQg5ola74A3lUEJhxaTOIfz
ZK+giutc7MTjwxVeBoxbHIX6k0YTdy38EJ4HZIjd5DX4NjzIeyk8RgJ2D34voriopbDybbtn7RUD
clxKL1GLGKkFev2gtZ38fE8y666xlgePlNqYoBeIZzKP7EmCoSl7acoKls8ylu+y9xWXAx5ZF7xH
rtuVyWXnSD2yWDPabtlepW1ZvgyovD38wK950xe3hjDsB5TdFfZEdhiWL6paNIisgqhrjXY9M/RL
s09lqjI+Pi8vCWDVB7e2+gVS9p0E5b/DuVb3qvaInOlyx9o1wpx5EDd4MPWsy4mJOEhlAI+pr3/D
5zBdRVjXyycNmgTk1IWKSfTGlR0TGU5xnaD6SMTnOGsF3yJpLAPfBN33aCPUxRw1mQJ71XdO17e8
Mdsipzb06oMzTjlA0HTvjXgXX2a5tCUyT6nRDPDsmNaJYDQUsNjtI2z5lkMnqsPuBEZzHjh+1Ael
vn0MYaa3FTmaGT14FmUAh+iyqmudbgDl2RpRWvFVx1KxVsSleOQK67/YU9F0GLOUzXXdc4ilXm3i
D/4JSnm+jYG/ZetkjAEQkLvbd1rrshvbUSZbeOHL5cwpd3Uf/jOnlOvVR7RrhHpls2+2kNx8pcBe
4QW0AD+/jjB5j0QwtAbmcAUXMr8OeqJ2quiyE5y7e4AiR2wJmvi/NlBjf0fhUT+urduayCYtsB56
jH5UncYnGp2on8d2ERYaIiaYXRzhlYGFmx3iVWqmjlpX70pXZFcm/gYQg074+nKvdNeYaD7Q6oIh
Skq+TXeeYVGOWzvoGxOP7Kckkjuq74WckuclFYfUSBJPAsmwu7fbmzrSXS+lvCKW7KUeEONKOOTC
485PfhohrYo0QUasluJWaUptfMjSN4Y8Vy5rp9yKgAf4r+lWcnfalePbKn36A3GaB/E8h53+SMZ0
AJ0x+soaDZOFmHeXIT8hKTUW0mDYs5krcgd/AFMIwNF3N93td86JzA1vpPdRz4YhnP1iEX+pQEvI
CwKexZfxcLRqbE0OjJ0axloHJQ4KsLxi7MLp2xBKCWn5X3cbphJypdztvH/vOwIzswkMLTuF87iB
BHoNMVzOe9lya7OxfWXN0TqDe+wgi65Jg/7iHuA+WhHRT903werlm60Jd3LR4YYxOegEvj8EKhpW
hiv4mHhUnNLASXZXbm/CphOhWzNkVlGPn9qK5S/lS4fEOz6rFJ/a/foO6eKRD1lynIwjw5VpCqD2
0YAkMMfvxoPGJrHJAm3MgyfwCLEKeqim8QdQUI7IXlqrIYU5GdmEqz3Y0HBEuvhbfZZ3Bfvhq6M1
IRPp8+FpxGnLFVJ7BROTHX/rDhaQxi0mkKfFj/oP1vKHOS/S4+QWPtRjHm3jeqYZu8rWBkSRYvJO
k1jo7a8fM9VMSEs5KM/Mt4DnA0utBTrGBEaUelS+UR3stzfGMqaKzbfRAoN5TUBsFQR1CE/+Uqxg
ZBrQc4XIgp5n4lFG8z+jK1aLBhAxWGd7bZs7C2i8wfg2ur998tZ9Ee0aBPOkSqYEU0YO5byr3rfh
wk65euCfFE6oQ5/lG88Fy6ozWah3U4xwBgm7+LOuEOGoUoqwRCQMeCadHvFkgtxFO684flgEEo4Q
MA+sEyx6zEsyOpJa9GhY0QcpEXxGVTqCTeV8P4TuLGkAq2BGGU/59hg0WraCteK7sVf5kVigGThQ
bGanTtNoLzfcp+fWUsJjR+Eayesi7KSr7dTSK0H0QsMFKPHQKecjYQpLNCrKRZWwAlG8K0IMjEYk
dMVxdzt0Sd95WGRZvxumFtgpSEtjprmxLSLCTEi2tzTgOnmmfN7Cs+QvNqp3iAypU26NUGuCxH2S
FqUOCh3sSESWJzh6o/vW8M/EpXzqAYCik1zCTyPkQIZrnT4cz4tuC6fh6mj0rW6DRq5FsO0xFzAK
knwwFqmMAMveVbsfLb/+pFlyiEw+NxNK27tktnKnQOAO9OeBgqpoKvQmo9VIUTtm9jOvJVrcaotQ
xnGrUnd+b5pS7cRfYhtqcPexKX/OIWhg2GF8ao7UbDNjg3O4SwzgrUbDgPkb1T/ABw4qN0i6YsP4
n26K6gMlAaca6fp64+A9jPb6+HI+zmY+h0HN/jB1do3QssKUbW/H5jPw4NcH49s1yqzulhoIAlNw
xo0dvuK76yrJuSAH6hgMLJuwIr6UB3R8Z1jlURkrgN4Z/asu3aTiFA5yTAF4nQEkxXzbcLrZPZWX
nLRPUXML8lW+0QGLWOYwtWKyfxSxhdKp+DZmASxpPqBDPwnonxbgwbZSWVDwBA8ReAxty0yh0WrB
HMZO+E/1RUfqLo/4fY/6rf972oqgT+S4xD9hSpNGZno342sEj8q3HPoLwk6Y3kUuZKscUlCSBFo2
CkRhNyQnnw0YKxsQTqaDDmpifXDM5FcaA3z0zHm+WtNmzZXnZFDz4/WxOf9UhxQ2+v+ZbLTlgOxM
vP8w/0rszWbiRRuNByv5skcN43/y4MsusUM6x2mv/WONwMN8VSGQkDq8+9p/yZ0xIOT6M4eHvIZ4
HauRHwXGZpLANDjudBaUwLzKn4Bzmlo1iZ7q3658bubVhqNZ/3TYumKohGIDOC9YX2TyEmVkUfJy
C9uJbKbv6QGX2H3wO/2dk9mYwhrh6ahRCFVbHgCY4flg+1tUSjHPRZTUnN3dj5BrWzUkSHxO1M/T
UCO9PiSZPclpU2T1TbcScm4WnVd7z+/Mq64yxcf+fVvE2qzD//fhicia8moXgblabRs2eFFZNUCz
C/rr0c4sTH2Fn7kkQDK5/GOgGW1lduD0bxPe94yB9L63PWV78RwAxNWTv5iwr4HPQlGNtKB9df0+
B7Gz7vJcIKzAClKzkDxcZKZQzkIWs0fSdtwagmL1tMO7prxw2OzRADG2mfYn3c6SlwkRYqYRYzuw
iTtxUvM2Ll36YXAMbZVtkwgcVQQHkpphDlfiehN2u6UEUiw9nWBIOmdYjnp8RLNWcMoy3cn38DRH
rXvfaR/V0skk89IJPeOrXi722Tj+/ffTZvFqKERahieQQArMfFA1BUL7fa7RTD+AWHBg22tkH/9P
l4fmHcM+vjdHxit5UyDDZ+ne86aLR5TQOJ8n7H4RXjAKI7Q2FT3hqh6lwqeHOR5I7jqPKUl+ifxk
PVWxSiLqa7njtDv2TBLptzXMYR1mYq/Oi0B8uNRMO1vl+lrlCAknRpCvQoifxwoNWavF4YY+mZVK
fjJOmsVOEfvcmApAmmd92xBLPf5AHOWe33XSzcsNdj6rifrtP+olFzHuby4tCzd4ichRvhrZSSPT
O6NDS1mKYKllSkDXTqN3eVeQOsAme7xLHBFyUNMfZzNlnhial+i53tkVdF8Vqx5f0vTj1o/mlysY
n3cepQ3AU8VxbRfmN1bgzINN1X4eVRNMgqy8PdGYi7A4nPb8YN/sh15WlJI6mfxrddONs9sOAykm
GcgHZk2Qyh8vHmTxdYF5I9OFsy3z0qHzW8+ybJjDC6DpyxfUJ2ibOO5XmKIe5jcrThKGSPtXLrSM
KBEDk2ahBdxWZBk882VT/mtHf9gG1tCT+qtYOXSZrlMWIrpUf23NmIYmGMGqzWggr0UdTopm1CSM
6AY0yBxyhV6/4MF1EHTHmudiwxOZ5JsHXiAUsddAHfDzrwkYgH/az/dQJSYYZ1JTMZjqsaGMkKsn
d6fWiGUyER2UQq4Fa+EQl/prSEyzc+4DntOd48ZpyeLUrkANIKypkodSCAEa4yF7GbGWFC8tIuK1
TkYCd0Y6noOxCZYGm7ksbHHHtD3eT7HMoS/+B4plvSi2/+0oSL3KLUUqsqJJ97LBV49MLrrQ0mpk
cSYI8JRFhwEjK1o6pfQqOehWlftvkVNnc2EUPpnGWQ5w2LJnUiQ3pScRF3IhTcsM+g9pKy5MqSit
SLn5WcYxpnoqc40cAfoCdYexFtmB8jEH54cry7GU+QRfRn/l1BhRwJjiTcOthjV4L0hLcLIPgbE4
a8le96nlzGHbmfT+lnqY8axfMC/rFX4Rs07xFQ/NLVrJSyeWEthemFhRv0tTcE54uj46ByEsSj4E
gAWMxu3pOJLc7FlxX1WfO7X4SaHT3LriaaXd7y27166WpLo1Wo8X/kNZnsoG+lkBr8bucwWjhgsQ
hfI2EzbMsqPk56gRnSlrUlHLaN6/jJ4uPAKUy8+itLlNw8tB9tvJQjbYWMymR2n9WWZYUHD+2gF6
LTM8sGgBuyiap0xN1BVdpdQWaUYWSh5daUHuZVYrpzuedN+f/xzVKAFzU3t9bYcPuCWE4NpQwJ9X
8RFbUNNLRd/wZyXsQYfl5gW4xSGdzvYZb1E8EbU7xUD3HhaZVAvZpMZJTr2Ng1+8HPy5uAqZ5h/G
iTALZphhMDiZ5A6x4Ie1Jm+RlRCGT+UdpUSpn57M4shlFCq25pZG0p8ZPWxyl2WjhdFPbn+4BtLx
tCRCzHUcaBU54VpAColIJgeYRb822+IZMTjYT6KgiWBoHbHdrPEed9sBefQtDZ5rS9xBJo+kHCcr
MCKCBY65qVuDtG/toAclQZzu0hrp7m0NTgyLpe7UaIGS+0MNMqyrm0SAsr47edhuwG5Gq4LVpHGS
ymLGS8BhR7IE5GeDwuBt5DdN1oEP291NUSJG+KNJwDdeNREenBsSDCVHwPRV6Y+M+hgD2b5+X/SD
cVVHY1FixZE9macDlROKRvsqiEqvfJ5nEr6CfDlnLSTr9ZXI/INzigtyHNUFkVZGVb7xUlLSN1ly
HoFUIT6Xdy8gm5kS/xXVnsE6M/QfujJf85EfSu5/PVg7HG+ARS6mb/Q44FyHrzQtS9Ud8ou09ees
cAZLk8fD6ExOAnJYwjUvAdWMHiCBw3hUgN0wTRrWQFQWypuNWF2heT2SpFIMqpASPnrni5mlNr6c
MMqQRPoQl1o9dehh9uPv5L9WukQYlBMjVpRY5/+aKrP6SWH3qOHxSoTYyEE0VfbxnsBNkkNdV4Oy
zklKev7LxdfJyUhvBawF0AjDRW19t38TfsMrPwZvzUGST2MqFgchGOVrP/+YW5z6+MmPUfeS63g7
CjB77Q3xmyCjqkRfw4q4P5VfrkXebprv/zg9KvBU2nve4KK2GXfTpjyx1elAsKufOsFYWPQ6v559
4cLW1fJ8QWatr2P/olPdl0X01ppdDbaT19LUH+woVjYGBfj+lOXXJ2LL7F8NEAwgz+R19XKbt9ss
QsqPUVjUn2uaWA4UqVnQKlU7tlqqzgSV/qTkfnDIgmDniIaali2jx8oqykXRc1QV15VgdbLDVRTg
7MKFAM2CL6eF7F+E4Bj6NKd/GwBpGFOsgA7fLl59FCLT+s957jYbvx9OGaf+sq6rIjpmFD2VIWJe
3m/7VQWlgfkRRtAjVHuJB13bRUzGd1JNrzkBrrCrzo8jAnufP1u2O2LJVZY11Wm29XKYhlB8ss80
H4jviq75EiG6ohBILXOyWfOm6qO4YhSRIaNN4WrT5B+uuwgnqp2j5NARZwYES3y9ii/bVaQYBr+8
qMrh7LHBClXXJhUDpORT9mTPggfIJJa388NnlG4I19F0ou/ykhrPLcC0KSuu90B3+ddp/hV7tY2n
dHZ877rYSKGbfiz572jY3BWAqg21NNASxG/k/3iiTC96/3iueebwKTRglmjaJleZSvZVH26JPU9x
Xxow8Vzr92RYDIjM1Cxxf0FUE8kD4/fPBUQhUZi7CUe7ylCPEipuueXcYUFvp6vOdlX19RGJxcnK
AJ3xPpnWW7BVWOmFiR9sNU46J70oSNksslVKKzLz8bmRakCWIPVJZAEHJULXxgqyElbD1PjKzEpF
INFPs/nWPckn1Rx6HKrct+jso2a5U7oin0bb2H2yPBj3xJ+eoIvoArOfiHHfCuW6+SS0QC2r7fuF
a7vClTZvnMuHs1sQeWrKfufiLdMcwz8wkHH8C+hr4/Eze9KdY9h3osdCIJRt2JN6AXRpo9NuAZ5+
hML4K5Dra3PkTHuLvYtqGY/88Ex60UPdn/dhFe11Wt9fd03vU0M3n+e93qQyUnbxJ7yKHP52bT1m
bneKA15WG7H9NcShxpkwI1xmFsvo31KAOSJri6u2PkTyP9B9pdius3ekeMp7YcuwrNtqjzoboNX4
NNihHvcW0eLrj16YwPZCn/f3CqaSYPAK2TB5iqfSqesKtHWc9iED5vaByIVPhbk+Yjjc/+ufq/BH
ZDBqZ0y6OeG9gKrYjGQX/RL4NBLvroN6F8vYkeVEqrxRftotvpQ67DmP8SSd+Lj6SduFoXbX7y0V
rm6unBvFqKSwSlVoZHnjJJvZkJspg7VONaaSHTlztOImhdUB4O7mAv60gltL611mZ3KXqPZOS3+O
8/eNjoXmIyWyaYxoI0kC/CKad1WFC1p/HT4awSIwOY+P9BM/H0uFaA62xT1lrBNBz+ZjPazvKqGC
KB3AOvAaGypzgf7/tKH6cPUiSkEO+4ZiF+HHu0N+/5S/UC/ViaVvqEk8wL49a+b33a4kih+5x+nl
kYUcLw+HCM7nP4RJiv74UwazJvtTUdyKzMyflLZkcteGO/OmKMNvXPjJk9nW/Z8t5FES493DkRgO
9AFu7gXPaAkoJrcqvBxLQ28fCcPhE3EsneHNDKJXgbqho/s1Fz7RuRNDi4OJRvY9ZjmXOW9KRLwo
q5Uck1ASjgvx/gb5U02Xn9h6usyJSArYG57udkoQuaWrhIFGqSKSN+zcx7OrX6F+WvdO6ooKGagE
thv8DIMuTMKdMLnnEQL+JI3YqlLfEujb1ikUXBNh7mL9MGFM56KZshS8KFDEuIGP+nTYZrra5wP0
5XRgQyD2IgOMeavOvjsDRHV0pNf/YD5Qvu1FAp/MFCvXW5N5khCvQBzWAT+OKc0QqStpTK6m6GqF
7Qz9ANk6PlLg0FNRERTPZyooRDLZ5q59LaJqnJmcpL3N1qHjdRrq9PK5ra8U0c2juR7Fjf7KgSV5
fYzr/md20r/U8GytI7C6DBn88Z5GDLWtQ1ucNsHP3ToSXc9vI0BV+GaRX9CII7TAGkIBpt5KL8Bg
hzGliOvzRs0itUmw0McbjMGP3AV1gP3+TAI4dKRfualkmFauSWuz7ijs8upYG82tHpFkz4Uf9E2w
enVL01bcuwkQuy/uWtltotn8tI29IAxw/xebkUbH6ZkQjYRTbgqoIDvCWHHjIQ8HtLIDeoB5yTSD
mjYJQq6Ieg7CRcnHZaaDjXrG+Vgw4rHazDCfaE/nx/GW8YaV+I+u/enwxT6zV8tdSyDzZ5dDsy9c
bKc5SFRGeoqHPCoX11BDnsNg5aBBdDuLp8Wi6PXvm92phEXvwaXnaZY/yIUfxAFOBXd47i9bu4os
mU4Hy6Jg382IYbDalmPvZ4v6ZuxfCB4lSsX83dtJ51QkoaJfPu/B/p0qoguqdRovb1eG7b7Kb6Pl
Ocac/qXlfPWG+IYE65nfVn6tQ1/DtTY+idBALu7u4yaAH1Ln5B3HyRsW5TIp8T3IJrIL6HAYEb80
32c6ef3Tyr3+/67dDC9qENr2Kz/uGDZS6kPSs7QPkwRZzE25jVvuxm1AA7AUTEPJ2yYL1RRGUgCB
OZFEVAmM49ENUL5mokXDRZeVHct1ASXkhFrlxbL9wnpX3cJm+ZOMHZwAZGYFu+5ZeR7K6fOqFVs8
/B//iMaDDFHXRZJowjgjyrbEEdN4kxCbnWNNpLAvD2rGf5ICF6VMgDBY+2lTfScQExIFRR3Uyrdp
WpwwqlPnWPfTPFtanWcac7evZYbcVbw1XZ6sfkwxAvClWlDaR4mN7L8nCKqL6eIuhOI1lfGRaXEp
0fwSlr5GNDBaMt7OKZ31Xcd0AS9G1mp2YnILFLV5JDi/eU6lFdfpn8RYaYb46qrPnyZ0kAX9+4TH
/MVdyDy0Egpzd5fzQEYRLKEElsgRmyMxwBwOar06qRDnTMbTnwXv/ZshSOcREw47dSuEDNHz3e3h
leqOR3SQBwEfsiFcnKG9LUAgm0Dyl41FnYsYUUanZ+nLd952YmeV/ovAO3oFYATQxswSob64Zl+5
qcHZO/gDbd9+K7p0cA2ppsQPSQwKsuYp+uOki1wtHsDtTy8Feq+Yg4R0HKekNjmULSqImC5idzJN
W1xN+KGfD2qgyCI3iVefd0A1U4LJrn3SdbttiUqLsJ+XBPvPujBXFGuWMlkelEjOVFmmcEgyOr23
IDEEEJjQM0cnZ6WDCVDjN0ouB05GBq4iMMYFe3e2GzkL/hH53p1eSDBCOyp7JE/qndsGrKRnSYcX
leDODwiXFC8cpdZZWbx1koeZ39vgt54rVS2D72oBwSOWjwUAcML4IyI3wTYkxXC7sKQi3G1pZxjw
OptY8kNCFXp3ObK81d7MEDxCx7EgHyBEXHkou6/himXiGU/rIwPEhyRMQlmjswqTrlQIUGWByj/S
c3IgUgwfQRnJPjQJbT2FBqnLb4Sj15cM982/XNihnKbO4Uh2jc4ZdThElr73qNqB3K12jO9ASLZD
E5N/kfOWPVf5XtZ+27d58WdDNYoD2BJRvjnKUjYENIZl293mVOC5AS46qQ71gztm1TT8BBuoxJr/
icHIHKmyG5yozyo4PW8gy66kBgnxp5LGVgc41mnvbzsss25YYUD5HiaX5difXuLdBzaSnTeJxSdk
4KHRVJfKTM45hg90QiK3aheWdN+u+SeQbrzD3IdzKh2APdMrbdNA6KBL4NB6qxvTtkHa+cxUhqK8
v/dxp2bJJMVhV08Zu3X2kYNodw7BWlkwykMTXJJbBBMIlED5LJOe12+lM70YvJoAmIOrZg9MgQ2L
rn1as6IC44brdJDrsblB6wwmEdlapd/7rEGr8laefFU/1nsufuNM4C7XT/kJ2pmNssqHIo43MN4q
0O5znmhoPpWwIEHVEsIy4MI5my/qulDA1Cp5/wFbo53y/aO/ah77dAeuF+Upo8TJs548zEG7FIx7
m2kb/inbSiOovE2Jsk1fiPB9NhZz20a7+Z57eYYCjxS5QREiJuaGWPjFQuL29J1RvfNFs3M+nGrd
A+M40blI+vtjMkw6RKvuvOMoHcG4fhONFDa/Eg5h87UbJG1WXpK0Q3BE88wCqhqwG4jtNMp+IOeN
MuV4V30N9qVt7MxE+CsX0kNac1FyZZksGy7JqhJh+5YebAFkGuyudfESGq+vDn/z0VABklVXRXsD
vhU68A5X5heNw3mpeoSQDL9sG8QxQneQ67d6riFM4r+CQUnLuaa7dkv5Fz7SWq4QpWf/ZOZmn+U7
sQ0Cdi6PZmDK8PZNakSkOmua73IeZ6KFI6R1aQkCjs/ge3UY9PB5X5d8demuWZ94ZxRJo10azKWW
PAL8Mx3nt+iNDofk8Nx8ibDJxBZTYBLOnFjGDzQNoyqeWmKhnwA8mYODeQUjg7LqQHVm2SGgm7XN
KjkvSHb2n/eei6o4zWfqeG5FcHjAe4SsBnkiraMJazVfjLgX60HOMBLSNbGs7/vPQnK+jvt8u60Z
zXSqaL84OtV7UKVdVtL9BtZk5LSbHGeEzZccI4nw4S2SUc3B6V8e4tdQNqXr2u2A8/wYgpq9ZfKh
JaQModrreiG/R1UeNIf5unOgXI3Nr9GoyEq0qUuMDKnBN6HUrIJCwkMQQIhA0x70497JxpRTfiMA
ZAPGuPiZyD8cu5rlPN+iqApHjmE4a5+ohbpIZ3dObT/01srCN2lox1DYKZQG6KA6KTiu1jhM0WXs
kDfh5vPPHElcPNhvLjN36U1RT9IibMl1dV3Cj0odynZLDGKE3nZ/Q5RXC7FXHhgvpqTAdezlpas7
xlniGoWrDhD4C5lIClAQcQoX2qk8UNxGFaCdIFdIZ4r2iQf3Nwf/xuFxq4yNEZPtcjnyBmy+hsX3
fpnL8UYBj9nTG57PFEiRYAk4gnBx9qEA15AgtfEM19IEJlyEkhAz9BonjEGhlZQO8w8sI7VIGKoh
kRQ8q7/dCVCOIo/h9y+Kw79v3Ajbrm8hYiK1dm+P04+b9LIg6q2rEpO+ql9xdSxUxtemPXzvJdoa
DhGtsoaul1ZswufKK05ZImIxFLV9/nkBbaUjCul/r+T7Wti58uWTvL+ttOaBnTq06Zy1s1/xHyWm
/ZsKCNmvj2TrPZ47wKcNmUEyjb/JMB9vqxdXhGfrhO7kjhJxSaIMJCS2GMr928mX5LS9eUEAU0Zl
EXTontz1UwVrnVvOcaFLMXvE1tg40t9DXDBd61Cb7XDgWoOLo2wpNyZ/9MbDSC1MQrzczP+Oeeis
Bliji1xrVC32jKJfKWg049+ApeJApOxhEfICraEje17I0qHf5znuxRbn7Dm9M7nKciNH1WgSUlOs
SkT5Cobv6O6dF8wzDfjY2zA5C5MylSnFjKTHkiBBC5tPr6b2IWVpsC2oKs+mD0HeBr+Wk3ffBEbX
6TkGOJwXvg1IoDmYFX3/tkW7ARPP47a6U4N4uBob56LJ5NKUsL/+T4FAh8cD34EreqlvU6TG78AR
KdC5uvoNjxeMh0Iv9nsdExBtXTcGhzJpcN3plr4iQZwBqBuKjBeHhjy67yvVtHxJpyAOIR3I9KAb
xC9aCqSJ7HxIS7U+VRHy/Agp7xI3hmz4q3/vd+XIr3eDwAWPgmZKfP4JFn8ZwtzNeDQaC6k+ABaL
phTrgD41EwhyAqA8ieQwMCCKd4ABmXRFpg6aav1chrKcpwMIzWWB4Dom/vSFD+8WOGWJqMk8lQxP
yf6Dyd164HbtPFshU8VfYHMVbsEEEKtN6xIwHWje8e9MsVru5sP76MFG0i9poOa71zfVhMfHgLmH
NsOsrCv7yRw6q/ZeKmlTfsI4yofllj4wKKEk+ZAvBxkYbQ4YZKe3ZNaFfyZrAmXWhEsXc1Crn7JF
x7FyxSpiXtILGOzH/sAYrsvO8p0lyG/oWTLpHG7aHz+GarHOWT/cqvSK0o0C4MiA5CXe37tzJyuD
F+NhF28pIYq7uz8oEpJL4KshDIu+65AJSMc5gfJYieP8PBQjBzMFPfEbKwg7Mkv8SteS1wS9wnOM
VOy09I5zhWEmTkDiZZGMLAxaWUUSkk6AOudNuJaQ6ADBLj0Nv2nMUAghF32ZrYjJx7X8DvpyLExM
NyUdZdFN/sIS+nYsWL4BrmYT+Ykh8Pg+/dVqIO+ebyQpYqkJXDx1W/KvByksfDgLOOG7cbY+z8HT
ZZZxBzAdLt8XjIzV2bHeQUxTyEY9EFUNE61Bd6M2W8IedPVS+/b4ByazgjGiCP5gSWoB/e5YGqgX
QcWVgDne+pTfbWl8YBFrQPUfSwxfQ4gNRLNh9RsxxpbTwgw2pmGzbLLMGVqO3Xu5lZHrypVf1tgc
/PoJBjNEy3AL8mAF8n/cEZIukHjtICvKgGhWNZxLoQ107XqgUCxRL6b4cMC1Rn8Du0LvQmKdF9cm
UteKwOGZkumYo/OuhNX0O5yY266ivC74Jjgl2C/FSN6Z5JjdDK2ly7YwGHQaSou2d69jwR+CuVcG
HFpT+b48DOZdYDqA9pGARss+xskjRWr0U/wF8TZA8N9ekpudGz0qDIPm3BIHCDVi37lhniXORU+P
VPSup8J8DNLbqHG7US+ym+E3DmMVwsI+x/y/d/8yY43mAPeV1hAMddQAE0UMDf5d8Dqn55vTAHQ5
ykKgaOjeLeqq/eeY4uTa03hnsSHcNN+OJxxAVz7qlJhHkO6fUlTHk2riPr2UUlBtsjK+roj5NHOh
HUXSh4hgzBENRtwInfF1hwn2d9SULjQApqX9y61BNHvWT3OuGPkMZOd/BYAQ4dKEU7SogknfgvBB
O3tjMX1v7s/hS/gRbsyvbnXG3VjN+vkF8GadUHC5gUiOM+JLbiHy889ij1aEHgTyYmwaMPHIf/5N
+2tKEY+Wanmq5GJmeMPR9YPsv/DOGAmOI3ALr3NBct4ME7hwfw6W2MIrqWP39sIVQJ6py9EyZ2NM
yGsugBmXoy/Ilq43DMk/jJUKH8I9v2IxloKhS13a5VjNPjLyPuqrSDT5MJDwtz2PunfuV8Npuo6C
EA06CLh8VxSynFqpQQ/qNCIwUfsk39cqIIqNuuLrqoG0zfSE/J6JwJjHMdpH/MyEkkMDtnEYTXvn
Ah+lYFtz3tND/xWG008II+Kj5/9XJZaUdbzGV0UpM2ESlUbR4B35b0G+0ToZIq1lgVY4asCkgXwW
SbdBfF2FO6yGzKMzHhvOp4pBGZZ8zfKP75NUUxzwPkyit+g+2LJSzR1iqVqbk/2Ndc07buc63BoF
sMc+PIAJDV5kFQCDBaocwo2AQslZu6xA6z6u655b8wJiiLCD/d7Iji2zsuiXma8iYjYjJOw+59hB
peyY0Ikn8pmPhEFVLPoN/pr7FIgxyAnqkBGwAE/yZpa0E1yuvrV8ejMpRpfYNaYIDvIKLvrYMdUQ
LNK4x+ZMjYfExF1aZJ8fxwPd3HiUt96gcAbyjoxqcts22qtjbpTKrMy7UJwXR2Z2oj3qX0wD/Wnx
MCZ+Ix67Q+IJC5h+qnJ+e+Rp3YP327PPmGe3EJA5Fzr0nmUJlAUiBTOPCRf9stvpwrZqxZE3Qgaq
jzPNe3sNMAmd5d/tv8q5yvlJhI5LHOLLYPdIfxmQOeD8jPOn6ms7UOKG1cxGe4j35Y7b8ekaGbuA
I0Y6CJzitfy6n+yGBeyIsfv9ovlk8JgQoYl3SuZw/3uMIWTFWPyXP5gCTECL9AzECbOrhEzODjPx
Wu+0xnwNCQrfiIKkKTyCu/KzhsZrwsNPoM8MU8ltW2sPwLp4WYOiYS0/KGebVQ64q4P116Wh8J7p
njIWEY8MtoN8N3UqEt1zAIh8Z9VYD/3m6ilIdklRj0RCpldeCgsWLqpAXbNHeFt+EXRTDHhqoOZP
To8avHLOgULm4haYYgZOK0lNXErwV4E1EOAqD5t4h7bvOhXwCXF5UPtmABP5QW8KadI6yOmIp0SY
cVrYG3iDpVkfa2u/abYVbcW55R7u2TKLyu45WgL8p56hmoEGsGAz8qGnn/LstkOKRiiqh1PuOnxZ
WUN3kEy7BHHXDzNJM3PKrmNNVD5LiDag0eh3QfOIGvKSN0LBRZmnshoqalBH+OQoCk5hz9VtK5an
LoUBGeWL8dus4ndEEIgt0oMQFosXr7Yzz/rlo+xoV911uTPgvPFnjQ+HNJMYC6hdv/SAqrxAuOFD
9N7rJP4/tmBysOJ0la8Lvcdq5GTrZcLtXhd2E6B1+GtrLLbjA2yuU4fz/0QIXIuGe5Fqzd+sPnHw
dvMUXsnBAjfCrYpg/WCNM/SW6aU5NFjpcA0HX5YJDiaq5u9IVuOaUdlv1I4FkQHyJOkwXVz4+zGm
H9QRdVLfZUzgpetSPYp1qQgex9hsK67v6EZsO8KHOOu8RuYD2hJ8uvbKT36pG7/4KIv1T7ecgm92
J9AALTVgfc4JAzbw9tMpH465CKadCtD3QSdEsn2WH2+45YtF3obleslD2K6BL4Nub61XnrjWbUYh
OzGi//50aPoHEe7+oeCGVNxiRzd7mb50u1Nq7QcxJxMmHCBBUu3IVW8KqDjwphsuH6kLXLojIKaQ
Ih5LHbzP2Bl0Ec302zM3/0BBeK/0YR81THM5UXbi6OqPAp5CdOG3BbijJUsk1EvlXAtkxMzOFkz/
T/6R1tANOsKjruycxvLP/kxaBkOVCo0ClHWa4Na/gJrxLwByI3C8cPPK7qL0Owpq0ppgfirtvK/t
Rf9RVL4cCuHzSaReayIct8OppxHu9WyTvZH7xID8+QGkODRYU8AvXRDSddtJOznmmPt5vWnS9VZf
KsL5SJZQ+G8Nxn554lHadWd3A5Gh+9tKB5ZkrSypH0egize3ui/7eT9SXA+vKgAh/90Seggb+PBb
QrSNc4rwQF4Gg2pNSL01qwBJPPgfaQVFfDW740lG9Oxbc6Q03HACh5JmL0MX+J72zKJjI8u/4ZPn
py/7tZzbhhVTybMagcVUw81dl/oOrxG6GS3cHyiGAa9/4hD+GTCp3DhBofqeb0RVgXCpGoe+IXbK
evCHOr6b3HPtKm86jJeFutEH3oNf1sTAh+ppaOrusToL1z2+wrDGYK4/6VL+68CqSqycsAkXGGgP
jqJreWVRL5oqNFfQi8cOy+ZqY4P1Ft/mqwhY+qyPGVEfIwJmOYzB02Lh4tnyP1BnyBExBRz/Owzh
OPEGbQ8MsMut2RvbPT6IYBkmoclvcm67WNvwzSIxh7v8rfFbxNOI+BfEpy69056dG4klTHnb8JZ3
SskIJcCwA4Qk2otQq9skBDR0Mi3oN3V6O/kg39r2MDKd9nketqblI3onuKfy9boChYTIJFmNBLBL
BgPROuVqqyW6Wj5jZupsKpYMgibZ4jNMtQ1V9nIPuwGduuk7Rj4rrTKjv5pNWQedqpZZ6nttMdZP
kngF37xgsvzk/bWkBwcLkoTVtWy/V8Vm+G16HYiW3zS8Q02Vj/oZV1dQWLTSdc0wqNGPh8K2EHs/
A9ccyPXjnnAU57EmtG3Htfdq0PSy5bWCSfVlPhKsCYV6x1EaHYqk/zodoOJTBvLetRUjuC5iC8Gz
hahxMpUFXLkOpeUjnBw0p3j3+TYTM7NIAWFtT0Wdx1M48b/ER8FvIHKU/oP2jl+javpUjoQOY4MT
3qqN4q1QZ1ewZ9X4C9FNPj3/uZMTvQHQ/kmElNnX3+gkc6DbDT3CqSX/4Xk5WhxpI+xPRJAqUD4P
rIh2WqqlX9sd6giSYkLJxdXppbo3HRLgLB7IRDNFl2H6Gn4UYhqfqyvYPyK1SFHVhegoWIhA9Esy
wNC9w2es0LTKBx67dVgHJpfqJWTNQjiIa662Fwa/sXWQVOzblOQVxmplHH+MM2JIqCRaEaou2gH2
xK8XvmteI/SvnN5zg4E2xb34FCsNWuJDFVHd0SOck8vdxUBwZ/KGSOwMfXPXKDOfIXX0mek6yxWk
JjKn8/KCr0R3+EU2O8QM3A/oievv6TzKZfuukecqJ3F1QOIodBqMYsojN2DZBFNd+HoTwhEj02Ni
Cop/lu40EtlZG7abfUkRnYzxBGpC8dNsQfP1CuFnsniYJRSfyEbGED9IF7QjPnCveJn/x2BRQO51
CWEtg8kshKtfSWfLyoKN+ZxzXWazvxHmvdEUECzbuV7Wn1ZsKj2qPkeSIeipKX0MkiQMVuCJmiFS
OINwZZUX1N3FVsCIX0YfMzlk5paiHzuNX+stVXIRLTd14Ss9YcOaTZcuhdHleKz7WNlbba9E5UtP
CAlnHjqZ+PcvgG7uJkG8hbEIXOQefmpufF7+z7c8A9mD+axA6mwEv8BVEyI37uAygvRkYKF8aKAF
BR9jZqAB0bRuP6WD5Fi0/6MtR6/2Rv8flkiQwYf0bEBxMWuatXZJRBvVLdJw4Pid93VEVMPHfgyf
Iv5bi6fuKyzP2cMruVPlJXITtczg2VcJqiUQ3DIWM1GgQLr5pwDqLlfQY6wPEPtytg7Q8eXEWfpc
EvqSJGlwu+9Oiw1qSBpz2xKxUoORdwTiGbsB0HeF1rDzwE74toRs+WdDc1RwC8RNewipVcSHdbhL
UMYRM54QC4AARPDQKYg65vRpyPbbccvnZBdv87ZYdv/tvKH+DO3ckDr0XPe9Q4X2+g9NUZA65vZH
qVHdlD9ZzCxrqFbiLO3bhIY+Mzuj9MpU/uYwvLQmsfVNz9BiIT/J3EBbR6FpZ/eJerUEUIMQGg2s
/zvi4/gTIgVkcPLIGYsKcf28zw3IQCBaVP468ByTDhK1EZhqu2MVH5C+JXKQNhuwgAZt+nfQ7lVI
qoQv4VYkhPoZOFf6iJJiq5s9e0SIo8IvfFvJdM9pdRAL/imO3042VPa2f2dGKg3uQDwHjr0ZztHa
hxLoSdPBBQmB94BGdBdjBVxQ0Nq/UGsP7TU62YBuPFaQ+IzdvHb6MzGrwBiXNPjVAjgN2RGoxJKS
tYfjM3LCeDSyNRZyauLFVLF9qgiCvExjRUo/3gPE9La3KyvlEUkEBzvA2KHePtIlOypdtLPtCmBb
qHmfnSA7pXJJOJxKypWFSxB8ui5oQv774wgo1moHYtbZt3o57dUZtXXkg8gXKdWZY5d75OWs60BC
5+K6vHD59qsdkgeiShYmvFe4MXT0L221hC/y7bjahQffgjuMmMA1z+ielmMFJZSneyGONlSqUQnD
oDWF3B8QyebfLNCq6Eq9GwQDgBtCeeyLBHhXmJ/0y0LaRyFnn4jnNtwa1lA1m9HwfupK22JqlWem
YRzSN1M3R/gneDNwxt1dkItD7skV/CVoE+LjnBCX+Z/V0Odhbyx9mMWlgk6RUgCSuZFkbT1qzJrw
r1jVX3i5U04itrV1sgiHNt6Of+Ge7XGqGtLifQbYKOX4UGcPYORczdziMDY0JVynnhBbZieq3FYq
OMBOsGkIwiP3Orj7EyU3u6KcLe0Dna05DHreHMxqOaJGdC3XXB42sVxCRncsDXAZaz+GAc1yS7n6
M8aOU/vMqiVIG0OpJATE0FsYrrx1CWSEk1IRx6GVQczeRJjDSGvkBDDepJdNz74JtWLhfZOz+Rld
8ROWcGTnnbBgYNO+DGuilAKi51CS6OptrvQ3MLVgXUP6/RzLMkGrdwKqLDuyx75wzMaTOs0iTSrv
JbdnJOy7YoZuxmjsCYHkiwE3kzUi37cM7L0BleeSI2muMWQvnyleDLufmDftnd2epYxmLMFYmPvE
C9YMw14FsQg5BRuMPEZnriDlGA1FnAZYh63pkqGYemJmng2SUSaAbI7cVRwvAZpYUROnPW4dWMGi
M9hVAphiEDt1/BluSdr1UAu9+O5ZXfaBytFVvQN1WKknA3zEh6V6iDElBvOEK5N8sXuqxFqPYG+8
Vu1I9uigTBkjZ168z7YPzNFciPksmrjtAiPDCr3G+Y0QyOxNaarESwz+6188h6PCWgLFn5B3Nn5p
3na0C+IQs5MQpfCU/nmflz5+FdrVrKW6TTTr5PZ4h6+3nlbrdVW7vQlWMn4XW0AhTx+rK384/dVs
VycZspzr3CPQutYLCsK3Ie00sn98AaIqK0WU2PN7To4cJtqkiyVQTZWLx4ATwWYvQT3iCsEj9gqY
oyZxnE2lAJL9uH00tIdOYLhkpJL7rHAh8I1ARqrlgP+DbA6a7CxBxjLKsibtfQeaHFuhcivPRMj4
ndWZq23oUCKS+2SzIQUUErIU/qAz64dg/afuZ5e2Nx0HvkkKaPPJ+iE/MKkWR9dgMZHjPTXAdOCF
JDW6AdawlKORI5TZPWrQPm4dPexR3qzW3axbSP5jCLaNl+fhzfR0tJW09u9JH4HZsNqilGxy+BvD
rbImg5RT2jzowFAiYUVaJOdHCEiWIRqNhvpayJuBFcldhUr4OM+CvefMPUHihF+r1dKxh6Ptxu7N
H7D61ThFSeyIqAWtGtkm4G0aeKeyOw0piUv3F75t9wAg1eLI4hqutQ3nnbsOkpGt5tGwCn10ANDE
n8O7WITgQow+90MkHyJYV+EA0YZvptxQXho7g3YXgTXeyF512ML/nRUZQyBA2+Ww+wKbCbgILLQ5
z7HJQ3T/Tf6Ber/WfMJHsSq5fs+wR07w4r1/gSfbiYcAUTVqH38mTFxec7a26Ghm+T07zVRpH24m
IS+JWRPuXvcMOSQHCxh74Q1ElAn6INvlOJ9fku/x4oL/Yk6IqtKlt2Rpz6duDJWg+wsIbpv+tqmX
/QmWMKmQobXpJHpNjhiz4Ufwejoi0Pgwxd+hJtUEUVErJAnMPk36aon9Qdb1bmFYsGUEYeVfcENn
Tk5Ts6oiryMgN0rWnoIAGvswXVJkXxwz/fSCPtacndC7PV8W8rhAFrONm9M9kG1aVNTHyytEfFWk
y2AHcD8ySwQnHUtu7EVfZfSOGuGCQ5yT1of/uyg96P3qkzS2qSTpCNDrI8tXtTw+OmyiWm/ey822
BQoODBqsRFYo7PAdxp79ZmkVCY6sW0sF0EhLU2DrCRGAyxlX2fNPmcvYgri9V4/XG/nNN9GBtE/w
SgOo+FMi6ywrgWedUH27BYn21uExmzPajlvd+MBTade7f2hhxLURMMDqqiuCNgHwHMlMIN2D5yDA
rrK3reKrE4CCuChJ+f4m7GwtTWYCvyyWhZ4QeTtLW5ROjkxnoLe0nbwz8z/DIq6gtVfVAFCJjhfd
1Kw+2+y1hinq527GPMb+Ft/EzyU7nDXRRJD6imdnK1rU8mnBWt99Uaa7dh7Y7NENLTEqPyeuQZUn
HtcisoycnhbvfHm65PluRB325rtZMZL48bh6o1ZsBzkHm2BM2YcFihqgvzQamuIILtsiZbDrttlD
filNzZ/5jd+aoBjMSLe1ZgE3f8cPIIpgNSnx1EoqDlKsHj0QqCn7JKJfnQ1+58OIP1lumbXkLzji
gzYbkc0rGxyscUlgUidQGajnxZrMGHUVZNeUi53Iwp1OonsAwh92dkoaCaqhlqc9aOFEoR4jBhU5
A4pSpBDy+RRIuI9qN2K5qGo+A6rbBxAlfND+mgN0KsLvPOIKrF4gDgBailU+up2adG5ibGCQOzU1
SYkKbhAMQBj4dP4ZteoFXh1Sr9uemrXL2HrlpB67lkrU6PgO2nJEMQuy9OJrmQGG6fIuffaTpq2V
MKC/tvYymP70H6xqKd8692iXlaRn/e/tfydUEuF3/HUPAu4CG0p+Yhp0yJXKF1qqnMWBwWuSW3Fo
MaBDBcYFHDlI/D0rQGCq/5IiSD08r7dolmMqO4O1/WHrrmyKsBeUo2kdxZCCR5Eq0wgjotK5ZHF0
NI722gyLUAg36mj4qeNI7nDznd+jkn7LJEnLC/xqgN6M97ro9z6x8akkVNeNsMK652d/rwJ0o0EU
Bq2wS/bnLWPAvpqM5af664U9Tc31CwdY9/ziM/GlOZnrgN4D1mQGRG+2y7i8b9bn2LYgz3r88ijE
8P1fq2nqd/eFxzibS1wiD8HEXqC/SB8oYMrIhE9N+stbO4FqcpeDUabbLCAaz69bh2G2ocssxHbA
airHUKRKpR3uofuh0KMd3GlIiPIuzfSCxkLMNumAPa6AdiXwVB7OkjwDeGvLz5ytoM1bEdsoKBdC
WgHXX0PGhMpMPMuoI4mN8iLniiprNrBEwWFrJGth0NB6GC6rAx5nQCbNjAusdqGpfFC0f+gs+REX
zLOT4otIvgEirqxd9P+BCU4zclb7yGXn7WzSgMOOfqexuAWj2wrCkyKWFq39a4CrsKPriS4jHJz1
/jgeYz/7d3YBvwRWpbzsDAxXh6ESp5C8W24QvaE+Z67jZgxBVzzXgKFDtZ69o2B6K++PBNAWp4Zw
vDjPyUiwukPlDI737KWXJFcILTssyE8faP5F8T+72ujJrfS7o/N84IgNucfoRQ22Dw78XBnsIur/
fzfERzyul+RmECcvSiPy5gwR0IjpGaYPW8K+740zGX4yBhOckstIQjdJle/JYvdu6h5h7x4ki1ZU
DxiDzTKjKBOAd9ztVWqLAeWis3S2GMeC7mGcjWTc6qyI9HpMHK3Aak445tN/P/dU9Q1g+dJ7chfA
pGeazX2qn/APye2+g2CTEBjT1hvloaBtCT46TResTKglpPFkE4VMAfO1CGNDyEBN7CHUQlSHIqcn
hoFnUPicIbJfzXYNdH794LRQpzgLIwEFEC79XaiKlp3HSDRYTciEkxxcXUkTpyMKPMpB8RD5CA8t
sRGlkIhuyJwrlSL4m9GVazCmhHRWgwz079OwungtpxCZz8YQgZlizkMFmFQ678ntAsbQKBp22qqg
Q0CE8wpeaXjjV2uvmUZJhP/AcivgOXhsf8WFJwLZv36I4s5v0cy3GP7azxLSkL/XM4kddOfsj2Ss
357tT4ansopjh8cs4Yz0rvMWekMlAx/4dp3hsKo50feIPtRjuEtru+jUKOboxLKz6TJOrcRVmGHx
kSeO0K3TXJ9IUWlJ0uTNTU2JsIy5EfITy2qJE8w5f/IZEhC0mkdhXDYRzJAEnc2E5mjScEmw6DjL
0eaGEzJk44H1OU3wLbrLcENqbE98z5bn1x+QPnRndwqAgw44Jdk/bm28XltD9rYWh+0THQYYXOzm
m3sQxL3ntclRq5H9L7MP7tQDr3pCGKIJobJw7NquKlDqhOoh94hSFvJxJJGFuLoZp0R9mcy1jq5N
3SfarFZjITz+9uWYMGf2nKBzjK6pBkc7odocBZZf/TyWB+7Nr6vsHjqxC4lIEU0Y+PC2sM04OK82
fjj9rWI1hHdGlXBTu/wFMyhzcDQ+DPLrc5bnLlRBzradVTLJx+IKcmlAq1NSorNhlSTzpxpousbf
+QLoRQ1IdWDJYt2MGMSXjZIBnrLtL48C3YzKUTKapGSMBV2M+JsBQJ4S7LJJ261MAYjkKLDtUNdk
psjG6Y2PmW3yfjK8xXm+5D9cz0qdEaVelARuZWzSB8WVzTdTBuL0bZNnQVP0GRBluV73uUOkySLE
zy5u05pq/eGqY/VbJD4uTuL5jiideYlF6vzuMq3pYmY2tAzo1zoPaGyCxulMYc0ROuPd0dDGlS7B
rTOs4jgzAa/2uzJABb1PkPTb+ttaLCOe3hWGpEoyCu+dA37zyh+f6dp5xZz8mDHTCeHYLwgDiaVB
ZrK6Lp575cxaCbGA1x2X4YW6tvYqWj+9wqMssD41MNnW7iOKOGtmunK+SROAFFzhYHVl0dB/GsKQ
h9HJPShlKS+KhswLGNDUPdVNuiPXQYHvcIhcuKbbDe9Nmp4n2hdFfG1g4F2OUzC3mIHUHHqHqkKz
Q2C23OetVih4Nep6jrVJalqUh6Sm6LbrMOKXhFm9Sc+3WVxHPxcmvVyfsgkslqCnk5r+3wjdDaGQ
RApYD6ynQA5SjRvbGIEgWGG6PCd/CQkgV0y8S/euwxVSmWqZj/vxmCSV4yQwSNXZ6qJyAHghHsHc
dW9DwGFOLzOBI/VD197UTGesqdiTKBG3Fwg1IZpt5CpPEshHImNMqNR9sowlEbrtHqd4ZLU/eWrF
nuzzwMov3dA/zhnDEjTvG42TSc0k/EBoHU+GW0OABzqFr+bBEaM0JvhmWEVH6opBwqE/6AVPA230
hMxUwTPf2+8GxsYc7kOYNNYeYHElR0Pb62fWidff1jsG+ZJYXhTdoG9yu8I6YkEC3cD0zXv00F3U
kJsyOywApFzfHD0T5rRRLgTjNt+PW9/UZkJ/ORnCcgJB1ukUGYPBoUFMw9fFwChMnGB93hWiv292
midbSt2phxUL9GEP481i9la22kMnHrflVaUn4OUA7fSp9Gs43QzFQqFKF5vyGU8glESiKLQhfNw6
Lvbx8hbrvUONzQ8Kv5MrplxRwnYynNfEHPd7InB1JhEeRTTe0jPfLshoyVuTjC/ViqwisqLwu6PG
5UVIrpg/dB5sRXOgRqSgt/9uEmdvwS53zTdCzHCmKVkETxh4Wwoob/nRSmjiXDzVF35jb6yZNIcc
EpCqiikDaJNaAe4R1b145nB1JvMV0Y1g4hnqoopHuI6HSFni0AzQMEkUg+aUhpykVJRMW9y2/EG6
W34vMhjyr2LFUeE5lwh+/h0cIbkFomnfBDMVUAgaXuYpLGOMD/eZDWnpPKDhggFWCYUTYpY2eEFr
ATyMgqICIlggz6d5/X/Geab3WQUX6vBLqmBoPOGBrdoOLs8zGnumTEmpG+hE7ISBvAd9lN7m/CDb
jhpMds8ir+yi7u9YUufjGlRXG6UtujjV0gM6KaxQJI2lEbx6NAXI1uGzTp2spX7TqiDiJNh/+PQC
LW+sro2aE+ZlvuQevBcLdWmDD4RldCcldr4qj30ex8uZwhc9hlhvXyVVnQWLrTA563egoNaRDf3z
U2Xruwl+nWniTs00yFhvGYFTOs7/CyiiA0ajRHGES0HUrL2/OBFTjDvuFNq+eknGwdU8K87T5a3Z
jIyy5OfaTjuXzEkN5q9bHW31dazp8sULRRnhxApb2ndL3AQ+B+5iSHFIQvzEffuXd1up9fo9psf+
s6boOLqcV8uqVtoDBBFB1PPK9U4VGu7sqUNzh7MqphNV6xs2ooM+csjIxXscYa5U7Hy0rBE/QDXs
lVLQrvhTsJti1dnx9rdpZF8YDcNSd1iLt+rP2ArC4QxYuDEjBBBQH0BLHtM4AmqYmeEg2rMdGuqR
UiW1tsYWiKQH8LBpcaM4qCuBL7MojWoPF007GTOo+WBI0kGob1gZbrnaE+iXuab5sz82qM+FJYsT
ANFJjsEHHsXMmH/BfXv/+PdsurocpnApdspv8WAeW5tJ8mal+E9KKSwCWdnMz02KN2i3s93DP2yh
G2QyT8Jlx6C5XjRR+FVV354EIb2IA/V+lq8lD9iFqf17ldEoPTUMRg28fnWYkKG2qu1RVlPg9PWi
xGSPV/mPHFHYekcedrzIDv2beR5eglkT4b5D/NOMuSVc5XP3h2Nu7HvllTcyjbt6fYHPOXh8r6mq
OIiYu9l29endMWntcOgRIkIeroLHkSE2Se1/THGWfJZlc9BbE49QnD1xHbNJJSLSmBnll08ne5Lo
mMY29kaw/U9fnw3tmhgepEhrjwiVhCPgI6OlKTEstkbrZAd2Z1OJCmR+TpJpQyVktDE4v4Ttb5Qm
Hcs/5d6Kqx7wYeO3hNdLQ8E4wBguGWKHMgmZKM07DnZ5fiHiSExBGYRLJjehlqeV9kU6mSrg2NNq
5PypITIDI06yM73LVFwyPQXzc2uPUVWSGKyKpMhY8iPGxPlBSrZaAizco0gLwKSSHRnOa7chjKoy
vZi388iEZktRMYrX/89lJdCdlgNuKU28SiaJuZJ1ax+zZ3aYn9zro8HK9zOmcB/ty4u6sH2Ops9q
ZiAA9+IthGlADUEgs8waYnP1CDTYDhNc5uw7rMe3JiqDiR5QSOni5RFLvGP3VvlGnTzaiUmBa10u
jOa39fGG1GY5f2BWGDOqPwmlzn4CvmY6nFaiow8BrJBVp3JxUFoCNEg6BCxavMzlAWBwxxnO2+Os
EfPdwRewriQ79+jYDjxt7yZHClh+qEVeuY3hg+aiHScEDt/QTdj/7IevZHuZ8Uphdfb4N19vl4wo
GM/FERNtwisdvSV3HjWzoLtd5MkbTdJTIEl4yCdb/8h3PX7nzIC3rOE/cJR1VIXmYOUGYD2Q07qW
1Vt3FyYblSQAaEEJwC0PaR5ysQiRRBQMeQKskkXLRN2GKt8Y7wh0Dkn1CfPBavPXHJuB25DTCwUO
2zsxemLai45XQv7GMTooyuk+JukUWJzpEAkfsRYEoJie3LLHkdwAT2oow1K3rXV2zeTIrHN9zOEc
PLh3JmWuDAIU5gyFWRWm0mlfIKu0a9/RYhrqkLnb/utGvnI5YX1MhTlQwrZdkkCrQ9Tm6sxrMGYu
OjTnDUwUY0btx9oz2/nIyqEx7Fqw1s2XZCTJphd9/+YR26ZRtM6q+ajIvyGZsekA3QbUlCadPzDr
l6tKZplibUJPSKLKWmQKsReiHTuVIhWAwniSfqACfoLUNkOoaP7Wv6GCAwG4GAPhBZtExnYMkgJZ
qEqszlM5+JXbqJ59LHebloaZj5T9XPfjzQYN0vnUV8RqsYYFWYS8C7LyTklfTAVh38EK1PsEo9EP
TBhhneP6sSRt718ZtjqhAR1K5CY8W3x6ITW1TY+AuU5SE3wK7mvaGKzj+W8kfAYs4Op6Oapp8O2m
Zv3ny09ahfl6mmheeKuLxILNB2v4/xHo/s8+uqu5JUowG+10izbzdwZj8PMuz4uEEHYLubsYL7Z2
qRssErB/YSRZGI1NUS1/43UJH8qtrgDMZurhwW4aCJ/1VLO9v+i+TENPCqUsbCVB6091TgxtsqvU
qYVytChheKmCWsHiSWbdzc1kidJsXWQVl4t9aFxdhmRlMJmCwGR4lSsme2AyOtWohrGFgGAjZckR
Qx60FKpbGQ8OPSUwq2gGXpITAPxQ9NWgulvlBKY4rhbltj5yHjAgo1O0m7Bwx/hC+QYaQguW9oFg
8lOjGcHp/KRmxbalSmdsrDT9H1asgXeJ7IbD3kwaXj8rbND1SkJ7ZjH4YWxmXliI/M/RH76Xwrcn
NbNr9Ot1+QSIGEL4jzyoq98PQDPg5bxKWEeXEt0EyyOjgWv8WBvmffTa5DjIV2bxl4voj1HhS5Md
mbwStOHtKixCGA9bAfqZlUbFBKYgnUprc42aFOUseSyMukJRcFo206Sm8B4bHoq1uz6+jgt10M6m
y1csop0GTCPavzPR325Ittu4qD+BKDRMhdmoKq9ADhN7IYFRioEfe5G+dwCe874yUKPbz9m9owlR
Zy/KMt0F46I5uSTWYjGFAi5WZ8PpliTJ7/nUuz72vz0N/JoFkkq3fe9Ku8Mv8OvObWflY9zayJFj
NSzeX5ixZhCts/C/RundzjqT91tCPntAyVHKXQGDV5OG4cflGhmwrCT9feAegIYz36+tNnODuvW4
LejHKxnIytPYmRuHAXbImD86Lbh/H9UKJ92fxFd5yaMoSA1gOCJON5NEHBzIqGHd1j1gltaWKKMf
MaNL5t3U/H+8niKDtAeinIHD9XQ2Sc/Lre7A+2nAk8aJf4zLNyOUykR8nxjidcpZq0VIDdD8jwUB
LYyGEc+TWCA5J630JrzG1mD6LDxVUzuhspdd2mxGDYhA61jhhAVk+tvVTqUG+MPuiYN4i34l29ye
1xngiuHW1QUA9b2tKIB3tBvwQED2A4rgfybjf6Dy8rKA74UcMSUzDlFBJ9gD18+E4PaN5S5ph4V2
mwdpnBI3iWKfpCZqF901bXbOjT5N4RLM+pUcZ+cTgccynwmmztl136MDBtijYqscQAP1CF8DmEZQ
xd3zFJT+e8quut199NLTQsL07ks8bN9MpBwcy6Vc07zNxnzr6ypIvFkfOYFptjIE13AlYH/BhNlD
UHiSBCsa7/L0RgnLmtu1Hd8wkSpfaYLyX/2QhbnHYYLcQQrBHttUu8yI5PE+p8E/6D/4/uSOwqJ3
ylRLfsXfj3dn/O9rzG0YNmJ2ScOkWfzkoc1CJ2WDhju/xj8gocmJ8SaRHcpdcrkPmqkKmjkzWn0e
GCv7gJzfy4ecrDPIu6gY5Ku83ErVuG+5lmS6JWLKeGtWUHn5KxRi0LWJqlb0eIyxSCmoeL61Qn5N
/LlUzTVQhjPgwoIN7I0yJbDAac6q/dkddxGDzlLqtTzHWcf5egM4S8Hqwj/KA4V5htdtKHGfLj2w
6wITO3c0J6KYWK1WHBnB4GvVSSaSZsBnKu0YeMMKKgQp1gzLiCzQcLSTy3YUH1p4IGepL1wvY0Ug
8WoH9WVDxbK2JaGgERQgTqC071nw5Bv9plP6qIFzclUXOCH1QDL6dNN7bDUZjMG4SX6EC5A7wovw
5osrKKa7ZkxfB2yVClBr+FpyEwLM+SwQC6Dk9VfyBpcvU0AqwriZv3tSdOKwBqgI4gc3HJin0eQT
vTMqINYdNcybHs4wUnQQF0raVBchNuC3kCU+/vkMhfAsDX7YyQ8BoKGb0ZYlqUQrR1Dk2zM+T9M5
sqS9iCMkJ1PEB3SGEKjbTPKFSg3mcY53mOSMXwAqTipAUOl20474gFgmfUc4mnB3A1DZ74sE5xPl
WMn5gH2WwMtEU0+wcPkl/zoTiouF2gIHFuTrdmQu+eZXNGAE9732gTrWChywX19EyxdcCrEEhjfU
19kznNpfBPpa6ElNIFeX7c/ZGb58T6JKKMdubD8nLwEt4JOTubf4sJXSs+QwkgvDum98YVHC5EOu
ckC3HrFb12zbs0HL/C2SXZ1B+qgnffZjYqH5RFTQmhUvPNdFGuK239Bd3nXgGycJHEBrCXGU/QWC
mKIzBlOY6ov9BFuOuYJS/fCUbp2B303SuMYFdn3L7LdUv5fGgRD6qC/7AH+GtModegTu3OC8+26p
1yKzwNXyYqT6Z3OwqPzClClqMgOyftSrwx6dCpsnv9MKKKd50/ljGS42gjI6pj/+XVMXe55RM7ZY
zZy0biX0Ej5OSYjUMEYeJg8PoiYs4dnDc1EqqTYCLxYjeDVkAg0fcYKu9Fp2P3a857yqs0zotwUa
KWLh/KMg4aqNdNP2SIdNVDOT3tAYzQJO4FQvqkG1hQ+rsYPbUip9GHYijkeeShhr4mgZggZz+Om1
XesZA81nAl0TrokoVHpGmDDv4KlHDV48genMhP49CTkrthPSpTyeuiASrPEVBT4aT9UdRmzNGxS4
lmQ1SBPxlmoTcH9QQISNw+cN5EvaG5clKbfpmebChggrjhWifIHMXnPLDu7poDvW3sivZ8S6ONIn
3usUeR74u0yo67o2F3iJyA5b4FvW4CsYY88anAu4KGD1lL8K6qEZbLQ0/v6RJK63ezoJLkAd6Web
fIHx54VWWIKgt6JUYOHGbvYqnQvQONyRd1Y7L7O25YF37PuuatutaKX/wsdlo1yvJnX7rcvVWlKu
4wOAeiT4bKErHJnjsSgG0Z5+2QWipdPQxABykOcb8A5JOCk4GhiUNQpsm+fQIZoWllytaNp2yxJ/
eiOW5GP2DO8NFbreEpDfin9+xptKD6bCjhP6hh0RvsoJNtgtE53YCvaLcL4E4NkEX2DegL2KUtJc
7TfRpRQZyk1Mvz97JJbIbGZEuq4nVFaDlEU7iappiKBDa5BG7k7CbBwDP8rFXL6wCBDwUHbt2MOo
JIMIpvy2fQNrX4Sgl2AUl9aVr93NGIGyEdXmXuRCJSASZJH6XXGeu4lI5vcpxVZhuhYrGXTVE2Ty
LujjC3y/vJFzwcrEGq62UKmQs9jaoKdQJ4z6QVp19XZMNpuXRbpGByVhz8esJz6oKy0LvriOqb/v
xP90nv1DCsYAwHXtcOCD4+gqcJiLVzaS1Soh4951NPYH0536NKmLB8J7N1qvLJvLndhr9Xn3JwCV
VNYHMGDE5B0kfAiS88UCiMxzt2MdSDLwXGX4/AP4s3zfc774Hcs8pjzT2aqNVcGZMT9fueQVj86Z
2JstaPmL89xOigRgugEanZs2UADMYNweGf1kzoaD3bv+bOjb9d5Bk031sii+XJZ1NrZaM7ey3gJg
H+7DvbsgLfFrcIU4JzhOElVeDEkmIXBziETebe5Q3hH7UpyeaI+il13ibFDoB1HYhWjNvyrK60/5
RECAs1SZI8F8eDuX/kWbzVIHbgY49b0lPDbG7V2ooSNHa2JOorlPLdaShbSSkZ1JjPXT+D/4PcH1
KuNmkKLecTLtOKsMnEmPtJ7s/gkfXyc/kV4IpeHzf17vPSplWUFueld3802DJkGyKYOwHLhK9PsV
T7/8XSlyi9IBCEOU2iUEOC5FgOHFr3QmEY8KCCm0IYoyNDwe0TMldHiFhHibqD2EhcgrMRgNvwPq
Oa9sC8bqZy7r6qQCxzifBCIYCZj7QBaAYuevnKg8ehl+G+3TQmswgPi37kH0sfWvYuL0c6tQhLpF
nWalZ0TlMl7yN1WhvCoGbwn0aElXVpUcea7JwKrhvRwtjhasD3wBdqa9YRVxU8d4uqHkP0LY6HoG
B6ET1L8nbHswm5FRArBx0NkHYKXi6ilAelAWpn1J6bPNKGZlepDjWXsAb8QB8tPf4w8k4RDS/UwW
F1Kr6fw1jgvAGDW64gN/nwNAjD87PQNFvJU957dyTYkLYOWB2uEYYvQHWoskjVslwSWrsu+rul8U
p0LvCVSmVri98rm0SMXHutk6WJsdijYNQZh6KfxFm6oUJbXNAvM++6XDdYC0M3A+o+X1Bl3jQmzV
RzT6xYxhiiD1BuM29DccncFBF77zhBzyCRZhTr3ArZMxGb8Rn6voJ/WAtBrEUdm1UTgO1BwzbKFh
fU8V5gJI6QuEDYcM4JNUSj9hN0mF7q3OcKxn88Er6SYAAU4zO39MKe8ay50re6i9M/d0gEFDCC6D
vZBjmqiJAUFKb7c8k18oXwxHt4RFU0hWx5LDSj7qWgvGYU1dQ5nKhrdsH0cTk39sFXznEMVDWtl6
qJO63mJoaiKLCzH4LdGhD7t0s7hG5zDaCyTrWnl5GUITHohIBSJ1ZVK2z+O+UBj6/GvLBM/wWpsc
cGdaIvtGZ0hV20zFcnqI9N9W04Ms6rFxkdUOM3YHiVG37p8hU2O3mJfumFeHtuUD8xw5jgZ6VBLJ
5tWlqu3McrTLQeTdrdxFn54RJHybr+DHq1rigqXDNSmSitREYP/JD9as8ZW7lzZaL+44b24EufcL
X+z6v8kfFvyfvC2xFDlAhQq63saeU9nWxwKkp02zSSP50bclZqYgN6BSQ1YgF+5zCoG88ZHOeUy5
Q+qGFxpIfKE+BtIIF8rKHj46/IyiQRSQg4zs8koZ3oVCyQGx6yAgrBMMBDD2maiAcrCPolbUnSB5
qUHezwVobjx1CaQrYoc+bh/BWZfXtj3ps0fyjUYU+qZqMlbE5OSD6ssZwx2LkZr8/IClPMzoYql6
8+BvmQsmu6Nkk2vMQjvCL8T6HhKtZIDJGIE5NVn2ecOlNry8xzypBlAAEYGKvN2PnTVCD2BbEkN0
VjM3vAk+3aUHSPjoMJmBJuEPHjQC+JwoLCgJCJ+hXbk+6mmM2lWXBxIt3aywnX7C2/h7gxM1NkbB
BZOZ7jFrMIptOAQDd2qFazQ3NjDoCNBpWLgQ2g2xTdqkdXyQLI4U1w7346tm4MutF8C3VHLFKFdh
haYnBFAAFJhyYJ60U1vvdOVY2VF+aQ7eQKRzyb85EbrbSzCZ1xyDojbJhxXOFHtEC7vyY+Qi0jTm
Z7Zhkq6sFxzZm8mu0Em6SwUpT0YZdOTNtr47ATGIyA9LG7NYZ/6m0YW9Mpp/cWyyjllupBwwl/gU
aFp7drNiQNuXQeGoH7kb0J1m6UiOP/MfROwETseLO0CLpnJxyJ1zQ5hP/BvgnCaq92xlXNm3+Zwn
qj3NGoGgy+7pPPrSz5WANTFO1ykbP1w+6nFOm0mjufHJOgie1B9f4HVJvMmVt/da8XS9WDJlPVE7
ztWiMYWFSu0ypDbhNm2O7q9xxXUJyYOgB9LH2DchYfqXMBdee+f5cL7mw7BCLF10PGCzLBi1tyTq
/U2AlwCnXe3GE+rU+Sr0HJA8adZ+IQsMvJKaQP1ggZyowhbuwE05M28Q1mYab9GSz/zuzBhxYc41
CDrpCn2qvat0giWXSJ6ggSEO1xoSQPOJnumEhY5Hiz80fjNHQV4n3n3GA4ZGhPxdGsI8Wylzmx2B
s1Nfvwte2ho03nOn7mBGMZIJDo04EVLaFUCw2AaDtbLTqRt2lteUWEnnMHbCmtZPzfHjgp7mU72c
jD0yd/EBdLS9Ryj+odNX/DxgmUvo9rOuDA7zi4Bwi0sna5s4hYKI7MVnu59sgUJWizF1sQVsGR7q
1Xxm34EEdW7zDuuvInqQS10WG9gpIyebMIALoyEINXV9CZ0QALE/JQH7Wd32T4gzy4ynmEvn91wR
r6M0cSkH1vn9vH6RHShr0jRGbeEmJqSkfOx+mof8McSirQX9Lc2TCxiEuPoKtBhkYrDeV38MJ6uF
UItPl7m5+azHiG6dvIzRHUoS/NRVmZ6E47a+r/2Tpn8hhmyRIc/r4XGE4EJmWz4cIE363atk0n6z
3pSnIJH7KKW6ZZ6+owfg7vmYaOvFtavP3VosyBm36u6BRCcmUZL2PzOQzNbAulmfWhvyusQk1cJQ
hv6TiVH0CuLMhOTM/6bbfI+jVPM9YEZ/xILbHnS4etidj8vwNX3aM8J/RGWo0S5kzmbIbUJ2ZW3L
6TAm3gwMviqHR2YOdE5jQtoCu3cuj1khXxbUZKuu7RqG3WJNXUhEFy7BrXXhKrCYo+qzJh4CH/0H
TryTIMVYNMwaDDx6PcIsnBciNAlU/ZQTH6Wv8MREcKVndLL4f90/q/vK62h+Ocm7ahp1DDGCKHN4
eK0MZvQv6Dmnq8M4tGX1H7aOOYskOTbV6GMt4kMUgSKU9Vt/AUQbVj06mJsJUqxJB6Wx0UqTHVUV
VL/y62z+/1EL15dz58ZpGhzcwPiCe7W+odGbw+c8HtlNS2Tm6tjctDrl394Xmi30TTV0WtoDAJFH
hC/r135p8SwlbGHjzKrA+HBvIbeu7laZPNVVN9cGE0xKsDIfhMogbf3kxgxITsV48VRBkfYnGjGR
W1mb7HR51CsVMRj1jC5qtSgSZNwgu5UOc6xCCuyTnEAzFEnAAlJ8rXKB2md1B6zA/PfuovmvOnaj
Dqu+pPK3qNZIU+l2y03VXgWbofBHT87PcczhwXfsDrJhTKGnXAI5GF1A+u8WeX6OPJVFXKc6ywtk
M/A/PpjSyH5bek2OFHx7Pk0XejS+eIdgMyXah0BFJ7zdlvRWachtQOhOPEE5LxE3vvEVIM3sIP5j
UhKTsWLb89trFsrogwq9r3M1wOmwb1SQwxTFJIJ/KQSuM8RuouSLMsPDoR7nRDdj2rpfLLWEbW79
O758ZSHtqoJfGLbKZfWbS1lhgIyw6kQjJEtV0OXuOeUSj/uPcnv4X9lcn4ZHG+JD5Ml79ByNHpq1
N4IVNhYLv/0PMJ412VN56Ii4B7pA4Ihh5uFkj1o7jiJa/UWMHIOE/nf0EVD5VL9EYgunOeaYv7kP
CUU/D6eG96GhphFBrLFmcDeG8J8BSHpE+EhtKmQI+uhzlsvtermeet2NDsX+eSke4gZszhEp6GSi
4YjdUKcN27TXwyCMawP2mO9iJUk7J9AEQPTKmbHox7Cl5ais7bWVOMXbuR3P/HxSFGgOL3rJUuz9
Lhq8b9VWeko/7zXiNmnShBfGejVlB/hT0YIGIwlf7rmctqIguiG8ByMS2d7kd1ZPYbfb3nXBpIMt
g75BBLOakoxofHNIUZp3fT0HuMWeb1v1Y8PqJLtjrPs2NDfRqBWWbGcyYbbsxhfFEP8IK9NTOhGw
996Zj7HAZss9vwDM1V/pcr/iMYwrkEycgib7E+Ui6M6JV5y/UW1W3DZcWQOuTBdBo024VAF0Ojpt
t1lsPR9P2dYk9SJwCrC21GpKjpvD7sKP/cIzCe8BNB01XUTiyIZYeo0OSuOhGV4w0IPK++3mD0qi
MMNxTsncH1nceX99Z0IZJaYxxX83GNpcZX5aHURmwwr8/fuXxFW19vTEN9u5AStYFOEW4EqyKtVG
P3N4jr/+ANUgUsz0U5i47zQVszbGkpTcFotKyV5GanT52cTK6CJPAFQARLi4Z5h4xxW0pIzlZehX
l8QRhLBhN7GTMzvM2nwQqAm238RT4JokJYvqBallfRD+bXVHIiJBHHfsukWWO4vTZAzXCEgMuUk0
xCvu6R6FnfwkeGEqINyomupXc71oTowYhDJhI7gi9F1HnQJ9edELexjuhg0Ju/uxfmaxXoo3PWKj
XSqmj+Wx8Uj+gcvF8q38PxFn84poPEP2bc+mmSmVhqKQZXKiqjhFReFKB+ydDy0HccOV73+lyznB
UROdAmB82ZVOH13e9Wm0ab7vMusT6OriY36NzjBsrDFXSV2BCkCvJShjDth2kbX139a6wNbZsp73
H/XKglRh7EtrN3g9MmQlk82CJGWPrCwkTpWc5rfJSox6GMcluVnz4W8Q2TNEVl8XfcvD7qihczG1
M0lbr5dt+DfOQ2BjvSi5KyMB4IBEgMiIArilNztUgNQ0i1oR+WVFeqof183qchFZHcta4FRRNOUy
PvebDBEVioPnsoWXkuQM4pKCcx7hH3ouNEhlzsmMH/UyR9gEE9zSKKwzxsxirEVJJUxL49hxBBgT
ZHjiyk2YRkEIsTkn9MWCu/OLi0SnENzmDXx5cQNlydDf37Hmv3gf5TrY0yNIQUoevSZgG4V3bG5u
GptlCEa6TQmcWcF9MFYyogtQLbelpB2F7MgEBfSHMKGvI59waPjHOl4D9Y5Pe3qA3/v+YPPb1Rb4
CvuijjqftLqQTHyLbZIeFLh6XEnWYzsy36VelQ4MeIrI9xuGf4IRiBxsai+QUpgbF2Am2MjwRQeQ
and7u3Q3ZlWhcpqGfGuc0wFvJh5HNusUJIVHnLqAtrE1Sm+FRH67M3pQ6N7G1r7WGON2ZafDGjqa
Ic2fs7foNN7R49UDc1XhM60Igabwi/Rf6XDHR8LN1ERrZj7W7EvjOcEuLItFjMkYC83Z+erKLz6x
qCkpS3CWomFXAxSa2+M1tIU28MOUpXE+DbRfyv6sJsNqpzJ21c0yz+xvQ9pJC92kwmPaTSiuYsFK
DflS+FrLPELJJJRlDRVBBXczsw/KwhJoj+3kmrtp8KXoRlu72v2PAZr3w2VN4i0ZEAILT59THE6V
MWOjPcHVHG/K0diEOZF2N05+D2KEYUevs1tkIXcc+2QSFxnAU3hNXYtLv7vDDKe0vFZeW9hSjmg9
LySR2c4fiIl3px7cqSnDTYdFfaXYOrYJ26k2mhuGopeBKSDvfBjyNsnXWOnm3fsL7oklP70d0zH7
vUBmSRDlXcWYeO/d9QJ5yHbttoCLZfldiyToeYXmbVNdyA1ugg4AtosXSxY0fqpozyWejlzO1sey
OagQxVFoQzyvzTxya1ce8B6lG/B9VPrNbv1zw5OmRylPrRx48cafmkvA9s1QcnhZ0H9lj1i+mral
1d4lDn8yqt0sRIVDyXfkcTrC+XYL1dJnziltpJ4s+Hm4tn/EewLWkdftZGzHmbetu+sQhJPP23yL
2aCuXEc3fQBOTXtEcVsDDLCDkRy8HGRALiv5+QjYP3CqP55A7K6ExFpdUtw33wHHtTpZOw/o99uT
9cBk4tV2Po1kUzQ0NNEb9ACkB5hBoR0CLXSSTvD6bqUSFSDScH3dZaF6Ftq7WkC/4GZBfAxoXA4S
jAxEx/yRNYxS2qcCbK63UJdi/4K030bWXUor3lqBbdpjRDYNmR7zXsknuxJbA57mPIwivlTpa4xU
GWxH7BKEjbWZfHLX3ArQkciT1SkpyCxryDif3a2s65M+GSuarYFFNDqkgpEfBwPvBulyMgavUjk0
lYQ5cP9ZaTghagBbA03ks8yCEJOeXaD4UhsvrY5if5ZQOxB1IBBVndAVJfmhU+H726rnxd1vI+5N
D4PhEbZQ4/Dm2IM8+z19tMYeWUEJoGEXof2QreUvBiYJxBExLI8smZv9xA5NkxtQ/TAvFh0CMWGL
bLp5KoWlQT2T3lHSnKEaWmz3Z6CkgKqyy3CGEIy8pQXU+8kHcQ5f/tRR8wP3vi8d9Pgfh1ZpTCRh
Jk8mClVDh3us0u0K4BJ4dEZXjh7RHN0e/gsNfNUjgdCRqNhC98z5wX7UIo9PLbnvdSTbU/lgcpmb
jZ7BvN7c0C8mlhkpDFDOZ3UHgesxKa3SD4WG4xtW+HTPT2A9sLJpoGLXRXfLXqF0/uiDbUqD2q96
pXc6h96B8L63XJa1/dGiGIPB6011ER/TP6gXUjuMWdKjoeBseEHeGu7m58PstffAxpiAWsih2xc2
AEBizB8bfxKFQOJ6k6GyG8YijzXP0w3h9CZkzcM9uV4M4nUGAkZIPDvDirpQCm2QhrQjNZqZJdU9
EYElKR+4NSs/x2Z9bCG03lW5ofs7tM19TFGCQeJsd4PRqG/ST9j5u+mlsxhY55i+c2GAxShqAgFO
C8tv9sMV8Lpr5orsqZTNlsmKKJaNsHvu4cn3kYBNGudVuIg1XTYnSyEqIbvaP/UMdPS/9Ya2u6WM
qpeyID67V+0cD1+tzNrRAfLkmnL8ardkrcgZN9ulepOkKKw68oTSnhf/TYqULe80UhWoG7GjOk9G
cwGtEqjAuXr976pJURF2h1axFFU/jPPDTpHT79GLP/HOZi0OXWspoPFGZZ/aFyAtvcKk/igC2gCB
uSFR8mPNhBgAPPK4W0GaoV4aPSft1fTAd5Fr7zNxhYo54pyCBOd3cOJy3L9tOALtLWp4eXlGQ4kU
ZAW1mUxbvB4DtMUqLt/NSJ5pU1Zp2j7KhANcju1TMXtxf/ycBMqfMa5gkVGyyy8nT4Sqic1E6rIS
YSN8vcGdMEbQxML0wiAq7K3PJgoZJ220NomT57AQWvYnEep3LgZBld5s5Zy+FWR6uFrn7O2QWFe2
lYEqqNOvqHPCN7YemRT/rJrSso8OJE9SHUfoCC1fxuZVxZuKUYJTPzxD25ghNq4VuIjxF+DqYn3T
HBs9AyQWFkkC3czo9xbf+yqfee41uiEulW30Db1Yf9NYSArJLJH/o9vx59x4G5thYgVFATpv3KHk
C6Yu0e6bdwetyZ3S3iK/6/v9CnkGMJlgQv/lmhbyxkebKaGQZwxKgWaT3XAPHUEQ+tEb3eFS84U8
NpWPbCnwYnF/e4aoO0t3eQl/BaFF+jKsk/5cyxvbXwaXZgT8UraAJjkPYT/Eclvs+/rNbnSk94d8
Lqste8HqHZbVh3OLW7YgIiQhIzaEGZyK+GftSiWtI+FDUIIwUzHznA9rmTK9hr0KN7ykIQbApfvD
+c4EtY8Z7Mk0iuMn66em9rzz2Zlab3iru9Ma6EN9CWTeBtTW3RHKq4KXuKrDKISJa+P85YKV/8Rv
YbsiJ9VHosARwTKWhkvyEH7U+DkyZhHBL5gj682a7p6nA0OjjS38r/n4zA79/zTDHQM3ViUS7kCz
eLMW8yTRpEiykqZbhWN0d6mxXs2wq4eVzkdYahH19n/Nik5RleNI3wT/SJ6y7a/EAz4IusrkBCaF
RHqsfL3gT/okDvtTKu9inV5QMCx/DChy/b1CboThDaE8Cc7ZLo6hzpszvSpmRQCWCO2Nqi5THbHQ
VbABUbB9+N9zMdpX4stqH/NL0TiNsWnMJAOuFKQfZ+CGkx3vtcPAgGgSTm2ovMn7fzPqq+2zM+5z
C14mHYsdCyy+OtGpDSW/Sx9fAPYd+Dd1XsbZPcoi5YKiivwpl/lAKCuczPgbcer0dUsfcwttAaYY
v1Ih2Owr4cUYY2VZfu7aCyNSjbpxT07EY+9/2xkQYL/yB4Cha4qBqf/I+H0taq1tZhK85gUS7VL+
mAgZ50l/IdkNMRjX3VzS67FRaRWgnjFKfbhFNm/l6fU36zmanmvH4dlcxn8aTgMUWuhMHinpv1vJ
DMYli96HMI8gDsjN2ZfKlLxh3lV5SE9d3HujBYddSuiNvtBFxbVvkOeQ+YfmxQ7wJOap2REVQQj+
VARD3bAKPVigiqVxfq5WJSgT9gKPpxVQrNeWB1fbHU9u0RaTrQGbq9COMi9LPFWdKSMz9p25F8rd
YB7zNS87EZbxp4uYGiUn4BiHQ30KY9Y4mDyAPb8cDVrcMsHJursCmf0fe1+KJxTOQhZLggCzTAk0
jTQQ7E7fxUZZLo1ajt8im6JRQEy4rXK3w1m5u9syijAllXU2MPrDFqWIXDOhRM/URLr826hRfpBM
WmkAs0XbK7MY0yJISH43ISeP1i/D0tmKD/gGoipCcbasOzRClyt4AEAtuDYF0O4OGqdRr+rnYPfg
6AyuB8bJWDFOxXPXXcxV4qYaPB4ajEzmalK2iIAGE3Qh8EGUOE4C+/AYVSvgxgbegQtpSes6ioi3
Hon0H83BiYnFPituOm3P8KB9fWmSUUIXW2q47wzgmGEBGr5jzd85hPhLufjWXugC2wedaDIKOt5l
AQtyY3t6H4EkCXiElg0OwsO/VD2ln/NFKGzXzw03Bb2vnJfoK18svvKOmm4mponZ+F+Sp4tI/F1r
i9c2QjuC0xges5MCgb0qQhw2YXhf9/MYXEkPcZiZ21KOd8wQgky7tXTBtyk8didmSIuYkSGL0raT
pIbCfb0BRkKd/6KJhHFw3oPnQ+D8poPvbMPZLr9RPMB1d7DOsBOXlscptW6JifVbdtOYc8UDuP/W
txfIP4q+OiV2qzzY8YY7Dhrx0fW8OAs+MXJd243IWblY5hcMqk8Wi98o7/ZR7zntIEA2m+LdWT9W
Qi2RNdTN2cvOzok6DxE92p73G8KU9RLxPs4JaOhNA5s2BelRmk5PuIz6NroB4W7jd6ULpHLLoNqB
a2PazPcV8FEYU7W/j8/OoWVS6rk2rLxAKPlOq1Pa7C+XJzI4nnuQuv5iQtm0QU/WwbJtVguNoPlf
iBTGZv0TPwfM0De2UJ+Jc7qDASExJsSaoZjpsnKpZZqI2k2/4gIC15btGP4sWyMYhfjiapn+ApSk
l9gtfZAuctlquLxEjJpdxDSE8PM6X5RJ+VBi9zjMCSJntrsg7cO9nNT9TvLg8Y0MOE4keOM+EhIJ
apta1OsNjabNRkLY2L/S+t9TgHthdSjFF7IRtRsxTDEcevNcLfPSXkWmgt6OCvO8vAI1w68nMHnM
tLqAzuU8cBoVU0Gz3hL5Lt4AsORrtLF6nI1VTO4qupyYqDftM4m+GRDKiC0xQIZA5yE4b99ru8En
ZTFY4HNdSJpQpXJX3YyDGbhtlDBIXnScrbXm3sUBfvMpAnta+yxhSV34nnAwBE6cLqEenzG1RfHl
0t97Xd8D8qHZKEwlQ2eqXitYoZ94Zgc8FrOgyQOrOu3OJ241mGbBlrorBV68JlmjAySX23nT/bON
wM/aySjVzH2EfZne58wcSvL81cvzvuXlf8nfJkK0THFHAfBXBpQDrf6MXZ2/gYJu0WpCgxmXCAxM
zp1Ja3zvNVz1xJneTYgosiDPQIhH8yniqjuDJ+CJWlEbQbDA6iXQqY9arbHs+w8+FoBHmuUXSIPT
yjstGdglh623L2Eo799IgAqB//G4QyN+HRohDVuW+eS7F70jGGjjMpoxE8WhO5YGVqK8SGEJjSQK
P8LgM5BKmwqu7mdMz9hmrWODmgkdb3MWWhcq+0/x4S2W+mnyQ2rbTQcYLkIdBjCU8NYl7DZe189/
moiV3j+u2nM5dBf5NOO6kHSWIShYdYZbIhp99u+zHjorWkCxr7nOvkGgyEBSz4MDvNqcI3i2ArSe
3fFcprEM9LfPp6pjaW6yJa6evm/1RTE7TcxBcz6MHPmL3so9zC7VYTOfCFphlpfKY8cACQKCIrDz
9xqimexDqVcc4mwrLZuN3IQOHUfJdBQ53efobqlCh6YuY9A38K49hahcGW7KETQyu8LSlXbmsII1
tAWxyiKC1fB05Rtk1rWFmXQ0g2XBwpI54KoxsdW8gLvmeQ/b2/BnW9TwOsacrJIZGuKNVE+XdpIX
YOLvB48fh0ZFdzkMm7d80Ce4CMkLLfQ+bC5uq/+MV45k8mAyS+8fA0dtUeShJvuMGVnKWAIGi6Gk
oAMa31eY+ojR47Z/PocR4tuZ9v9m5/aTJhCsw0nLuifXSzWOdUs+VTsglcLtXINOuVcul94txsNu
kqCBOlnQJ4lcxrAoxcLzAwMERQxuHzFiDjxiBAOySBl2TOtcI4oMfIrxf6SJR6rgNx6svD3XLNtH
eykayPnXhd5ixxqHm6eCbcPxxN5MBxzHvPHJSqaose9vIcAPgwnzaprxnUlpq2CLmdyqxU3StO2J
6Bnb5mmHxJo0hyECaAiRNpQzfCj35mE5Gh38XX0RNXvB+NT+CTXm+PhRWx/vlQOxCXdq92AnU+/u
hV9HD38A5wLUGkMZLQBvweXWnNJYVWzuMaQnUsStN0YCj30013zauoSXokBF8N3vttIQD8FZ2p18
PVEkEwW3qGsOx66ZCGGxHyUkZ19fqulMIOPaCyu87DLHuKjBnUPuMpA6r+yFJBhSH2WoFBz42Dju
UtHz67CFtLCQwd9O9rooS56C+jJoGESP3+ll9CsZqE+JOb1hicc1qa48XV1KPLbn9RajveMqQDUA
ya5h1ezM0TNxXThpTxDFVKnx16wNMYgPfC94BJy/1clqc5IkCFMRbl23Ofr6FaIX27R+DIsXBepq
yVD43XS6rWa32pU8REr92z1nqHyvgR014/qUjAmH217o0jiIl5Nj41I6ozmMpj9WYMFtWSrVmxG3
GL34szRovdqU5Fsboxeg94MtO0IMnhtwy6hg7GuUJWaTHLM8F3PYe/w2vVISOa9Sut8MIYFVJpP3
hAoNct97CmloKKw3sTh49nqePUJl6t8TdWd2Smnh4nmnSPGB/jItiWgHhPyE/9KGF944U+Qnbxe8
VWbGLkxk4ZOp6GCAlKsdKM/d2Ir99Gkaidp3ilH79S7SmVVppCR7Ku+fy/LVySQX4l3qfaPfz7UW
OR3bCcA1s8Jf85ZogVz3SBvrZ3EvCn07aDOLtBErreui9XW/O8hXYFK+J+BIvOQoeoPNuk7P0kQr
RazIuhcnSf78LkHzSHjYwWhZkSVTi+abGe9faOc6yJForSafJqNgHInaZ0XMbzL+XL0CdlIni2Zl
OiwAKYFyi6xaGPxoXiwbSrsEC+/bwnUGK0ro7OBXAlkVXVfJkfn1tcxLmZbF23Bu6p+AFB3TtEGt
2WIOLJ+Vfwjvl6nriSvCY0hWjVe2mQuPoP8yvQRsBbmK/0wENK/cE3GIs4EoxGNDeClHr968wLJ9
Vd6xlXwUhC761mKej0bOZB/rWfU1lJgAychEJ5N4GSai9S6TLwFPxhJy+365GUFbttI7nqmkIcKW
FB2lFcneptCF7XhGCy6BonnypBMdk3Yd4+cvoY+RJQ15pacD67IA2QmhMzcmczuM9sQvRBVHpnCL
1xq71N85JqqndrEltvk6/ylwUc/DpbledAFVBaEmPqf8XEah1obhXyfYc8sqtPrVEEY4LpI4zh1b
VoPRN1kp1GQnWfhmKaDCcSPr/hcmTedLlWpvqj+hzs2k2n6B4u48hjan16LD5HLqnLeT++SMsd9t
9gkXW8gdLlh/D084/MxVUKBVV+q0CIIrU+ClHKhceHV8+bw6hryeAcNI2Yg1d1jA5d+ph4v1fL5I
t4Tzop3SuNkntnoHPI5WIgM/7Siy/vQD5Plb9xM0fpHqTyCOhX7Qh2enXkuD4/0FWKy/TfFLKjEe
MApP/Wjvv/2xQyctOACqFdr/jRfloIfOjaT6pzcOfqJi36HLXYkjY63B+xFrpRpue+rgepkRQ1xJ
U6VlEvrLQjahjc/XDOuvk+r9/YNx2Csp7RqdhnDzi9fn7LcH+tlLWVQT7nAjNaQtnxiaYti+r5IY
FQLX4XMRw3STp3t7wJ+MYA1S1rnwwVVuY2XShbnii+StxdIOiq0wAJrWI7Duo39m55SBmIBTjrN3
t8sdeZUhiH7imOPvh6sWSBGmaBBl0+CtRj1weDDcWp7Hul2gmKFiR/OOoMHy4u1VZTkqJaTjaKet
MVhiS8tTvWJGkv9LYiV6+QBKqNeKrs3X91QKiSQPNrYbFyP9tJOsiBjJO7W8ObTU4ER03Cl7UbnC
n/E4T8V3mOYeE5RV4Rn0n7vXqtGxdRxJYzVv/nFtfSmIARte0F0Tcjfs4f/TITSjPyKLgv2FFsD8
HSqonWI3iDppCfOrkS7/Q9CGFjBxUprTPDNt+4mz9gi3FSi1hvcprSaJ8SbENDIgP2AiowEtGg88
awM/QMF7t9DDUa18GnsqhnyV4js3VycHt0SBhYdoPX9hwNkFRxOZlNkuSDZ+AK2mAG6R4PatSkcr
w1/Tjhi7AaLMg4NCHp1wE7Wm1dXcZuH8P0cTciSoi3GjvY8B5jvP57EdcvCSgaIrkmkM1ETLzQab
fifoUZaOVUeiTQAA6GyuzlQiuNM2vUrc+Totzwp9+VPLCVcd8mSVkBF7GY/Fv2HcOZ3qJCBRHIvm
H3Ba/OguODuXzdwwxosGRbJyV9q1sio08c36QZEQmc3u7cwhQjC1D33NE9VrqsOT+K+ei7+8AZfo
BEZmLIVW/G+neEtmSEipT1zAil1CzMtHYXrFajH+VIdSh3o2rb82DUoVM8AcSSEyXcUz8neDDSCU
e0jMfLGaDpMhCoiCVb6WsnWVFDl3qEvdBXrcSpqOmvPztDsf6ANreQ6tbrxEJIxTWUocLeMkQqxH
FZpkUm6vzIVg+Hxgr97yVzjWJNTtGuY7nf4iapQB0gtIs8yNx4VQ/O7RdVSkunMpo3ajWOUJSvME
5rXO06b0vcNCepP6pEsW/Aq8jNLcN/die1WOc7PquOugojH0aDEDB4/kEvwXH/6ow+TFH4A53/F2
rB8rS/vEXEd2OOeP6YOkGJJaaGxiKxpRXOhnja8jey3YDqegUbGyDKo9KZ02I9DRVGMbNsIoetK9
XTJoyb1oXlpAQumxmRgnAhBBH2vRgLVtN4KTUKjL0InY3Y17paYGj0UL3U8hy96qulvY+nrtbEAQ
dzdsoTCmiOiT3EFeg6DYA51D8ly39/kwrGQCm22SKQd6VpuKyUlwMAIV/BQrs7lFZYVXxLmKx2C4
0Yq8AmusrTV6ib+Y9MuZsjBgEMUbXwFDkK/c4ujYGHI+u2FnLtRGfQg0378fvxIbT0fKXqUxkVWa
7jBu/z+LcJQXRh7zULWFcdiDR8NXr8+8bRQoJasUmQo4ZNrNS/aPcmcLecFYCralI9qUbixoy/x7
e7DlNVjLzKuVgIgQMcd4p35JtKNw1uAMo22+TakhMnvWCep2JsPLe8ePyUsJAlYkws7hVVXsZFrw
N35Que8NGshwSktrW1SQ3D6Wj1k6ugIFmcj6CoOmBNvkJcQcPU9y0BVBE1+ObHItEFE31Z3fT822
cet4z5Sqxn58gvAmgwUTQzJw+G0j+8cF0Kj5OK+sdLzShaqkpTUjqVUFNDSokcUx4iDVWOSPlrQB
N+YAXsdA5dU6m3n66OhdfbNY6Ckx7C9ceRLIVqbP0YH0sQj2lP7AR3qLL48S/P2Evp6JYeCX5ecd
dUFFQu0g348CVXkRU8ng/buWJ1T02QDEFfsHFOaKrzxWDxJZFYkxIaP1IWrZ8P1Stay3773iSPde
c1B6aPVELJXtzGXOS8XUf/aZq95g3tHcgrll588SsWkvXSFEC42EXf3VBwwgXqFE6WdPQVSVqDo0
ZsbUWhfMmyTMqFQCpRYv8qdXvY9tMrb7dN5yS6LZwHaJcsIJ6HPkxviVJwG5Aua+bI7wbtQiK6d8
zwW6rw/j+LhHdki19ToBg5vBoX25jhTuM+mUWbCXg53pFzXvfMEmTQlWLJGLLkNpqItO/aofhhXM
AhgJ7PpKRcptMizByBKY0yGtjBPo5PBd3aA4nVszc4D3AF4B7mMUaT3OwS3Uy8b0R7uI9pv9v1XB
PNpijIR2HGxF4cP9fC8oAlOkRW1p1jhzlA5+mZRiwyngTN6b/u4fKGPX58db1g4USrIEJ4d53bOZ
SfQVfPMvqTB05c1NQL7oK29ENSo7W+v/vj2uwFk90p9a5+pgfncNeoZ52AyV7QKZ76SWhKD860Jt
WauoCyzyJPmMhPTuO6WLB5+c9uFkxX2YZqizIVzkXnVxZfs+g2HmVDdBd6d5DbL4V13IB7psJZLi
XQWypNZ3LdSl+UAeV0nchD7kepW5+CyacV1E+ZrlGx294K0E8zbT5LLEOGF+Gs86zDJHTkyBinrZ
1GyeNe6XIY2QL/69iGUKrPb1MVHzVgiBoU2ocMfJFrCeg6CbEvXQSQY1hE5MoFgUpux4IMdHSFUJ
j1sYfwCI5w90z9371dVuzHz/jmS2UP0YwkujxspcmPQLVRosbKZTJcE9V4m/XRpE+nYW5A3pNWTr
b8YGb6fg6juvX+jOWnEqgmNleiuCxikD6QZdNerUUAfk/57so1YteuTGoHjGFfXhMeQIOz+KWFdS
4QzuVNzI2pf065OoS28NStQSED1nxA+MQQnFx13FhXGZsZVf2gdPMKR79Ecjq/9kUOzYoCWrLCgd
Yc2EJJl4jIC37GlUrP9vcPCUbx5C+TrrqA6Hb4Eqs4d9z6akFXGXHj++lAAs2MY2WsfhvkXtFEF1
06Lw/En2kCZPc3hwhSqF/nO4QhdKPWJTbBB7xfU2o3uCQEYV7KYFwpWSkqry4SfWHMBWHbalmssX
NYsJagX3gnCCa51GkTdzACH3s+k+AOJNWuRp0MH1jE+Opk2gt0W5QRAng4Bfov3Mh7LaATLtNQ39
S7H9m9i/cgBKFmLMxGYu00oIq4zMfdb9pgikH+1y1m/2JlUHEpCqQ1ibiqV3Nbf9mZ41Rg0pTArO
6SSRPQlUN0ZPbQQnYRFi4utWyLibiDI9vDSfv8A3XKjHOX1j1YuPJHkrtjKXDHdbpTpiza7MR9iP
5Q93mhaev6sdGkY4h/C1vk2a31QtUQHNHRahJjKHiaTigw5anLQKJcuKf5+IfbqiMAFLhKKq6mvh
Q5SvRJEeYOUZh9iVUQkhCIGGfmtyPVZMgaXKL20WQoqun3rCFnw20l4fUyH2Qq9ocJineAZHGG54
paSeBTJZn7SkN0emKqciscDxn5KMysF6O/jlO59SoAky2v+7E5mhJFxNlBJ5dAqy0qiAEamaHilr
Qc9nQLnTl7hBa6/Pk+wV1V1CrwGXDyIGRskkEkdKHrWNmVNLChQtBosTcjkoWOqZ7nfyqEiS3cHl
srfV6SA5xyJF1ugfsdgDMT5qwb96RDnPukD2WLrOZZ2Qou1g9mW0RgO9yqMt9ZzJUEHO4c/bTtts
PU1JL9VryHTsS18dNEIrlfka6b5qmwG9DqeXteb3UV8Q2fLdx2c20R6luD0BSLo4Q83K0Bgvb32Q
J+3aRrNiDd+ANXgU7FL1qkMCvKm/RRi4xLuIQGrmaGoUimpRitNJro5KOnWSx7k4FgLp4s5/d+V1
/paQYRxN0QPUAC4JqlGNFOMydqdJWjnE0LDqK+VybkaZti5nQIXo5xPFyFqohxiNBLJGk18nrsoP
ZDE74P9AFX9eKdmNWQ3TmAkWAVKj2clb20xxqOAuC1+RTJ/KQ3srN6yuKodI2+PaaHPw87VXwi5R
5SUnVl3Ov+LndxHq+Qp5ISb7xJphDrDUC3ppU644mFCv9ZN7nWqbuUGMPP31X5RCHE/9hAaNDPSx
qi5Lv6GzMOHRRbyBfckI/HmfeQC+tNjH08IZonygnergpxmIJ95jGYwXsQjX9jMr2aCRjmEi6ob6
WXL+JBvooQ2vPaMIymSfGxYgoywwoDS8WUqF73mXWGFh8Y8pnFyMjyjepmDkuSYgj2B155mWcuU6
dpy8I7oDAFdMk7rM9tgbfiJ0eQ6sllylwa38HWA7Vq2a+4bWXnXCVpO+PS3EQwTV2ZciDataCXCB
IAoInjPzCdoXxWuGadXy7fMZVYtES9V/f3brCtMMUI3plRsNIuWAkI+UlcU3Wt0GM2s5F9HZpeXM
UIQjOIXXDnkjU6L7+U2FhvFYnJ7MwvIlGvsQj/SSRcllH2eRJdRcgJLVz07HSJN5ByAISE4Y05ao
kRTpouvuh8LCpLVdkZRRHKlOkpfZdQJOABNfdx9u/Eg6bVgltdbsV+QxZ5ZbBb3182CP4FLn1AAN
EmQU0aAVujjr89jNq83i8SuGE+CYxjM1rF1+SPPhDPjYo3jIllhMw5mdOlAyi3w427fvWQ7CzUeA
mddpjsr6KVe9DxyvA8YZYYMjblx0gweQKcTXi+ZgodI0ajUskOgPWV1/Y5RBHgrAgA+dqoyGJ+tF
w1sUMO9yLPjcra0d2Ta95wbS5TRRDmEnZN/Q5JAe8+7J9K/94zlpBeSv/80oRTEL2JDFuJkj0E2p
8hVfUwEzbdtV1lPUdff0Of4r1MaTGizrgBOzPJUBJMQ46nQDkpw3/YhoXpe++Obd0QQT7LPEkZv+
e54Fo8vOUM+rFLQG3Q7xfQnGU3bdg9DA5ZlwBpQOOMkvsXTMQh1VWG3/n/p1GFwf+exvFPIZdmzT
CEzrblPNnyvMdwQGtoDut1Dv5Q54VrfQYp83cheeixMfKD2xmiv27DNT/n3o1We2G/acqcMh2Rg5
VaYGAg/1rCHrenCrlzGtlnB6run+AhmfwigpqwZGS0QL4SHIhb5dLzQaBC1vfJITKYlRdOiU7BIy
H8mFQp52P2jDj94qIz9kvzkXAjqirzBbKa0haeW4Nea9TBDQIPton0rqPsELb1/Q8aN5KCswVxP1
XfdXp1B28/diCYzGUsFyAlXLb/rYAQHqHlKlOxVuU1AsEKExoYYeccX2Ru2bvW+U2eYYbWRedUre
g9xzQXcoOsB4wP7Lss8gYHzSi5CVcnhJ1YX8Lgj+BKFl8S12PV+V9yW5sMqXC7A+eUpZdIJVmIs8
jBqwPbsR4lWogRf+Y9pLsuGOo3cEhV/lPtAiwF4jcoSgJm5jZ+0Djfh2toTDTTtSnMJmm/4489P6
9AYAihKzEnpyoJTd4icOJ9CRovUhxyP1tiETiV1FxPXKtI8160FU/7P45uiFcIH3quO5L/Gm4RFF
i7i+gl4GMP7iV1JNeHB8F7GGN5yDYACAEkOsrM6ev2oz4/ldtVP49iPLYixyEFF4l3jPr8juri4o
sYqOyG0/06lY4gfZYqzk78kNo9uKMyrKtsQhj7E5q3+YPqasLVK0W01wnewIhEmJSa4bexpYNxbB
U+LbPAetEbBxhOJvTSJojHNg60LRuxwhfT6s634au2dA3NvT8fQsUB4VWsaEIK7GwoAmpeRb/4Sw
U/CGN2vQVHBakM+B+aff7377gD85kIAee0mCiphqT6n/vmrs3HVCGK5v0+hYwg/VOBr0k48kBS80
2u1jf900wQziATyuzM7D9FVC7M3gnS6WjUv8eJua2TvbqtiWBeImw9TGXWopaxwbvWHCBaKknhb9
SY2JmRxSI/vV7IFILqByC6o2TTcg5LHUaqpPOg6AhA8qGu/dR4I2mLcTilyf31Yc4BULpzbHwdvN
iooiWSTo6MkEOjH6ag4VG4xNnSJFICs9zdT7CXAaFfF4aVRSwHm6s6c+DRyz9Cblwmas2ewnyGVC
cWpHq767wtXheGFc7DiTvel172EKu+zU5/eQVih9zqvdMhOX7W//aYEhhPtG0OApajr+kzQ/VHtq
dFeVke5LAR2MpKzU3kvyrjb+QnxjTTGsAnN5x9nva2IuYECrQozQ2BaOX/owbYYWMGW50x9P0keL
OXeKr5jE8ZxTVThBKL5TH/CFlTxcCqaZdHhea4QhZgbFsZ9D7lMu9WPoKJu9f4xg3ShHd+1gfsv0
ReqURAtwDnJX1Mzhq26WovZ9q8rF5tq5pzMMjWYS0+z3+L6pbBDE9tKOEgb+5vIqQ2sTzm8G8oq/
MkvTLmZ+9tmISU77NEAr3s65VYAYflY7PohsxUG/YCOEllg+V0Kyu3vtrJD3/w8sD3+JakvnSo5Q
/UFjoKRgk1yogIlG3IOCO0UTwx5xocOXI28MktrUzpZwSljsMUt263mUdG5Mc2irNHG70CgP8d2D
JU2zfWlXkiX0PJ4p9dtg6ttGmbYyK9ANTmZET5fImunKzK8C9+JVeYF5MQrJOobN1oQnEvYYNkAX
DArpmgZCb4PTeD4sU6zJre19fzlAOwvbHaPs3ABYSTOs3nilkiQfRN2f+oFS5xr4dWcB6dsZ2alQ
rqavgoeHULKaYI3V7Zy85yp3SV/J60KhiH+zAS9OYSLfALpMERmj7bZ3vJ9TdBNblHHb0H5mWHw5
4U8FFkUYh5a3BMMxKzBf33+MGxMpK5/IwQjN8+138uy++cUZ/ovLgXO5QgjVlb+dG9mrJ3n8NOJP
oC8ZCVfeRlOQdDBd/2MkxUU6w95tcsrFbaBGkUt9CUR9+Bx6MSBAErD++OPRrx7jH5j7zrCmtMCE
0T+636TjlrrQAt5ayFee7GQBx9f8QcPPLd3fWq+gfQMWKLj/jp8viFpIdLXG/UJ+oLnB6KAcK9OZ
WRcyeyu08E3QvHMGTdhNpjVqtM288a9Xw1ofMwuq3KcYHJKTDzg4RZsTWs+lsQSZQ3tXct6pQIcC
ClA7A1ZFVmB9ICjNs36MdNu0hgYy29qWkGebdnc8edBJCUfA4DlKS4p83UuX7E92nb4hmBH/S6QY
oWtsekUyFD6/O1PoYv5FxILZ+o6EPWxX0lt+DUVKTwVXCo+KO6JV/wS7t71r/jvZVn0jZLUrelOs
v81ZgBxVQyyhgBxSSIKg0YNGy2VbF68X1p8y/AW+Ezcx8hZiU9/GuENERB6tg4LSDRIwCl1PaQS1
k1PAqWg+EdSP4AfQ3TlWXZpggFMJBlqv8tkjnvH3EA64v5b2SLFgmkq1UNw37/+uVy4XetC0DO7b
goFS4Qp86yqUsmWo9jrGQt4c6qgcu9UX/zWlV/rLuMld/ZEjfiuETHKjCwVefOuWDhgirAmDHLKU
pP71PkeA2MSqwIilmxfSX209ZJydpefGuYUDmx6p7SV6MlJrqrA2ZUAEByuqkq/tp+G5YZU4dbX0
ehwiaejzu74+2jhRCtkLgLdYI07chfrHQPJrGt5o12TgoGC5IZMURXrI8iQWNPPgBNJNTSHKTrMP
Yq8HcLobqXcCGk/3tqP9wAEggDuijN3/coIblCUl8XJvKTb9B1snzuUVuk021uVAOUskDU++NWSK
kd4TP/Wpq1i22pVPhp5m2YOa9dNnqElAPWQvApYTAMJiM69mw9S36jO71PCQfvTodpeL1eoaWEP0
BMApUQqikPcElHI3zEMAn5k4OxjL5kFxad8zELUT26/Kr3pJreeVtGhhXeFwWtKw4DQKj04++gPX
BsXD7VL+zVhLyGY62HtxEhqteosZ3wTa9xR109xvfIeSEAarifnsRh2sUn4Jg1QW2n5CdREkyAdG
DwFpJXcE42K5yVXBDIVUxI33BEBqoyJ4oND/OYrVcnx/KPg+S7xnOCG6t6GNpT+VBkwxTpGwyUtL
kId7CeJcPISRROsa4ej+4MdH2KqYKCckfd1Bmg/GlP53+VjX/GAl6tKV7CMwTgpUDNPvaPxcfQB6
kkZl3ABbaVu3eKYWqkadtJ7S4qstbxhKR9CU8krPT88HCZeW5ykw6mTzm2ym7H2r26Agpd+oHWjM
xUcUxAAepRd3gjwqPzxavwDgGj4I5hGLs90aAM0dZ7ZqZef4nGlnG4Zc4jUyfdHwQGnvMuttOXas
0SzRjdixMGkwKPsW0crQq7p6x6nCBmICaShdEXqQBUkxf87KvBKKEtq69sN3Tb+dKfaLJfs20iLN
GUNrtOo26EFk/FiSU2RvOeONGt72ZwzUT4zX4roI68C9eKFcK++sNmhzYTMWI2vdPhLedSgXPSoK
73u9f955UGTg/stKp4ksJgqdd9IoO6CnwPwwgMvY7ptlyMSbywotb6yZJ+mYP+sW2sFDBtNpSb1m
2JUPagtOBqFkg+6G/g9uScGVUGglI7qEeSWErO8aj6tr1wjavH4mdBM/RkHWfdWUoYrLqv3/dXtX
PHrQ2338Oc9+mCtUiAWAf9M0jtx2IjwTLw48gqikwmAOuolMBt6/POxfbFjt5IdQ86g6LzbEFi3G
cdJRwg1LYASjSJPX+LObIhaJNvO6y59oMbuY6HOcrp9RSn4g4BAUaWs4s0JdaBICkYRHwWxtBo4z
ACAAH6wN7KvyiEzj/1OMhOg+eyc+1yLkni3NcKewv5PrZgCQhGT2P+nKh+6F0DeHDDCiGRVuLzUE
eKEFguBwbY327tz9LD59jHlfR/f92mMrkODMr4Ag9xmCDfF/M0xqljZtU2Hmy3VBoSgDbXt72hUi
qdsS3aHHyyz0mxcVQuoylO219YIivq0mXJMDyt8uQRD43bQDfbngvET4ukdQtzo30tlUur0HsS+/
rgB/BLh3e6mZRqxRrbL8ywngOhETXtD8+wAhOdYCln/jUzOr5P4JFjFu7evrXxGtps5yclKa4HKk
2ZXNsShU/2OqhFhivQvaudlHKo3zaTYKosNq+GUQD1ekOvjwCD+G62vdZgTSRnrWydVrWZtOtWUo
0WIbntwOc+bEJma+GTtDm+Cnnws3xixrZR1mAMTvJ0gOcPeZ61Fri0Pf1tvZHycxfPZb11Yv0gy4
jgGOM7e52SyCgtg02uyUJe3eao0Jifm0GMpm5zSzIk6hVdiSFYRVnRz2gSzzE83OxxIl7onI0Hzn
63LM4jm0QC9DRsFyMmsGNrA2AqF9jmCgiF5zL3J0Tnh1vMG0RK6lW51aNI9Ozij2DNLuHoY1j99C
lOsub783ZEatOjcGfvn0PH99JKoMWuUHt4za7RhGhNZciki87LWHxlviDfbpA3BpyQP8fM4vaVvO
ifDADD8X+Eh1M72SKrvOpGw5HJOC8q18V5Lmv9Fc3Gi6Gkg4Svwu+tp0ldd8Oqym0qApIq6Clsfs
IC4cASr4lXQMSbwPXBlBoYsvXyrFdAdEclz5scUyKYGaBWVKuYISVf1um5XJDEuMonmLCZ8DWcMe
p9Xfln9I0+FbdNvP7+QQrl98XGq2x69uDBXcVayun2haWWq5g3Z1Uvk0uuu+78LFMnnyvP2HI07U
A2b3cRqXx1cbBZIBZ0a/J9DuEOivVZzpWt02STZha1d1VAZMqsJZCQz6B9ABOlBINdRyqWqQGbPB
CYBM2T4H5WiSy9Os2uQbrVnqis/qpM4Ny0wd0abO1JCS+lfgRD6Drif+XJJRcm2NaX4ZUq0aHGhR
1fAxsdXJN6wZ9iQ258Jwp4n/vQkxQglQ98RryzHHCdlB0MQGLmghXg074GPmzjue7/OOyodOcjyh
47t1Ork7TKkVUaBYiIjbZj0efGMJdqbWOkKjk2ZUQbpuIG4yMY2a9xdtyWHuOAOzYAL6zXF6PEye
XX5vZ6FEeWzQM8lIpRpGQ2A6Q3b/qdaC5ymAHIfQOKV8/Aph1NHp1RFDrRH42revE9fWl0IW2yGH
1aZFFkX60dYpSaRootZosCtZgfy99hps44TS1w2E2d9w9jpWkeDa8urRFPFBLpN/b9zGqvxYBdou
YDHC2qAzSuQhKsBpj+GA6VhDwmKfesJd+lXWoRfueedY0D7/YV4ZsvOprdbeLYxAuIBy54LbByCi
sbUUfv7SzSE8Vn6VvnVFEJeUSTbkgwr9J6BnA6eFUnw5FfYJ1RWFcQtfX0N5qTT8k4obgWXcxZEe
dXAMFznNzLeXlmRuqcHyQ6QR1A1MADImFeqiXynzg3poOAQslrJoX1EWwUwEe244jNyyFBlx8Krb
7Y4aaIH2uKZ9PRnOchGOgwSjC4xaGpAfjoSoU28ifrVhDoq4loExYTPTMDW3sMIjhaopUWPCwNnR
CiCbuQZEl1z8Y6mQCbPL3+hmXZQ+zwupbe7XFQ9VtxFyztMQIeTsSYf/T3ovBW9XM51qpDM75Gtr
ifQFGOmxBuDV3O/Zolap+ck4EhfaxC+KmOhVL7pz95etmO1/Ttjf9EwmCAiCnjCxlZ3Ssa7jCO8y
np5217Jk2Ko26AwYRORg/SYOa9X44YeDZ4iCHf14Uh++CS6NVy1DYliFrem+D898icfn+fu4HkJc
n9fATu99CTSMvyiwZVlPi0kwdeSWs76F7Ra0vzoZn4T/o0YwVUpIdxVoeWppOBmccd8y/m29zMNN
haHfO2YEaHxfPplBUCIMLOTYz0fiQN42s/PC0ydA7ZLyhZUEPmei4rK7rnkqDe7YOJ49vHLGBJOs
dTIUuGwrXZxkQSRf88aQ8yYzNTn9sAAF7AP0uUa8XqQy/j+dBN+jerPJ52XzzAUSGNDIYdUUooHf
veM+qKPV9CXRHDHkAerPH4F/W6igPTR12S7dQUQoq4w3g20iqJcGR++xp1Lz8Cdeot4W6ODShlZb
a8StIEwS1+JQv+3tK7ypI+iAP6Gr/GMQ2qciuCs6MYtBE1CmkEHe4eJqVzr+FCyO+bAPBqEpQ+vE
r36gd6f2PI4jmv7rGj8hzwltJFAbdxejYXadldD0wN1fraGpJPEaJ15UKfXlw53vRX86OMoPnAyH
dFFu19GzD2qHHBiF3nMe2KE+PktQ3zHPku9drewP6rBSMrI4Qmi+hhMcxRfIwhy9u+3dXhSJEgZI
l+0btHIT5lHOr/vOac8NWqIQ+voao/usDjFdnyV2EE5F+eg26VF7hUIv+PKZ3UopkSQPFn5wjHRO
s4uL5kxSfU/oPcyUdiuugbS2RFd+VS0hwi7Ln0NRIOj92dPDaDWhtKgHSsQ4o8eiKvTGcfrX51wy
aCRcNBqfIXy0bdnQMb2jTE41lDvhGjzstbq1LcXSYTSh36YCsYYS96zqbXkr00p0DGpQbzO3zd9A
l+52B5f2vbJqO8tjbnQD4iEDq86TgjW7gGv7kso2TDfoba0jYG1vYBodEDWxVUw1yQOhLNg7p/Rc
4gey1vPKnyhuBhF8HkMVeubf6svczEcU9r8/Z9LKvCPi1J8R9i8taqqn10c5KxwXJGUfGRonnhsk
rsbKw2xIXKW/CWD6R1/B/JFEGJ0i9CrhWWArCFBTSSnyb2+mtT/EXHDc77htCFqbE1p6Vt/Sg42G
IUYsHOVPK36oaD2xVWa55b6xt79aSq6ZGc4ZhFsWb92CMHL72nPCYgBOy/VPJSTLDzzq3iqnBXK7
kJxqzA+j1J+lnMxP6q0sueUoyCnN5hKu0Fkz2cUgy/8gPG63bClv3KabS3IFibwd94Lnvi7iNYG2
MQhdpW0CYbmwXtWOwy07pqAPRnMVFu1h24VIOZj5W0G9/1w29In8yZx2yuBOhEE8fmR8pNYtQfRw
SYYKbIqnKEH60eb+S1KdaBrZF5DtiuTao35+mRMIVwYCimaMh/wfq70Ynxkr+Lf+N0VvuV0SUpwq
qKs55kCy5yWQ45Jv0C68rh74W67bH8DDjaTcNgByLJj4svCToId5P5hm17eMkZL34chMPiyb5lwJ
c5e6qneY/UH7J+hn51qjUSL8TTpIals8VvSSw+ozujCrekHvtAhw+gKWYKGkQIsowv6hQJAy1Kua
qN60QNEB3P/5fHxbfZMDl+wSD950wYkZHxHBJQdyRuHFgzxqOm204z5gScQD9VHXJdNJehdQr1Q7
lXhtzemMiYQf8BCm2ksAUwI4Z6XvU6N78cVbPFvoQVUeztR8ZSuvWtqOplyKreTH94OZYfYvxj7y
5yR1XpbPRsnz5PK+yfbQV5V27g5x5gfh5OMHUTC97KICTr4VnsV6c8c4N18EDT6eBsxVOxm5XVQE
UHKT7dfEvWIBpyBxa+TuJfSSgCeTX1DVvfdl13Jf+d/9f6joyZXZgbNJsD9d6XCRmF+rbIQSjmZV
7WiXHwLoFmsXQ10hxPdHX3iPHfF8I3ANZiuEIxUhDXCXw7kjYaRxz/XoeUJ23JO0Tc688Lh7sFha
bVsL0A9ALQ5fZ4h7oSKI60M97pvP3tRDBRuZskIiLBHejFerrfBi0zf9yhxsnapvQ4v4iTevtBkw
VF7svAHncgmNiOBuLBzRpU7scaEz0M596hn4k303XedW8Ztuci9ryf70nbBsI+vMyRiwxo/Ti2va
NDWRhOnfOE9ueLRNxFJ2DIzc9apEKZXJLzWle3AWE6FlCZ9qYB0RqVmxDcW7qilhcXjlKRbkzPAQ
Et17KYpxKzHYjq/vyPrwkXKeiMQ5fddTSjS/7yV+LWfYdO7NBHq0h5HtLWNcBVJ1yACvLDeKs5NR
4t3qTKkGzU5s1nC4h1iBuuvVVB5YuwnRiKJ5UZ/f4suO1THXa1lr8Si2IbRe9l72hPjbHIyNa5bH
ySgLsvKnwQQsPlkPDFQRhUmlsv7OLPRqyvnAQ4TrarVyJlunyKUea990G29aUT5cE2baYz9Taw/Y
C8Wi23eOvm3HXfidrDAjk269YCXUiaObonrg8bJ4SGKe9jM4SOVlr7p2eN5ONmjMaQ1EfGEgIuv3
1CHZ+FpcU/fRQFRvj0c+0IH2UE8m6HzfvAQAkLNhNkWif7gPPLNUfpaC8CzzfjaJt+EHpL5L6VR5
qkWC1Lh8DsJMqT0XWhw3AvAKg4iKq1Sl+oTVDRwqKxaidEudkM4rxJwcOdZTmSQ6wJw8OX9dLcmK
ug//RgIkiEn9X4TgzzVw/HDOu3VAcCqbSVEPWgLFSlG5LdcN7jCKQSYeeier6NZ7vhlNQKkbZ+Dp
5ybD9QhqdHgitwdqR7ThrapUnU6xM75oU42TE59QdBzM01Nt1SEBEs/sehEQpoV/pVHWJuxwc3ZS
ofAWCNdj9yirnH00Sdf/GZliC6UXr0X8+ev0zEqg0onSefJqOF1nEKOwsM9wUUaG8v87hopRUcAj
ZqPH43j2MR0fRHgOb/t9hIabJ6qmq+oxV0rmSvnJvnYwykgoQe7omTFA7zk7flcq43hwoAtDKhzK
sh0vIureCzxnswRoTEfxYUQtqPaFqLZzX9hdGA7BLIpV11JLABePi/bd736AG4/jnINdxHpll7Cq
6qBB1SZS5t2wxBFk97ImsCjMUhJVHEf1JSSKyAWcHhxMLyegcEDlRjCx0mC11/2lHBg+o4sTl155
dPIp41QCFawbXPZo9ejx6u98SYE/rZ8pMTX853+lWMI7LAFnqhj1EGh+LPfHuLrEkUvBBPw2M26f
8VkbMTOpaS7VHCNV8wo4BM+b9MJV/D+mOc2EKoJgHjbe5+7R2DbzRpazTsr2ARnB6Ge1smWfQHrL
a9Dc+5kuxO5XqZsDxAsr2uFOWQ8poP7XhXoMRjNHrFl8hJ7QvHaYZxFCp7DPQ1A03r6tYJgsik4/
sUR0dCn2hqOk0ZGS+SWL6g34Su9xgMFFts8+SOQkmPTaLJH3htJdT52Ho6ESQnl8SyMyaVnZc7C1
yKGm78sXkQCJ4Bz28xujizSMFZ+vZtcS4D3xyBg7U+oAo/dYqO0co31XHFxUtXnqjCF5gN/BlCJ0
7yEIC41al2FLlRaV8+qPkmxMWuYPj/zY2SXRSjf+q/fHhOOebaizKEFBdXrf1JX1noIQ7VNL5nz0
LDso0Iwc1kStQJ1/UjCmHSx1kL/Ab69X9MlF4YZSnMTfbpdoaMgaHGUU7IQSoz/+DavgZOnrOE7H
UzkmqX8SKibTKP2pwB3ga/ruZuMPbN8eYGIOlP0oYtdqg9jCnRtatndo+5swg0wCrJK43pzGX9Ew
Oft8tEFOdowvf9zLKh9/LaKFjRX5WZXiKJC7LIjvy/6GeBvDdnDzSnptog6jZnVqJpb+4YnfVo8f
PA6ycHZzBd3BwIBIgcjkWyZuWSx81JgxT0ZujpKlKQGcrcxLibVf9NaPJi6fRpln0NNxMEth59CF
XJIDB6NApVWQipIGPzC2jWlTsK542jz/X23r1PbqZrvvhwgW+15YaMUmyGr/dlDdCtgklRG/ZLkM
egj4pSTs1sw8iJUFPTIesOmCFgEn6c+z7YGkAFKgMPcfgb1m5HO9o3ApDhKgLg56iRSp3zk8J9ct
ObK9/l6ozHpQC/jn17+DEud3E1hqzOT3+55I5ng40s+/020kpXFyQCCs4EJE0Rw42b/bzFia73kJ
0wqMzbrmHj6ImlvZXuXngt8usEI6NTyWQQGzcaq2Irv2X1mIAPSblgD7tFf6r6DeIuJv94omCpdD
BJ3odI+CnZtm4gqgyUhdLrD1m1oNhTJ+y5jbpa/YpXGn0II+GVtrsE2hzHiwSmbbICg/Qc5Sf7iW
5dWC8+3lY1LHuwKukmDdjFyJDJ7TlmUee/fQto72xx2+3p2TPjsVEIFmnrjSbCAR9gFsefgwM4v4
7cKm3a+TtlDzbS7olYZTwHebWf9Pby3J0SmDGlEg5uJHZ5UPgqMcY7gj7l05wKivNakdv0XJF01y
hp9vjNiIOrk64noZNYJUOSK0vXvrN4oTL0Lq4+yq/xbhzDTCUtmU9C97xuX+F51pFWKSmzpwvBdF
DbNyKZP11VS+glTHem63OssHhpQ74bvJIFf7CFqCBFqjF99JsDUQBAS889aM6IUbPpZzJE207pfO
uwaCNr7kAC5VgkmbQvdYjexGynXk7OlCPx44TjgUas/E0MYXAYB+V0iD4C8qt/sAGQOJ83yVHCXg
7xIsr828tyIxCdqW81hW18pYIuy0um1ZtkhDDhpj4DZPwA3MsYo4rY0eBnZHw66qkiNUvv9sUHKw
gGPz8tQKEJz57vP4kBrcKt42Finj2PxXIjyhkNMfQneVbf368hC4/Po4aZ4mKvoZWBGKZlJl9RxO
sdv2HET2u04RPE1zcQTJzoLc8uRNiBXJaGZIHJHIVL+T30p5ToDavJ07fuUujKMaIU5wllgm9b37
0lDTEsnmkjblmd2AJzoLbGRG/CSAZ+Y8S83J4ieo39w0kZ44TLPk++9C4Xu8XJGgSRmFaL4P+nK6
9qp95rmEYFAoq62+BS7fntyhIOoI5jZfFcwm9Issu0AMS9CIDii/itlJFxo2SWWiRLT3O6IVbnnP
05SgS3mUT9oUF7Lr6EipZ9Cx7CePjnEoOUEsrCrtG5Vq11yA117GH/EtTH54cYXhCgmxLhGmd2EL
Ih68R/o9yDz93BijaZTSbXZ+4F01FYBN6Im64uX78ScXzx4CMzYx02P6W9PrVtGJASBzcR6UJJZa
CIcK39fN9DSafkC5ETujCWKm50oxmpErQmBx5e9uJrOqucyPloih2LaaW036T+a0EE/4ZgodjlI5
wK66sX3pbRc2sXt63HlUaGEnwlBjlVfyiq2lHkoEuNp64NIJ1XyNLDqLgxOyZp19j+z1+KRuHjJ5
lapDU/iYIpQoqnFdpajWcZxBjTr1FxYXkuMavymj8IaKCCILUxCP0I3RntcbW+phpyweEqbTIMef
sddj73ujUwF5PVTRX2+cNC2erda5PrxRelSAh1k8bk7EOD7V0smLQxRgzncj+nr2zU6rkd5jtZBC
4zbFtx3DSpYfCucfpa20hCU65+ha0zK17N931/J6rY+z8dex2CDLf6UxnXqrZthhxNrB5G35UTt4
C7zri6I1/T8o8WHNTz/HZFE2LOYwt/sVriswOSotdRRqe/1yLvgQei6gdDxm9oR9kHZqCKvckTKF
HlgRzoZm5KTJg2gzSn4w50H5S4V00VQRMZ701tQK6JhU55GWWqe4JKy2sj0veody+CQkUIw4UEz+
tTO0NbjwoiWPztVrFTQcQdWxSyAgwNHbXV7h9fq9k7k3
`protect end_protected
