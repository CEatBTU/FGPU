`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZYOr92Gq9ECZuY70EjBXygq5nDSjp4+zC2Y5a6yqzQeRCO7H8anrBdU7aQydVRvTwhnQGwrIAFoF
2t2SQbzU+g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vs7yxitOXg5+ZTiyQ8kjvddK/VYkW4Fx6qEWlX3T+U6Ay5Ft1hXhf3YCJoRdSW8aE5PRV+viJiIy
0xh9b9JVnUpUZdS1FR5PcZZMz79HFTcmk6IqmtzVfEE73Wxgs7h/EKCrEmJdoWZaNmWoZPoQ3i/3
1+s5bh5+euQWJkDxi3w=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nipWPMb/eTjvLfd9KLpZt/DDW0G+xaO0DYUj6snF4DETt3xIJe3sWvSK50iOhD6Zim9XyhO0s1lH
350uEhcNoPHH8WwC+KvhBRm8tQBKKc5bfxVXS40AHIiWGcdYLrGMUagWCMvTGXVmm+VcyMUdiIZW
2kZoYQySogX8aw6Mc9U=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uXQ4V4PLJs2toPHv2Eo/G7oRjXjJU4P+Lm56f/50svghwMYFSxK4L9/M99VvmICMWMPzpXtSsGdh
6FGXh/iro71XVf/Ahk8U46Yu4/mJDO6gkd8miRf/PiKd/rwgHtMMLk26djT63Ki1OuU5o9NbKIlW
iL2aRlrg4qkSOAcfss0I4DaFQeoumBumdFHwm3zMRcO8JMjv0pHziQrRYsIj8bibO8eqBe50c8F1
H44px8Ap8c+WaNy3G94pRHlieAE2xV/FRXlTdcZAsPtLmQR1vWAjgqvQDd1mCYyfStEz8xO6eqqL
UEldaCdQM+8YVaY6HOgB+DvSN9ybub51zLgFdQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a6OGA02SNN4JWHn+1O3SGnaCrC4oN2/Qt7lfv5WRDWRk9JvBl4dwVuGewwIYXMLN2tJti5XgOk9c
6tfklhlESB1HljvSoE/y/DkztAx6YIcWU/J2dfk84bDbxcGRtkMwgAP6LVPOaUBZcHh5M2GR1kQO
NxYAsbzFejsgqUQMNqlO1sX6cmgkcGy4AcZ4vCVYhkzZWAIT3Q4sLhimiQyEl31piUyk0f/6kzY6
QaxtjGsWR8LlAhMXzTh8WWNb00A/DBh+bdE3gPvEPmeOP1uN7GuamFt2Tx73R94QZrb6D2d8vD28
i4bg25a+49CSqDTqUxZFRYXz+ht5YxdQLuQLoQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MiNuJqySr4DBk5dXHxJmrCfBEmcsuGTZxtlSKJJkcuq6Hptr6AoGog+m+AvfyodH1I3hD+pRuGEz
2Olohkd+VAQyhPpmAvfO/TxfZ1cMliE6zkxfzW/cQ18mLKpZ7AsM2HgpX0dGInBflcbe+3x7yiey
S/37YPw8Rfxbs9GXUJEp4yWvzAyt3H/KaUth4GQfjoR3c13v9J2bMg6RD1VS5twPb6sFAp5xvMtw
FvNyaxqXn41iwRq/OLx+/5TeXHVV+ESdAO9XJlFbaef3qGWWzGQAerTYySDcKcr8rw1qgg4mGLv8
VqA/5Na7fHxJO/XyUqRdNpWkUmdr40dkw48ALw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 122928)
`protect data_block
9TZ46BxVWUfdRYemo0VggghAYI1bY8CQW5OZ3cdsU9X5X4H1FVgJpewB6QWPbOKg2rVT9WU2AfrI
hIlTTdfKQipF4CdRTytnTQ6yxlIy82PVh464bFpQ0atBq2vtPyoPxOYfDNzJRoO+x1TMANHkDO3B
78snvyTxQPL3dL6bGZvMzBGe8iCqQzvFONJri/jDSIcCt78bMR2rqyhSAywjTvF6QAe5HAyubuKi
vn1zM1VoDVqMi7BalPDRsfXKolakFS8uqU70yjUBn/liDqhiq/ZDJCZLjo1i/Zx73AAT244f0qbK
9sKyY3ERoU5cLHgQoqORxjxt9NrhaUALqYtn87WI4mJFjpKDKmu7fljtwEkGvBITQ12OFijpSS1D
YdEU9YZfGjf2hT6CoUcevu4r7BT0aSF3fjrhO8b0vcEB1T5rQzXyKIbFzd9GZzWKOSrvx5cMVVzq
pvtRU056JueNZFFY5h93T1x7uw1jAMoDc0AIvcl30OkLVtUl15R6WSyEMQfc38Z6+pU1le0N7Vby
mKUgLyTlEBYfwHMW7IIrni8IYsT8uM2oZ1X9KCeiKkwTuIf0JQJE1da8maSKsSnwV5T0xj6QYGzX
FCK6Ip+rYlnbvN7oHRHbnWYoU3D4hQQI7MXoJmQN7BmE/4XyZDmjlYxUROAT4Z3Kq8FbRrcIhAl4
yZehpEBmXk3ktLUoWsQ/5OoyPttf6CqjG4ciDllGCbNihVYXMCAs8sjgqK3rBaaBQ9+X3bS49psr
VVOR8qNxwMdnrlLnZMa0aHxK4WoLcUHPIx59cDCE5168kUG8WMmimvSntpZsYRaFQyrRi4D43rHA
s5RDKyoNGN3b/KWWFrT8iH0pYU6OZRrJ32DdD7YKr7qTEY8dFIE0fhvVYk3xRsIbRR0RCLbH7ubq
z0xmyj61WCZq4eN71th9Tz9+az52hvcpdOab8IP+pu43JmJ17Adv7XsOH7nmA8moKADZJ0Mze7aO
OejXwEoQ2hEZCw+HPnsKcycyuamo3s31F7iy7X/32RVgj6SSslFWKDdsXR+o8XSpoPHjzAtRRgzo
RFgronLSEiYJ7G/oJ04qcjQR3gyRUfQEKf7PMZutlY1rBoOi6pkVHEfffIKPtq6Z5Jy/t1ozpmlj
g9ArhIDrk181u3iK/0Xz2kP6Z36HtPRz8ozqDIKbc4zWkYQBtaiS/z+Fg78Rc/VL4tzh+K6Xleb2
LV6iu09SsbYpePwybhfO+bB4bHXyCRIeSzvEtmcmdQmfztErCR550Uv0mytb8XbQE0GQ/2/SFPEF
Gitp74wepUI06mQoy9YL6Yyf0thJURIdpEr9AlennzDq0Y+vH3qkBb4jwgDMmJwPXs6obw8TZHBx
fCj7GehBMteS5GHqMaimCYb/2rr3OmgVGZhx6un9R/4h9ro1hat2GudJx7XrxHeM/luAfubAVtWK
xwu1GZgYz/rA3Rus1fgGyUs3X1nH3qtOaE/TnX286/kK8ESDlsxEtMSr9V+0JSO5q+cuvyyxr4cu
bFZof7LXRvJpApHfRvjl/g9r4gPuAeO00AFWJoS87S0i/jnVBxcyKAUTyaR/pO8cTYEo1MI6fAKN
intOZv+YTqh5K9b21lwXaPx/40tMsJuV/8Z/ZORKpAl8aAonmGBKo0gmHgAmwsBm1d6hC3YegP8k
SBPXgNgePcp+0XX2xQ+/MEydlnsql1AV2bDrRwYoTKIkGLFqkbEiNjO+33JmCiWBNWyqKBTBt5F1
RWKznWZOoiJtDQh3DpbSCW0VMZs2LEqq4vmS9C9atfn0kfPjUI04Seyn6D9kmO+Ng5NNWuMQrVyt
CgSjZsNjMzYHH0YjL33HxPZlt8UDWegzXLK3bs00UQnsas9m98N+i8UxCylKvWGWGr2l3lJ2tFQa
py/dw4xJtwIKhTkMbVNDFr8duCySXiEx8VCcMIH8ecHpKejAGF9Hxmo7euzwidIEVr8XETZBV73F
o85lJB3ye8XdQwLxgD8fZ0zxhkuR1Qe2kiZi8IgJ3BvGH5VTq8CnosNw9hZ2/RzeVVWvnMSt6ChV
BloBlfaK6RlpBZQKt4l3sSd3XwKLN30SwAZPnfQjlPv9cHGd11Op+EKZ7LszdJEeK9O62Ft19Crn
d+VcW1da1ChJv2d8T+zE+96tnrlYAZSoIbyqk6OpPRKR7rajV5I6uyrj99arKpdTFBDVd8+Jf1i1
yjcV+wzP+F+leoV/fe7bRpMLWcb+2SLEEQsrGc342lEesRzKBvgd/TPTMKHMRb3IaLqZ4ARjYAWz
qSxeaYEZEtKJxCXEJhmAeOPpwd/FVhzvSzVXeBb1rizChHgOUujLDQKb6mwgGgIVhkycr8ubwY45
TS0VasQLr4g9CjbCIOktssCEo2Gf4wIy7vSRTrHqrmPHkMxEvzyMB/JVS6xSfqdlfPKRAxSTh9lD
rShx+DeQVtx0Yw7ekUZxXVty+088p/pzlrWurum6RIvZ5JEIUaTvgXnM5eiHgCF7HTvbuZNuxDzm
fDCUo6Gymt8l01Da35xJ7fhxvQhNe0rY/C9zjDdhhuVUZoEZXtUhrr3IRKqJAwn6aWfcst7Av/zq
nrhEu8WGxInSjGYIQFs8qlym0SK3h9vbZsjsu7XKTUsP2r+0oEyuwiAVEhOPr8W3xGlNUj84Qb4g
p6dHy9RoyYF9StckBTF3iOQ+4v74p8FnOEhZCnYtTE0ztx97gKLTjvrFgCJBe4wB7TGr4tr5tkYB
iZJ835vDSkzK+pMCyJPRTHyoeufOZpduBOixEvGl5BJ9OwyMAzHG6fX2FXkqV3y6K1luYAHC+/tw
ORBTFN1WyjRFV9KIflVCsSw66xqR8Wn6rziy1Z6wYzdnTvuzJsFvE7UJaDQSYQl0AHNeeMT+DnTm
k8s28e01pSkzNae6rPT/yicD6VxWbp3NO6qp2ricoE2CQu7xd/RyA5dCbVTesIBEuPmIWP9UTiQb
4jTeYwK7Gfz4VpzaenPMCwBJIOI+P/WFLaXevhKx3WMGQjcsSZTEKr3pRaAMXGPWAm2w3VFZwRT1
zyf/wbqQMPXSxjDqHAFqtvhmTTxAqHESm/eTmme6gSjF5wXcBVuErDu3foyImpjrLKVX4aDjMl92
QeLXNmdCl7nC2gRvydzAgGF9DqAQMCqqQGHTQK9o8X4YqW5z8st5y8nqHKyaQItM0aNw015yQ1oN
5fb9L4c+QWZar3rsBwCpNlmHfh3P0Xtor2gxQzj/V5MIikoL8dIKvJYe+OiWV1igSnngF2+HABFD
lZgCI2HJxwDDQqbdAnJqq4daue2Haxa15C1bJ0Kg7N9vk/srFeTNKGlCrGx4Nb145iCmMuXZipvd
kOcdkR+FzhWV7+0tPYh1GhIy4yV1808hUS5UJf/B9uQd64y/zuQYLr7J3Od9gggV2fYQ6LTQVct6
qWR3KPL2TRsgwDbendEqwxBWru4iTfwjJwIy19Wrlrhug9tkj3tbLRI+pimqwD4mIpjEzEogBZrb
+3/n2+yruc7b8ML1QjChbgYDT+LcK821iyCrrlP6kYE5628yfxqbkondYi1rDfPihKw7bNAJxmCc
s6ElOxrMSmNu9BMUF1uXMNbrqyCud26cEDvNczNba3FtAibe+0VUQh72eBJm6aUjhWgycMnuIrTI
XKuldfjyzvT7pKF/QWTkI/p+Ny4ica/NFZUUT1E2GBtdZwBxswVAt+gouDFNHt8/aHFl31m1V/zv
EHmDduFaS8va1JUnDa87HN241W4g9gu4YESm4oIbf7v8yCN2AfL2jweegwGXB3lN/X9AyV+brEAK
tWlDFd0JapwiBVjXbiUurk2CQ2MdW+T1e7zRgTPbEkhIZHgOyrd9iE3Rq12TRqSMI4A/ugqCK8mZ
1mRiTB2jjRBIiGwkUO66sSdoenwGbi8+FDSy65h2F+/pI49atVKb4SFDu49tEj5f+8XSNi3tmWED
WhU68TxR9PyZEj5MwGJaVVHFrc/neigaVLFY/38+DpFi+/HZpeeLpjm3R5KjHqcewUSirDvfZBnW
+mcGep+nylJ3ak3Wvuyi6Oqfuj7+hDt/16Xlh08WhzYzjsvkEmh67dlzsfSC95f/6iP2y5rg2lPC
8TGPByzBASVRRDh16gT+2iZuzNkGDD3Ou+RGNVoM6/55aGrjvUCs6LAq+kXbotNwD1+oBeFvJVcG
1+sEH8KzEo/9o0E1hmvEBqsXbH9gwt1RuHNsJ/86pbwmQMBTtMz6Qa/KlwazsA6ZHusxZ9kYtcA8
ae1+Ch0xkVoBvnTMr1mRFacWKTxTpHOG+y7Vr7mFJA4WF7v6cu30xywYNurh4eJHvJ4g/Chmak+a
4Yw/f9b8+NDc8f+Y7SlELU6MlWA+0MivbJ4u55h9MhhkR4Ryz+YFmV69boTp0ZyZ/ywpGkuSeeWx
3IuL/ThZFQxmGub7QUl85BGS/MhGTNg4WfuLDBI/lzcJgpzqmTbVTRZhfPokzbUxr8YQsEeOq1OB
iRrWu4NnXhqRYQPLyIt41C8YXfGqHCksegiIXbPOj5YdhI1aRaOVGm47ehRlpwL/8Wh/tMhn+eps
ELG+G+b/pKW8ec5x05N8jxmcOmm0MUFZvdbKNQfHJ3r2bk03wtTc9L80w4QS5S2/+7T7cG2rX+L/
lIlEk3gllQJrixghXi86FysnoaLCIL4W9ZZhIUU7gecvY2KYlCTIUREdLzD2fAoHHlL6UnbX+l3S
9YT6WSrVa6ilxhtyQ6dbguNBkI9wGJVVVer+tl5zTQ0zUq5DQhv6moW3PuonPVmPtc5cqSCFBLvr
bwSUitzxG+7FFNL6ciBJow0R9KtCoF/fSjZ8tcn+g1beZxfI0pLwD8gAHnYkdFMNqWEg8gbTB4/C
TET9bDIT/v+tpOMt6mvrpdrYVMyg3l3OUsp8dYB4/RQIdc1jLe0PbeCXLPZ+572WyYC24HMCYQ0Z
C0wYVF7Miay4u/5P6g4xv0rYG2ZSo/ONXZKehKgzFf1ajMWa63VdajB4x9boG0zCibbX4qrmnekM
33ZcJsUzzi47IOBJeiLBgXk69gJhGZQHpt6TVZDaUpFRKZbKxHXhF+xZbRqAH1u6DVMhA6tyIDWv
S4V2rkiS44PzQl5Egf6Im9/O3EzXA9Ie6sCRQuxCXYq2l/SKxT9NIz9k7BB6/0rVxrG8guUgLobC
3YnjAhfXvpjVsHBeifCGA4Y45+0Y7yAn4Z6KjuEPaBMpsraQqJlq61//MRzK+aVJGyXTfyjlmS6B
ClEoJmWkCmoRfi2CrkGS0ScHexWbeNuSUkR7hQLq0gboMpVUJVKS7EwZsuKFdoFeuUbWqejQ5ZbD
hDBBVLujAbS/3aUf+x5Agg/d9mR3CMsgED6+o/wQhMINOAupDPTGqa6MG3R9pw+NEcDi+9L4gAH0
i9Oth8Ydylq6SEXciRgFvt4M+yBu7r/57CxCTdunTvQtXUV7iyEYplUOdEfMzs+835AflxGmBOGZ
dt6+2oYT2zxSbmWMCyml7ZdIlbkJGti+EVNVVgThn5fevU/6WTS+9HcJmfW5hsQiS+/s2LyLJY+D
iMSxXz35CW197OkRCpihhtQcL0tePwjd7MfmVjhcWGvUQfmEi9PH/aFPfKR4wkjcjMw3jLmcKVCY
NBk0euq2Rvpdxd3PLo8RFdAVSD7NMOTpgD9HsdcF0xr5xe3wncweWDFZxFOJnIcromWYKfVRI/Nd
s1QYv1UfHdOP0NvhufeDFQ/cVNdhGwHbXMhU7VCbOlIQf6gvRRkeG9JBm96AYz3ImrDauiiELvsn
Q2khuzP7+lA1tlmQ5GyDZ2UAkZFuQHEt5wrnGpSTRUEf2l6cPrX0DWbEata8nzSCO9aOcpi2l7uf
ZsMZQL4fRPNilpkcQ9Nnf3mQBwu/yjnvNv/wdLjCLeT8YYW9qZ6IveBn1DUxqJqROfJk+Do9O5h5
2kY0F3rbdGTMvfh5J2X0e6VROjh6ePG3FKGeczQI13LSTBKCKBsoxYynADPTv2qqkDMzjk6c+dBM
Z5pmBiwEWbbQt01agKh5FLupZkU9zhM5DVMUwLr7IkKOCpdycBRHht1lHe7mUxw0Jp8/Ooi9txIs
eSSf1jVrQJXqA9ecIHihusb6Vc9CfILILHIohkohWDNu28NkrOscY+ZPw5TmBaCCt5LH5K7w3GeB
HwCJf+lf/KN9uzgB8Xtytw9hDQOG/UbcT3zqPE06nD/DUACusvanptlVwyRxRDL0QSFhEVgvVZIS
oOoQuaUyuMsGy/m1e8fOQup7ds8Xjbkkc2eq4s7HawTg5YCXgl+Ea77GRQV+O5XOwtaW5CpINVQM
Qzjbt/uUmyr7YJAv0sixZX4Qo8apFXbRlv6C6f4UutRcZOejOuMCws1Cznrd8UXYAT9m+7/29yhG
JnrhpQRqxa/dv/LOdL+f5zlYwv6T/ShPgWxvyIvLNd0idqaNW0WQekaBItfqDv5nNOa+fyKO8FO5
SXD9oWwhOkE4seuGjWx/5+qQtkCEstRgvD3bWxmzgcaXCRUIRD7GLbDQUUQBxedyioHR8Q4uFaD8
EdJ0wiIWkpppFu+74wAyeAtuAI3poeLz1jsyAtC4EYdDYIDtqVTjIzh2YBafix7Dwl6jqNvtYgOM
CQkHY8QYUSvAjAJD6tfa+PbVEeQwhMc6Y11QcMq2k/V+h31B0mJFTnt1qivy9/ck6UF2A4WaHXH8
09e28UlKw7dOOt9E1R4TOVAnmiG2yojBZuS12vrqRxgN10xpAPWEh3yKr+HLmM8N/RwNDFX4JvUY
e0f5l0Cn8LzC7XoXtVck7HUqF7/+OxaPhnsl/ISHUsB7CoHr7qhkjMCpCvN4xwHYRXi8Zln/ogw4
55dBydlRjtJ+bNyiIHzdlJ/fa4JUjzI2WXHyH1ahydpScuqbFLlYY5xz2ActVN1QynOOdHlxZ8Yz
jx9AcPG4Xo3hphSY4e/hFJzjU8etSBfkycrYZiD+fS6AUbAMeT5vt70uqHeeBD/0uGnUASvOxcxt
KtWmzB/TcWkHKjyvwukhefme9W22/RGJMkFqPbIbZtwi9rjzYJ9J6NC/3WO5+nEzzZ4BCPFR6dMl
izFhFaH7mney+cWBFJcRR6cUlEYi+nAkF/v9Sc70opcL+DEUWKxiQykodm8V62RNlDUpaly3ajJp
kcDlOe6M8H3+apYY9rXdM9ci2gnGPRSC+I9BYMjRKGP5sfVjY9KdPqOY5PJLB0wb1qQ6aPh228mb
WB5x4465wylaqxQj6aYj1v3p2F5Ajvrl4JtjHYZspeWFTuemKNEZZMLJKoqAvC3kVFaQfRk7aTUO
XEYz4AzXK3/5bFCBUuSvkxnrI4C5xX+2Q67N9vYDBUSismK7SRzaA7OLcFhYoSnDWyVgRalqL5JX
V50MR3sRMSp4TM+P7RmlFyTJj5MikmLIiCA8bUM9mikN409gz8pd6iGYwpCQP4tacEx8Del+VZ6E
lPWxncFDKpZQZGamd4ytPQlG5ohv3znFMwduszQ8I3YuZF74x/PJSfg1BeZjEwBoGqGtKY7BFxDw
7ms1T79TCWL9/8O7KGEr9gr4z0AVUMfxmagK2/eRyyJQwNWzjuMZ2eohM2/k8ktc2B7u8VDuOUZm
zm6xYzyeEd82FF4QAVdmFGjz8WhDNQQbU3RSQF9X94EGwMNeosj21Gf6aENTptYTwf43uuoNc0BA
b1cxgGFG+p9ZpzY8m91esCE3YqLMztnPMQx3gYYYBicQrssEZ+9MP2cBdMOLhSvD2wPJpeZrvn2C
P3BHMjy80HsC2hTaMBWDEIL1/0fCkrhGNwNQ65/kVO3V5mK3aeOsLZqi4IkSo62ul2ePuJ8cp+we
UVv86PbOoW0VUuoVAvnyWlVYmbAb9i7M0dWS2Ovs9ftP2tDTUl09CBuoNcAaReHAY4kVtAVUy05q
a/NVwflXA5GHzIoklKgOU3IIk1iiO2xQGmZc+ipDnqKdx6vEcNGUfq32/jbRORR6HUlU3/D1kyjb
ikvbkzstJm0Q+38D7fZ+JpynTvM0+n0mMxt5yElnbFe66LCbkfDMYAbm68vCYj8RfIq4XwtBMtXo
SLoJPbU0PhKI46OLgllkvDNcBYEXIhXiUF+JSH+eFxMhkt3j/JcaNLV/rKrAqUgY/31zapmfTjSt
UomfXDPraU4ciwcqkfnf+RxgIeY6bG5IoK02Ljsm3WsjPTGJjtPVKtu99oAuPt4B//QB1T/w+dff
NPtE6iEzaLfyVam9B8nT4n4lm3hcS+Sbhs/S+cX/sQOeTv00hGx8iyq/ocZ1h93McReYiIQLYbRr
yHzbVOGoP8lNZKFXS94oSvDnqa1npa3ir0CKnwFzHRuPWL95pRkaZDwllI8S9Y2IUm322VZNfKJt
Q9B8gKIbk3ytljVwi7utElTrCOrba6RDmvTOrtwwdvYES4uTNQpg9RC3h/Srxcbomm9MbQtSNhFA
zM41+iTXDTtbRC0+m7FPDo0FPgPomH07ZFZBSHz7sUnuAC2aw3T3avYGGy5nj2uPwOtb7Ac3ZXtQ
TIhxWDwJjxJBxtqPl1D2JvsNWI6HUle77/BOQuXUCDCnf59S+lprayzeF8atx5yM2FSMkP00fDXu
hVA15flMz5+wuyaUqu9aqTS/V3UzrgskCq3iQ8/cklz4VtGr19jgY+QDeoZudC78vgSpEepmomzk
Jxi9VW0zq0YXam0IehtsZg0XmWG3lBRBDpl7WkBOJ4FCVyq6v1yUe/7oI4KhsEaRmMTgPIpY1rxe
wQDGurX4IaVSFmkHaUqA8OmCu9EpsoKGjEGB8WKh7vknHmXL6lEkE13/J0M5eUJjuoTVqLxEwWX6
1CL4LDipXs+uRweaayVgvD1IXZRudNl4pRm9W76D6dFwa5JcUw9MdKUWVnjcHIUFnxorASi9GG+q
ifDzDxWVOfDP0oNaWgQQzGiCk2QEOIw09wtWMglKyTFufE8gqEu5gkDZo3u+JdBz9XBQXDFYXb0n
fSfoyuCTBe1HKG6eotDOwI+rKMZXZudlcu6DiXYOuflSyHbYSIunCShOKglQEaaqUD/edPipi/H6
Tr/CSnBxRDslaEQ8z2oJgCjadkRdvEU3H6EpHmCgdefKUMB7xixHqUT6LYnVRLuN1gMFerltv7Gq
qPajEOvIRKnL1CGgxnD30l/ywR3twVsNNDfQrT/mEZg8vVeTmwaVwLoZzBuDSMWKy52c7Du0QT/2
vGjuLmuk/YhVa4PgW+eKrc5NOAtOh7IqPCaBeYn0YsfJPpCLF17TS5MyKwCcTvmgCc8JkQZPBq/t
uMLkrLJaHtbHiAe0P9b4NVXuXucYWg9ag1lc8Mk5RTlWqb/TZGm1g46hDbbf8BnfGPxn9xpnpUmO
7rCv1HdukVl8vSgF8goN4BLFmfGyRkuFsLrz1ly0HHtbHLG2ljWXo7V7kS+mRI+pum5jAtja7z8W
CDLP7mQX5uu7m5tCW2Eq734E4KsQ5NM8sG8NtF3yn5mkKLBQMldUett/dVCYR67dOxpe1s7wnuWM
IACZmRvipnWu/Ir539c/8BFvmioxh935OyUY5rE+WY7I27WdG3oWoU6cJmn/his0OUgdZAIRS7ys
mjN4pUoR/DLZnQMgGSpahMlTdrp0lCeQgBw7qBhMAulVOnJTK43D81cdhFjaXuom+P5bUUef0UIU
bnDIuyZbxeJMRY3nUa3OB2jQS25FHVcmDH9jA+ekRSfd1uXkD3949bCodx3rSHT851vLkVK+WhV6
qgUJ7YmWNVWEm9Ci4EfUa1J0cav0KhRt7hPdpGE0ErYEwSwXZWUZ8z0MKel3fQBrF/ItOu1TIZE/
o3Yn5QDOq3H+XAxwfpiVwjYM0npiDDa42Mwn1N/94uG3GGSTzwi8jXXy1XVTk6yjjLMbBbNyJ+kM
3VOfKGXLQsOggbCI2qiPF9T6uEP6jnODgPHCMGkCtXc7DdH83aGlU83aqs/vs1kNRROwWMozIosu
YeKOgwC5ZMkWvsPWY5mOilA6ZcBkFHcTjLxs0U7rtGXzsB0WVx/FsRM2cEzlyIxc8hbLlha4yq4M
ZNFyo7IX15s9iOjkYnsjVUsQVcapN0Ub26woT4FsmqvHUi8zDUxfOfoORhYm86oAp84SLjwbhSh5
sVR0Jg70t1I+h2fqSHw9buCi0DW/Ed+f2s94Z6qPgsylB7CrSyLDLl6wZWLWC4+tG1SOWfm045S8
VQnL0FKghQzOr7dMKpsFyMYcFLdsUw453ETXOmXt9EQhmgaM/syjUL9bHGtyTnX+B3Ao0TzBxsbP
0pMx3Bq9ekiBvKkveXcvzOUzHvYzjg1EcU0WZiUvTXv02OAAXAv++YHxHaK65lcnHpLFkbxj5pwT
zXu4IAmaQJGBvKG/A9Y3CPa8+fwRMu0b9puLqKQYtXeYOekthYilR5/M5zCK0rGUT5mem8W4mtaU
8g9YQtT1gg3K6usFshfjpqCI+Dd+BceNcmSocvPf29EkGRZtHa1JZtve4k53iZU4sroqmfeGEBqQ
8VPx4Cyjp7oZO/0j+G5P4+93YAApG/ms0qLEKvHUzi9AtNmReDiAZTQAkkG9XfaTXC0dSMUm7/lr
gVUGsCcXfMbnacwwzZsqjBcaou3CdC9bg2lTj1Zz9io5AbJTXLIS6wve3/X6OacG7o9l+EcYn+AX
NDW8zbGAtmq+j070SbVubg5/zQ/6xsOws3Zz1pHaTFwgxnoIZK8UfM+z2YCwlZSfaX0f32BqfmPp
sUr3uhIa5zFfk4+HkLJLKpFdHYukqul1weycp0RXTj2exuMniT+DXHHiNSHGM0TKG7nBDcz6uCZB
1vCiWb/N9CpsC+IzQ7i64YIA22iKDJH5YveYueZYWCHY7XEQWxS9ZvhbknzfYjVHEhJ4ecnSE+ik
xK6mAW92oV45WC7Myh20qluao30YSCE+gHH3FIq694gvJCJ5azObmUaMZYOVRwcXVAq408X5/ulE
YmkV9DkcocZv5uTVdFQ4lndKI03ZPTiBS7OKfWSm3S6hWhV8mIk4/3cr3goO8+A0er+A6UHd7BlG
Rq7zfe1ZKyemeEpAfqfv7fFZ031C6X95Dl/cbgKVfDcujM1HyanwwN7A1Qps3zO69eALAuWRyp1p
XXlnM645ZKrwcUTxnHyPThtiT7vGcQ0CHzg8YdCQpGbtKzy/wp3ClkhnzLeiKfS7S7wLg5I/WSlY
88P3V1Utf1YKdHxYclktIwvjvuBxI/3yvfC33aBgGbfiJfRG0b1tLqCTsJW+fUViF6J0ndCSWkx9
tcMVsca/oWqp+H5sxyVch3IKRpQGOrJSzAcYt/RppAVSbJB3tyYCxlixgZS1l8IwaZN4YJKNAyiw
ImPTQ+fi0sVQyA2v/l2XJoYjj5/H8cTSQv8rPTlJJynWBXhMi+HCe2SUu9jEmmxbRNVnqu+PwMQb
GYK4LvVQ+lXPVjbbYaL92SH5GFnkC9p/bm0zoI8tGjAq5veGNbscznPRAJAocPmjna4hnoPLTbEQ
lpOpTmd1lcXGXNOLH/Z8B8j4jimV2HcjV3CfAfMTktikhFYjp0IhW5KfPDWVJBsAkzZbm4or7tQY
buLiOkasJ5MH5yaox6tvibh5yJ42Nt7kcDbcwKAQywW0qyFECz9k49Ie4/D1arlkHf4zO5gC4oLg
erv4EA0De4f+LB1Xn1k6SFs1TSWQxQ3y/u/6KjkXKZzYzqKgJ1Xx6GIoxvtSpzX7DWK75+ugpLm/
Jt3Bi41WrBRXyxOLChl4yUOioRF9nOw0qCxW3eWGr5PH35kSXYae+3NqJqBH/O2Ehg0CeLrQsFBl
LV067JMEHpYstWBbWzS2hr19a2mg7DGhrttNOEzNQA3zVlQGrP3Mma34arzDB0G6nkf9aQzjlZp2
RS8OKmzj7iuvt4Nwe9h2kzE0PichoZP6TznBlN7E1uSyMVybOz0H+prWSyKN4fEGobkfonqo8NGQ
atsxrk9PMo4EBFKOLCeLavhgJvqgRNVxZNXHZ6qPoJIzoDTNJSCRdRB4Bo25Yy4q7h7yEaHJPjml
n6889QRj+v2rcTht5PnSsI5nYBDYLX85tfZ2b3RRoYiM0My0Ov7JIaoaY2WVvFx0UTy3lBDtuTUr
yZ3mLUuyMGT0J1hRMgNx5MFnMNyLMFex9jLKMAnTodXToKGrm2F8i/DBVYhavCG/Gb7oatJC0UUV
qXr2U2Kd0Ub13nBO8/QIyPNjpNN8XL8PEwFZA7lVwkuyKdJjvBsLiP9b2CwkrbibEMkAwb/eZtAr
0IiWWl4gnfZWi5UYdFzaD+3C3PpD3y6xgXSpjrived/B0voG1KxnPcqyjYj03hZZkbAk+zluw5O7
rQJXiB6RKBWo3y2j8QoH/lEFlgFEPPn+kU3C44kBhq659YeI6/LIegGyZd9N0TKDQdBswguXHppb
zz+t64cX6hKwaNA32wbkL2aU1kdZfIhpNsjUHN80VPcQbe438R1sev+9d7d0qklR+ewdoF/cDXzS
ArnxDIRCETNjzUwr33D/RqiNG2jadqt1/ZESpE4SAL3+WscApB5Co7vlp0mSbvO7UBDMONVoEnKR
W5lcZVshQWKiaIrGYqjktDOOFZRrBc9Vua5gSsR29LcKCp91RLLWNbY/nZX3IhpT/pPc5hdFRMuv
c4s2Qo6TOqLxgdewSHbcM21QuxqlwcDhZPyD7O0lavd/I08NqQHci5i/qLbBYxghDMMkDLO9mx9G
bnhyAO/YccVzLVrXaeplPYu6Rct4bdV0NM3ciednsHO7U3S4x5gmCiSbci0yv9l+8FwYLveNgw7d
DQ7xakvuxdimZh8iDD+qh+5UZo0rlv/58zo973PJ76STQNqd/euDRyzP4EfdosWC/Giv8j3iZLbV
naR3srJ14e3mDVfkmermy1ECrk0ipCctteIF/+Vk2DM97bUvzd2hGEKT0QZ0lAZygUA9oGs+I0NL
O+4pl3DFxlRpRJFjQdVteMZgY8OT2aXC6rGQabpXv0CskGXGR1PixZaIe+cDVp9FbHBxj6fwBPkU
Lb7ZPDGmzGK0xcim2floLYPglcBZxRXL2QwGpI7n+ZFztrQa5TaEtraOQwOZGWYi2AY0+tUWtx4r
SJOU1i3vWRJxok7IAtnfJGasN7eEXGcPj3zAx7hdd6e23EH3gnpb1cciz9uYmmyfcJ/bHkId0hKV
mJUcFm5QTrwpM6PUXuXh35yAiH+O4Mwri2Y6U0NxHNmj9yKhG4dVa9tSNDKyaYAbF8TmhHyBnMjo
hKo8uUGx3T4xqJ+fvioZFL0bzBmbamH02Y0u3UJgtbl5VC+6OYqSNddYo78IJw5eJSGEStZUTdx+
rJzx9RD1pHDWXRktNX/XDfG6menp3cXBNe/3YhbZuNnH/0nb/qP4jrI3k8MNXP3RHV5g025gFnkt
HMdUeP3i9Hinx6dezA5PHPy+lmFXBUCpmM/EgGBGuoEXnmXiMGEmZtOtjc0QcQohazm3/tKYK6KN
TK6bq1C+xtapRBq79T9U2H/1Tl6d1gUatjMbAoE0/v9he7RskPdA2ubBayRVbrHnzuKeZpxv4/yx
YgHQEmXhgGV9AKVPlI26TufhFGaZutWQoQstf2z3cBlGom5xEaNytnqFC87L68ij8GWf7T0rSKWG
g4b9f3GsGcGaOZrEoHnHd4TvCbI3+fHP79+1+CxK2ES8aYqiJq2xxlU1viMDZu6weuemRqi9FVP5
rH00zy59ZmiPy8nJ+2RJd04obldmKdrpJ4UBNGnTKL9YC6JGzwzDMQYfn+HTNuz98SFxq5vvVLen
5kxi9TBgVl/Twly0Q0CyvUD4aniPIUrTprzzWSjoDi5nbnrfoXh0qjPqo1GjBBhqggj8bEo5cO3T
6lHcqMpzvcwMG/6TzCkL1zpsHSvZHKSW0BEJWMqgnMB6tlK/58KPUkwCkhLVkFTJ813o4ntZ+X/u
BpU2IiDrp9bXoXnWU2Fe0JrA+L4zszBxcj4AVRQq6310qm71TUxJmQrcbHn5PSibg72wL1ost9XY
MqVJ78gO5n+UN+L2uTkdgQ8Llycb0l8PiQHEFTZnmj8SQxw3CRfpo1jp7GVsAwL+LhcqGQl3IPJ2
0THuT1e5L/6R7XKVAC/zmumKVNjTQtoV+TqMAUI4zIskFDszTX4tUChBqPkzCcp2IDAnub+hYUxP
JERh60daJcEK1gU7XFWuZ2c4vp2jv0lmvKREgHMLkkiY0s/VFhQaLz65KSp9bW9Fid3knh07V87k
oLpVG4Z4I1WIHuKQqHa8hz4H0MYLXNHJh5ZlHo9o3iZiCuVc3XkR5cEgn5Oh0PUCvNwNcdsMTpUD
AiN0SF7o7y5U3qGgJaexbjL6Yt4KMFWqwDAUXisu/T3QxEpv+LHao1vQOLK1zm5ylJchA+4kR6Kx
WIu5CFliWs7I3sQI8PNSfej/tMWq5QFq1a5t/BL+4oGPEYO/OYRY9wAMUzUdcKFvDIQNr4wKS0FJ
dlCB8xR0iSkQhNwslgwdAUr0VDa67XDronanKd+ENYmytvzZs3xRL2deVSXqp1Z/zKvoLsh/YGRi
oiKNvKiM1ty3CORxl2oZ5H2M7aAex4GJiJeZ9BadKuviV0/CcuLosTTe1rMhpcb3/ManMYD3NZoa
uMIYC5E42qrkPoUrDS/0WT/MdUnSzSA3yfqnoZvg6irhlGui2KKrK28F6VNxJCWw1EFWXRXf2MH+
8WlbTc8Fq+OWr2AlOTUXge1aQ240yS8MZOFn52IOp31psn9nIJ6rVExU5Ia8jT/TJc7RMaj4tZ4T
VZBftgouEgpNrEthgvlUjI4pnrE+rtnzDXgPYx0OCCaYbSBIPElmZ/a3DNf9ZTqrvBve9QCnxjCt
RttBipdNYoLoLx9qR1Ial3T0+3sDnGcFp4dN5BrV6EBtRSZSBB0VMdbWPXjNDW4fiJ7eP/uu6L/c
JApYvM0Iv9Icn4hitTBZTaeohN4ANOzWaeoOzPUJPMN39Gdtiru7sd/pZANsj2Zdixq8F2h4nVKg
xUwNaqFAGs9NnNfc0YPUa7D6NT64OypKzBoGEzYnaq/xBDA1hwjmPkpVsBJKbXykLZYCoimvOlfw
4UwufYyCis1smHH1PGk7DFaw3xpD2TPjY/nXhzF8mbB70JI97IHGbM8gTOVp88FJyR8DjmmvUZpf
au/J5zBY8YfwuRYzFDSvLD22HpQhWox6Zr1kopYIfiQQnSIUfoOF4Jrx5MhI1w3RlR+1zzinI6bf
DulmucjaXq6W3EbOvoeXO1jTSaAl/L7nRvMSSZcOTPYTKErb8bfr02Aw7QMNtVntbfObvaWCNiYq
4kIRPMOMZf+LZwn3VF/Qv3fXrV0jqLGyBmPj7V28fEFsLUDdjDAkclRH7GgPji6IeWfI7qM3SPpX
pex4OUHw5/5tLONy9l1KK1DCdsBsNFisw194jfS8XgFDQVpqr8YHzoQDmq98hfuqYqzNX8bAL9mx
nJgU9cDENnyBlHYiBqusiP6JTw1EhVss8YvkvEgACeuzHq3yYicHGY8Qg6e3kBvQcXl2f5OF3K4P
rdmd7cvsjo8a8taELOqF/VnRFCxHsZnyQlxLV79Od3vBS4Cxz8O3MG7TQSmrKLMN52eLOBy6oF/9
z4zfntfYyUEHmsN2fDFZOugDUK2mEn9jRkbxwWwgJAfHgwp9Br/41ut1eJnknJcRnzv226O4+v9J
U2OizSrDZhpLJz1JiF0zfkWAyRfVLys5DaCTx0tqk/CQMmIBGHyNI34Dly8gv2Uo4S7XSIuEFbvz
6Lf4NqfQ5iWDdSAQOZHWIhIVcMrrsrCu5RlrIyTDErmVuybzE+6xVPrvd2Uy/eSb8kkKY5IYETTV
kEHH+012g5fwGpssfMhrlS1YgAbNdKrhMj9ANV2XhOLY43DXWX5ipSUnpS7CAJnVLuUciY2XO2BF
hO1PSfWvSSH1GRPNUrjwXf7nNzDwQENQ90YvF8qxcmA4ar7C8KoL8/WufziR1eK9mc7vqdSnFmRy
r4JoDuNJs/tFEHNdKJar/BvpTrDdu3ZbNpT4Qzn+W6JmtJv6+AB2RpWJsGWNMZJ68dQTfXcAE7EE
L+JPYd1oBUI9Jd2jmqfvhZjA124CwWHU/zPHYOFYLP2UFdBxgLtDuDVRu+DKS3GXMQRiGrV+cEwn
+XB8P5BCOKhG+Wx13Lzt3xdjLWu+AK5ksz26WRxsZr3PZVAQIw4Sfm2m+lqIfL9udJIVzqEpyhxi
DUmgvLrcUW7bJ8zK74foNoBFNo3f5AziphOzir2YWxDOsCpEAQlkjCg+IvGS3+mWVg3mJAINlsK4
u5l7XRXVJqCcSOds1CZmV/lojid2B9EiNDfxK9+tuftHyi3DJQZ84sDrThICcOf7xbicV9CiOhrd
LtM65NLmRjRZIkjVrMqBZrgrTkLM3s/Qrigd9pcc1aJVluY1X/LrQrBF6pGF3qit4Qy/HjXpYUcm
KVxWt54zk70ztS2ysxkm7v3jnP9a7WaJ5MYFlBGDlgHWEM7h3u/kC5sXopFzbWVtWoCDsnwQAkHP
7j/4KZIOEaC3H6GYZxjyD0YWwydkpvp5kmAR5W66a+j2xAR8pQRI1BsQhH9gpjT1Pmg7gqOAHzOk
94sXiVMTbymi6hu8y/awvl/FFFahhCZkF2A2Gl7ei0gBb6L5qanzqMEM6q780xq29T1gPnA6w0EH
Rza86//NACV486o0mLEGdQqXnoAepefOEJwq5E6O19F4lsEUVRSv38fP9Xk5FYTgmzYGa+37XvLu
BYMh84+Ve20UFOBhWyJZhU+fr74pzCkLT964Trj+CzR7NxKdURs931Bb3CviggT7f8fXPLf6dxGD
DPnt5yqUiCFXS1DGw+ICJZw4Ig2Rerym/AQ5tfZF37FKvRwKRcb6hA/MuMvOq9rtf/RSzG/n/Xoo
EfMwFOPNTISzfiiqv84oUkfruaIyABoF6R73rRzpyaT6fLWyiY0wDFcWrW73Af9M+zzWgIec/FZv
zX48APcmogas5MvOgfWIQsHZI9ny4eBs2xpJBxehZ4uRGpOODhR2rn79GHX1tC250DcXDaeWMKZe
IHAMV9bMNHzaREwwkd2HaIQ6jsxFadI/f1aIcz3Ts4F206AjqAWSgnS9L1ko0sgtp29G/4m9hGr1
mblyroqmJCQOFun+Te8mzpJHfmO2WxIiQZN7CqJMCsh7VJFSG+0JND9cM8bgwJgb2LNw47H4YvQD
VNiuUB80PK+1lATh0LkRTWrdkNP7D1ZG3AmF+FttTlrpgk2gy5F/B3htMTFLIMQrSSFIJJdZpzNF
BwgqyR2rnLIsSjcPd0VPWj+FPM9L2uklOdgtc2WtOjN32g62g9YuqOAdtro2mdWZG80L4GUqz3hV
vUccS2LQwc0Bz5W1EQ7UFzxz+wg+w6SUhxDan8HMhgEsVydsjegS4RkKMwhKhjqFKtm5BJaR8TjA
zkK2dcRqkVIyYfa9PEiGHpJP/bRIj/o6jpgubWd29ZwId8CB+uecWx+m/MZncs2ohNNEiVGvRncs
/knt7qhYw+s4pTvMpiDG4NTYO2PIFypRLiXxnlopZ6asvyQmooczeb0kOZOXNhlmgPTKy09B6a/p
87S46CzYgkp9PJ5tkZyfxCh8qP+TzBlBjq3NaD+7pNlhj4sWdR9bvd4ZaYaEjSG8XMscgKCFrLjI
gXS3XpBo9a97JgRNQN9PE7u1DsDEYSybQcg7Yir4GhYSJB9zaQEO195iWcSCbaKU4/68GIC+Ytny
jxFnVe7ZxgUwzOfsGqDrJrBVzwxkN9NIazXLEHOlGEWx0Uchk3Yoo1SR5uwpb376NsgEmpDdJ+2l
7EBjs8DHykWUkksu6ipaDBJS1eWsZFjV2K+IXEzFTuDwORrmgXM0llrDzSX3EZL2X3MSXFUZqqMk
x2113+sYbLjraljALgLxR7P8WNgYzlA3NPG526nHgaErQVqe+RXN9NRuNGJxSYRDyUi+DWJoGdf7
bJiBw1f0UCdScYLdVdqyJnyBitoCoxRCexxSpIMb8hnkXP3QbgCnRSgndQbGnkrXE1FFOzXengLv
N0I0Q0D0VLGtyQ74JuiEezKS9ue3zOOyvV1P1C6q0lSPh8eBateq+VVOJPAE7q19rKn5Re2yuudj
PRwsw2fL08Yrcyfyr8SX3j2nUVilnmWGdwbrSQqfChVVkE7Kxmpo7CMx0K+hm1bXNkFzdBeseMCk
kU1ZxVmyHPFm3h2rTK/moC1gyShyiny1ajfl36uo/cb5HOmUtvowrQtR1i7Y72Vxvb+DPQvyVMZQ
5NTMHuf57bSwt7KZen+G4mmk/x9CaIVID3BfMgueDOjjG2toSbGayEC3+PTWG3IH59ZcBQ7oUpEz
xeqQJl6+3mU8VoDYFJoAzzXTr2KYZFJDVwCG/PWKu7LfUEZ5XI3sh26joHwGyI/QWSl6N2CNlFNh
LaRg2zfMuJsjonv2e21rkM8XrxlMyaLI5BeYIEsYN67dJRyPRuD52EY31Ct613hQ6IkyvrzSvHNy
anZLTmPsVPbcgIjTRGQFEAfpHTuUScex/HqNKu4Yp/kPqf3lnn50tg2B2BKGpaatKHsEdr0HJ1sn
DYba3IvE6FLjM9VvvTFk0atwHK9z2RaReYkToGtx2EZPBfKYYwEil2jiv17HMoAd+5thtKY4D3vl
3mBmCfCATJ1jB5ZYaMEsCDiVgq3vD0F4lPAJjuoj+H0M+uSWZtPJU/8eHLIHF8nEi5FSK3qW3hrw
rmObWog7zn1/Qxqw7Fj0PNISi5fQ8SFWfD+GfWKN1YEgEbFFFUhUdZDGhErKBPL6swkNLDt1gEzc
VZYlw2dy3+ho9fWT3KlDATayNYzivCH/eqtM4/uGpCX60v9rk5uIdj8A60cnitaEKtp5GoLpOXKO
hdTMbU8Y62qGhJ9v/KOKuPb3CUPrgx0CU3vn1Vl27QXD9dP6AZ0zkkM3q6yjm7AtHWXshpJupo0g
DvELRKM75rKkINBGw+2y6iAKJ+NdBqtm3qGB35YMGacmrQiAmd5kA5sVuIyRhHVG8rfzo3nAWaG7
EVUpZCbXeagZ9HvguAbMK1e1Lf0ExVYb5qIBiRiIqTED4fvvte2l25h9Xh/U4wXQW0Puj21xEAYU
DFSvPpgQxJoiqptVbHs22jYeG0ONTd+olJJFx4gDRjrHN91YfWA/a4fxuh6xXxJsaKHrCymKo8oe
ylN/BsBDb0PsgCJbtgxI16c7wtyL4n8WU3GN4QpU/O1MmL9HSOsz9vnDLgjzTFA+9aim+3/PnNfx
Z3l17O/wIAKFmuT3cnAPFw8c/EdeYdH6pBJImJhPgrXb26KeZRXr0W2//OOZ3Ew6rX2pr6xxs3a8
VVji8yMzwGjBKzs+OnLoq7qGq5iGGAC90FEoFCKqajw1XXGmeF4AbkLXy73svUC8eN/UvfSZcAiH
yRQoy+f+b5FtD49/M88btOYnmMAXbFxvk0uegALmujMk3vrNMLo4Nq2tny0P3MNSYk7fo3cotGBV
6CEffKy/JPPkRUEhpccMEpxzKpqjrdPcZQxwdx5nYtMBAlsI5Q2RwoHv/Yzqy8gPrZq8S+HDViQI
lewbdVk7BczEDswW7SGqs+42Ra38tZMKsF+Zf2fQPCWcRcvTfT9TLA6WjlWJbhWt+Xmo1qFGATG5
Ct7XOsUOqkLM6Z2nL/q4/eljZ1Vk5+SZkX09cj1yNuvKAGIsACg+Z6e0dwxo9bkAZt/NUqSTYJwS
rlCi8qGubbj0/PhsejaPZcQC3TIUtL4PlW6zUkddjx3WybmpduaDgJ9gILW/N2URxxn2e6sy59xd
VK57tIm1NufvvitQA0eA4K0Ab2v1JDsosiZ2q/1/CvM/7/REfL2qvqHI2I/48XNsIYUgPa+PpVK9
+7bEamMNp5WzLxanul0VJ+XqVAK87tDrqPDQU2cNYefGlHzZveHBE+IuM1D7UU/oXZHohA2vgAQL
0Kk//vthKHktwMSR6meRBGodILfHdFVzExh82fb1F2nga3l43+dV+VCqa5gfX930cyFWXDgAgB+p
bXVnW3dt4NmH/icXggzQVQnLY1f7y7PP55eXTYLublOdL8qH2cPNkHi0bchC7lYStkP6smZ62Yo+
LiAw9eiewBgB63PQjhkFsEhssIxW8bZrpGjfIK4OBh1rxXl707W8fTzl5fgVBARTcI2BeEtWNB4c
eCHjEioJfvejhNMfRxMbMsNU1/T3uf1EyJz7XEPo2swfA7WD6NioPFwzVN5Sw1UBJazGyMrcnqG3
4kuEFZOGPYyX8dmaRHof5mGyJJpVrR22Ym/LkxJRhHnnATMjVaDQlADihpoCSNlsSkooV0XZcmcT
7edc3fXgInTT6NAkUN5elbwWcsiYVQNg09wwVfcuengKU/rBWdCD1TaMucUBe3i0p2OwqTn3hOAO
CKtVBbRvMebguK+Cp0T5Xdowo2NjVb4lsXjiI+pavE0kpLpRbWuTjjjwlp446Qrinn3+01Xal0Xc
3kcjrEzdPZlOkGmyY06DJpftFxmCf7RGdQiIAKNz0ChwoBGL2quAW2NnxYHVYd2CEYxgmvBJwxBE
6o+gd1d3JztVMvXni223lTHGPIOqRIf3pNxy/dvCveDWEKL38e1LNjp62hTrBmpkgjcF6gj/0TZJ
vMDYQt4NIjH4LpE3pibW9476tUkpPw4XzrhG1uiAFNf3bCQ+tr7/ZMtpBj7pQY0sGcp8QPPuPTxW
LCLPMOYd1qgj1d02lhX8/bEBbDf9sOaHtqhVDKT2ol+bj8xa2mXui1fPk6eLd1b9bB2Euqvcp0tL
0l9itzxbEDedX+rTqcl9giesTC6oxzqcp44dMe4gkcPjUYKTp/zQIohMaCmGhB9m33BA1m/tRoKQ
+TP28o70+x1lZ7mAmpcjElzA9U/2eAZzNfKmBqdzCD41jsiRjErxmzDJTXQE3uo9ciiLHMGJSJfa
zmQ1Oa1/DGGC9VVvKZmLrj0nwihJ89CqV0ee3wYuCbpZPAWaiCGwsfwXM9Dl2DDDh+WSbE9JBEO+
9NFMLqauAJimsP4vgd9nw+y7vGLouKmpd67npXLIf3rhcdR6Pl6PsoQZGB672PWH0P38hi03J/jh
42fxPboykSaICZ8tjFNpeletr3DODYqOys4RLs7jYTCIzddza20FodtAqXUzObqvxevKs5d7ZihI
DrVq5vM/AnvthTYOFhriSwnqukFJX0uYjT7dcDZ9TvK12gXeCC7f6yiTkUy8ADry+pwFAB1RlPQ5
Zx6SpbXw09hlf4Qg9ILXkFJMm4mMMfOtm9o9USi7cBSYnQUYmx07w3SMK0KkvGn2nzYNGF4VgAdM
kZpRFtUspq9PoYon0xgiB/ZI4nJFO4n9dAMgiQVYDzKAhZxrEPD9YHxACkpYmSOVdmIwwfl4zVrw
N0URrZPRYqalG1CUCvaan0aWDgKoi7ZpZdBPFnFx3W+I4SWMI40DJWxqfpL61xBM7lgZjoyWSSSo
OMy/0bsYAIPEjsg2qhGAvvPkdpKm2d6FnpRcoJrtx3/yz1hO1Vos626qJ+85cRmR9hatquZoAW+9
ZaVU9iO3y0lIR9SNC5NOkWoQYqzBIEnMWCbqeKDcvsJW3w0HczmFJkp+so6RjOevfjS6Vr5JSke/
rBhNpNSaDSCHJs0ry1NOiXP9CWD5NINcTEPGyC88olHE5bCKkaL1N9mQP3Dc46YOQ1rSKVjVV+sD
kqtsTCIaKwcp0LSEglgsrHaxINLJEbqeBrdoLk0jI6mlKhojL+8g634iJ9ty6SQ3PN8bJsTAH5I4
6MA8i4iSQ2U2PwKdVZKAnGZVzazUGOMFYf3/lqxkARmm95WVLJBE83Ym8EBBJlsQGR0h3pIiIxh+
vgEvFiySD6IL3Ufvqfv4bIGP9PLOGSf2ydl95nPDWLxZHUabW7HNT7+c+oYs/jMG6t6eFSngbZLb
bp5FMBq7OUBwwUH3qliIAHDXpjZyhNxu3FWXrciTP4KZXFKViCTZSeEws3IdiLr4vJ+aI0J/rlus
dzU7BP7trmelYDAYwd28Aee+zZOb9tYTVXC2VRlgowAJRGVezkG+INKhpstcvchG6oFG2fmqT5cd
nuxiaK6II5b0j10aTJloKTOP6h66dvdXP4H7tD8Cn7CjEO4qbhXQO9/noX7DLh1/CfCkBWK4nRjL
lLcouaXM3Uyoa+knAG4RAY3GZtp6uG3sZvXG4rCfq022vxZOQ19NjKqxFEUB8c1H7OupT3RrThhU
s0UQD4RnE51zT3TrO/2bmYqUp3IhceeZABUKvEp0GttvOHEIbYrh0lxdPGsO4qCH+DL5K/OW20G2
hsLRK/7cuFHfd8nXM3mxjEaFR3ykWDEnb0mCF3CWVPKjkEv9rjgklVhFpTqdvo53hCJdmy0SdYZM
cfK4N2VzFvSwHrgQtQ1iv8baqwYYCwe2kgI0pFpvaGwJ0oFMNoTzUZQDXOlj/cUZlFhUXkpjKCSS
Ao+6Ut0F5+CmOLIFElzmME6SM0KdjfReHuNtljWG3bPF3FNnZimr2hXKvLNwKCET3TyLyq3TrDs8
cfFUbBYthsG7MmR2Q+NF4NRDd+WJTplYCcvQ3lBjvuX2C5UHY6BeCIBgHXq0sD2RPyhVFt1tr1pv
QFYIbnKZXM1taecKfZcgbJp0K7trGoD05/m1ExSnUj1hv9SyybOwKdURUXlE+DSsAxZSfnp2m8dC
uadVtaellXuI0pmekauBNUcFfGjWtFCLQjnTYPpPL422C3jBLu4gwIvUvl8Vsk9+PfIQXr1M9B/p
T3jVO+LDjJf5J/Sc/72pog8uL8BipGbDs+8hbz5X37p/NlCccUYXFprCG9/U+hxxQolV9xue5p0j
t0/QN6x/XLwsR6FOj7EsKd4M2pklaIj/FyClBKpvbBoRrEhqC5AVxLF4DAvw+OR7oqz0Xjqjv12D
1Lip9jids0LdNxTFaSqv2EhedNucVVd9T5nzB/MmuWP7Xf/JKe3w6pAtuaUyS28apgoOP5YZtwbo
i70cKWog9HyrJgQSfesGX04uNtFN6eaCRYZwogpIMzQ+KLuHJgY8WYzHSruOD5NppOciM3ar5iZD
Su6bBGupCsQ3dNkz2w32q/nBNXBt9RWGSkvKPwekC89tgXWgk8B0rlJNQHWAmCAMzIbvdQE3b9YA
+TsU31sv81BIL05ODXnuVoO/baP9+gORpl3VuTblEdbee4QbgddQFGT4Fe9JpGIogirqLBFlwDRO
YioWw9SiGGxD9FkDtqzhch18/XUbVWLDJ3KlBqhHpKN1xIN8sMgZ4SCdV6EOp3zN/EXNrKBznhLP
IYP1D1on1eRl7PFXAnFElyCAAv3G8CR7bc8kwqQrh2aMYt+bFJXRJhF1974SwRGjhnSNS9DFoEsP
9bEBjvsJI0iowYLjnOfCxW9bRvHsWlsXjrR83nj78QdUKFwSdutamdYZRTY1cYI4F/K5i6tL9R/u
eu4xoT+1H9iY0Gu0489iZGPPHXYyULjcan1hRgc53kTw7DVT5DvpIpzIGuNnw0Ha+3+/8G3BMSKa
TaMQZ414o5c+HMBBwe2HYMgnnjrdoiQ6hYRq3BQ810ZfvK0NH+q87fl0lziwcwbyiASrxwvK2p86
6aNGbstrOD3yiqwpem0KKwWgfMEIoNRuvuXKnWJzNKAZAf4yq0Y4fud/bNeqwS04OKu+xwS910E1
4SfsBwa5VF4vMA0A0oFRxEfoIEtKw9EKbTnnzWsHze/FsukA7O1hrDjOidgf7NLXVfzwqwBRtfXY
XkoWEwXdB+b6/3QF0EROZC3HEbufqYvcxX8h/Cgk5NAZa9Ap9TuOuv4ElqXY4/Gamb19thypvsb/
FbMawNGgr1h5ZAz7EJojnEMaIfNbS0laDKAFoGX6fKDqZ6qpSxWSvY37GgDKQn3ZH9+RxDbyOypx
y/nmlGbj7e0YYV9FijJjgrVo/ARyqz/QN4eXnzIiMp6cgxTLzZkJmI24COdh9LIVSoz3uyoSTX6K
oslAL52J375756j5QsL0JepnFCyM7zBNg0wTcImmZWZTyN7ues2V1CkRxctt3wyAnD7deWoqMNhN
RvryS07zqVEPi+Sa1ymJ97r2dx8zs6xnuSXcP3zWChzOpSBm15DkemRGCKJWJ37OyUGQXJtZT9/Y
bA7ytw3g5WMVIhMBbotIkSFcgjlFXrn/V6yH92gtI+EjPXGs8cyJ0F3GFYZ+9ISWWg2qqFDps6Ma
bslAFsbWRHH7HS22VtshAomXEQKXwb3QY935v69OJiFi2y8wODOt4761oEStKIBFaY40c24uypag
TNb9K1RnDEMlbgnA5Os06gg7VXpLiSY6gm7kz3N7G6oAZaNwi/zMupSKaoIzyUxn9hW49GGZYO9t
/ovlzQy6K8q03znqADaFUZMRjoLaAjEnyaDqz0h5Lrx7RNHbGxj16ob90e2FKHsoKAsP+2bGxkZp
4yYE5jJifj4K+Q4ApctH789mspcJ84i8orcFlDNUd0vKz5cVLR+d55fR6MgiBp/7vqqUa0I6wXPY
ZS2yiquzz0CW27w9spvbneofzTnrPTLCGUqm1KwG6Cc3eoftTKlhv31TQ76ysI4XtAMgfMj7CE7W
EdSGqWJ9l3fyYtduKiXbsDRWaLS5vndVgSuzknbuMltwSjI7RHeMB9etuIoh8SJI8D2qDZq/WFsN
wE8RuwF+1fWtPi1ci0H7cIbGb5cwHG34Wa3nbcWJfFcfNbCNSJ9rep1OvC5ihyxf2IDmlS0qudrn
Lhy2JigbVb6XU+EkoIfy8KfXuO2izw6FtBzaNSYieJzVOA1QGg9idGt6Geku2H8bpRXoXBS29GBP
qur4sydPt+oeKILGiLfR37cbaGQlGhJvef3OXrv++TKJhWEOfPgUPs6w8P4pZH0T0MfqZKSaPQq0
feZN894JfJikr9A1XsbHRX0GKQj/Fx6LLjWUEOQeyK/6rLD4AANL8pXmquHRHpPEFIQcHgzNkQfo
zD1mcauDJyN/eM35OJjS+8jD86je3M+91hLLPMEBJDNUB8EOOhmASWb88Z93LDiaPCuBTMNQMCa6
FvPiNMOIGIEHw89KyoSN/8MR1uhpwQGcqOJKAIvKZo08m8m5LP9L9a7cHK9GhNFEj7vY3sgiyq3w
VSXwbZ+CzZzK7dHEwI8+1RcXH5ELbGD2aCEv968eVNzDGbCqMrTVVo7h0Msjdm2MrPhCZ6BnQLJu
uD/eMpoV+AnT1oZVQpMZEj11WQ2grtoejEt71Q8wWziUEiv1vigk5Sr3kj9YLq4wOhHXxSVSdi+E
dbMfAhKSNqWdmwbxpV/i2ZeYkVK8HOM1JJbEoFFLS6BifBAvnDRdfPy2mbUlcRW8KVzz667UEMST
i2rVbK9mX2muCTR2iajzNLEtfd2R/GXN+FSuD/KWeDmvScslnFxI6MsA8+sartkJx5qMR54Y4xhi
4vGJA7sb90VNZIpS1Am2NPmxo+tHe1CYNPD5DtBpjXuloydX2oapoJ2tKBuGEh/uHTq1+YnWCI4n
kipKHQfNScVhbl94wxMigHWlKTERtPhMDxZg+/lAf6d+xDabLnfOJcruJTU5+U1/tNFTfC11TQ5/
BWj0rc/EqWad1J8LipsyiMK8otHMxiNFnRowoOvKkyknivhkhBZ1Ud+8V8xuTb8PP060AfY2BAkQ
ZD6MTqhvjFAfN4x5rv5HnNLkafC+CK7MXSnGSODfZ2Xva0JUURFOY9jN5JF/cADM/jQeuKtSa1wQ
hpHh3opbw9/ABKeMnkbJXZTF4IJ/ohaLWyp7Cekra7H8IaU+kqXuwLA6IQGSY2OYKQjGKTLWz+Ts
fAUgKDMvTh5riEBF88OTayLg8sbX7pXUUERNOc6QZ6SRQqQctbcBQcQwvqBABWICkHkygui7AM/3
em4GI+SoUGButmGJT+xPxnEfc+NAIhqepgJ057cDBxJDSuYD5lD+05cOCD8gz2AKUgLIKXOsz9J1
q76rBffdMc2YkuAk6+vSP56C2hQ5MB6f4xNnvy8n2avgoRVd5CI3ECODVIAOrNM3tJYgRitLwNOF
BihvaumHF3MDv80g9waKlHzRA6hIxcySyenKVsndh3aw+OmZhAceCTQPM8hCDKJ725X7FW8uuSE6
Uw1wDv5ZldLPeWp9DTUSumchIFeJcnd7wc1HPmV/MRPtRGLWKHp9kJ2EbR7yT+/N3E75ha57G60Q
Ty53blvxQMqbBuQK/wZmyErH86rtCgGRGcYGyQBuYR0O95FoCw4HM+3EZx1+vu5JCk6XPrDMpWc7
hO29ovHlX47WZn0w4Jdh54rnl5BBP8Bqk0j6pPL67DR3W4TuhSUbYIs9p6FCYeE58ZI2a7wKGOe+
9Ku4hbia4YSXRYcLWVzOR4+4ROIgOUzpDnP0zTB9QE9k9/VfjV5SDSIKa76ZMM1C4wIboyvdWcGD
w/RbuCGaFIOvvY5V+rBQbiib17oLQz/r5iQ7NcQ3vzWM3sFcmirgrlKA0EoH94OmrQRwI1tyVEFr
aEj0vAzhgpNAhNErHxvNaG8pgdA/Xlgq4APImI46CY2BPorW0fTbp2KFPTkibOjBB/ICZaLVJzU1
O7ekWOLwvWyhuv+36rcy7ANEznYeVlxO6IAop/WIw9wQgm3TumTz5VlLH/jZIELAL/NTuu0D9dBK
UZ9awlKBIuqt6+aTZxde9oCshWmqkT1vTMZF9DkMPSQ59vKlBV2ftn1J3Tq5L3aGF4CiUMFLfC1j
yLA01hi/u2TlbC5thB/aO5GedfsvyUUIcmYv1JLPhGw+5mZ7MlkS/yDiiR3W4r428qw+AeRYsycS
k+VDdd6nbVC1NJyB55nJSHDNdrHUalAtiDosQ/U9L3YV1oQCPkbESXeZqzkBFj5nhJ/bvblB01Jq
sk4H/6BCbVmtn2G7D50yzfkDRBtJiWD/8aHKTYhelRX94ZS8XH4ONK7mK2rXjlog9oirVozG2+O0
Mnpsr2Sn1JysafpPrqAuAIw6LsvUG4wRbkLqzEJz2AlE8pXz6BmEQfu6KVAgwpMd7k8JRIl7IQql
vXTFk8GkIA4r+WPQ3di9V25/XzDtwkbMY7+AhYpjN42iRZZ4mpgu1XLdo6h0UkFf05JmUhsvwlTE
3IxZZZDxEBpnX2kM+WpLWiYU0ghcaoiu8tpwx1xiQ/p8MvT0ylVsbaG942uMOWPW7v5uOTS92Jfq
aks2JidUWqBA2zk4NzM9Qj62a0HfMx8O6Sbp5K5wDjqxk9OuJXGjVvdLqAaqOS+kFQABOSohgi+y
ytdCv1nDyFhNwCjQyWJa9AqYc14ZFeTT2RXmQRiXVzl8B1qt8DZ3pjDJzO7/klx0VKITKGhbCqqw
HgywOEdBhwggWuWuqDro6nEkTXoKwsFZ4WCl5BbaC1m8HkRWBoCJPN3Md+ofSJy0/fTzYEYiv00H
xvCHhVfDgY0VMm1sIgV8h/6NrxdX0FQVa9dQ8/26DJ6urK511W460dArFv9C4hbrnBKZkIPjWKr3
EaLpLJ104rOOr7GfMON3eOQ4LiPMQCQHkf+KfgfvtuNQrzl4FN3Tpw01YiS77Dz+yRugS00XHuWh
l9mW9Q7XPDDLS4aab2Q6Ccbxp9Yc2T9YsoZXO9L34yE6oawqbAhlAhnqgp2WODm6NVemwOgqGP70
paT5hjSUWnQj4RJDOUNVVH6YHDgL39tKqRWoTUwHXgvFB0MQD5r3yZjKKJMU41Yt4JShQ5/006Mu
El+Nd5P6t+eOdZKJRm3usHAP5Gf1GY+PKuRxq7lWR9ZoqGxtxY/smndpXWIsbTJpzYGEramSsJ5y
BSxOb9MMTtSX4AmE7gbh3qr/pG9hQELx0qAFhSicVP/CvcOGHpoMdYq1Ty7mbLXPytJneupr7Fkg
BmEh8gT03TWQ7iFQNfQHY9+SFKQyXzJj4bOfCFZPe75IzUJXb8m5uGxzxoyMlWO4gWYxrKVySdX9
DV7/E41KOI/kL8ApCckW7ztYuYaZcly6qoUqZz3zV2eKTyemkUXXzuZM3fec/exvjmWK9uvANxWi
goXaGqpDRGcqnSNVeFLSRllTeO7ryq3Bq+jvOg6WJznkBSqp1GfXnXQmYx6mhlqyA9QIoTU9CC6N
+butKcSR9hTrFxReOV26XCSrUVPUvuwzWs00wShCx+Ny7Uhimonsdi8+VbmFJBKJQXpOkgNRTqLP
rnPkmbeGusMzk2g2SiYGnANqL1D0HOOiWosexDiktLl/+ixsistBcP8y8IkDAw9WIbWotQKPtRhR
AY0c+tFV4G2poZR6fRmIjc+Gglznic9BVdrFwch1oS1iodl1wlbP7poCNm0TZaNnH26Ei89zvT6+
/qpSVRP2kOxUvoA6atZA1yGaLuCRM0QqiVzBWUtrJQ9xvEUtaXb6Ij2azuCh387DA2/7UUtXdnOL
Y4qNgfoWqQpu8JjTSWT3NgNzVxi6gVHdxkiHeQXA/OaK7GIPCondozRVJInF0IwLiMjtDUUFUU2n
55SB5EqHLIJU6HsC/FHU55LYtCqHkANWG8LK1FnG6iR2yv8SOATK1o5ScPD1A+czOpWfR4DL8fNY
5Gbp0lnt5b0GcCw1ZLyJszsT/Aa7RpkMzLp1RTPDYsqW8xuHtKIbSn9hAQTf1ZVK3pUCPxyKy95l
pnVyW0iXqCxIa2K1Dcixv09wcGv4C9zUXtDv5En8rDhPiLIa1uEW5NP44Ro/ceHZoAT/Mh+50+TG
rgvkGXXhWCQGqunFYZeXF6XNixSRabo53K2WsmKLnWRn2OyojQ7e/x0utYeVNbwM42XSwITjWL+w
M24edjbn0PT590OMxhCgsZMFCHEQF2Tcv+hZGyrYlMGkIL3P38in3PIk/HlgD0dr3MNrz54zE1I/
ZQkOE+m4o5x+NktvD3Y7yknRAZiHE/ipgio8pPdp08WCEIJcB49hh3PLCK2OXCyUOilTjDjz63kw
jmOkwfij7sXIKjPfpGClk5qCfhaZNF0swAfv1OIQfLked4WxBq/DehPHE8yH9y+w3Av4JXpLM+Ai
Hbs2+XZGVLjMw6tL0Y41wOdSdCkHbxiJd9kLksNfoZrJhC5z4hGPXUoqy/5oJgzJab769RcwJE8w
oPtry6dV5TXsT6mUTi1vgSRdi6RfPeHEhodl6c2o0qYDGnp6g1SiLi3awqANXc3BnGaQbI8i+CbK
1IJhtEsgGdt6uqqKgv7xHDQvxhFW2XBX+WMgKee/M2u9Wax4AiZTMCXwszK+ewetYA5olJO/VbBx
zGk412jqvWMsr1d4t9hvwLpK15bcrSjg+DqvmLCzKX3o+eozOFKBaJuyUocIEkCqysfU3/vlebUu
ZvIzLG742cFptS1AG/oBzMUfZnPgYgVqYSQiqQZMjlV91pWYs0NxRHlLOH5G4Hfcivg7kcJIql62
LEIzJ0MCwdO8OVI3mu2wY5J3+7QzyVFoqcsKUR0PLIx4kwQi6hu26AvUBq9M+bHRcGhwDtuOONUc
LpNOX+4Bic91wSqD200g9HjPu/DDenevfCmHHfZd5DZDYVi9HeYFVirgfqoei0Tm4pY25EDJgjEH
Kys1JVAwtYJu+zcPNzWSKp25iXk8TjM44PYImoA/eqsOWjtSsQdloIyMc+9OUIrwgdFrln2DYosL
O55hoI/+0hNs/3elix8bOLuPh7YHLWZjYtqreUuXk/CiUKC0BmuoPhKKKG45mysANfQDQ99y51Es
54o8ieMsxZenYvRC0+Y6SK+RHKlkXcu2Gkjm18Dsfmok8TXQcGRk5Z1uLxevqHGAoM5WXLCOoVHQ
qWiuBAVSZ+Sb+MKChmWFCn3/tlpVUAmbip365qAzAgnpauvj51FEMh4Xp3u4pl4Gi/RIqgJNCmVH
vLb+sJD5b5I/qiBVAMNYqN/vjjO2BLqjIlKxbtQC4Wjz9UYai2wv/3U2CXzXF2QT1xqabiBjXcrz
UdJ6xrwt9p3oZ/hSRFfiXZiGPo8nwWD0qUEu4G3YJ/kKN/ZCttXe8tUyx/mGIzqXXVN2kJiYI8W1
MY7CouLFN3WsPPAyoJkfLsnfskRcVjqKL75dgS+bx8fjVPlNsXOOl2OO6LCyCvqjQSM5olRS6+5G
BE8y+B3ayjDyEEvKly0olBL/BeOZlXrLz7ZNqM0g1Q2p0wNRW/pk53luaO+JMfNmNGtsevQLm086
ymmzTw8QF2MowF1/GS1jkPjwAlNnX3bwzs4LRwGUEGVYqKRim8O/CDJlgjJR577+BQ3QdnAe3SC7
yDHvRElqP1hX5xpMFsWpkcyGGkq8v68k+C2zS2wgGFeVH6Q0A+oT5of+kyCjApfLCIj00YZdJrKr
tuZywY2znpzfd9GCDVTRD4Z6eQCNgYAfvO4GYZWbCNcFpUj7uSPyzRentjmZwfQTxEzdWufBTZtZ
IZPqrkF5ENFrfWnAsplyhEwHaMSjoPwWHKes9SCYg3yZaisntdwWUFvMqj5n63fH4fJncmqrhGLJ
0dWlNmU+7VdHO2KX4dRBCj6049nc/WzmbbU2KgRGRZARlJ4XHZvlHWwlRa6/Ew96MmdfkOFLGrVo
V9GLzLY8WUwqPwf3a9N8oLwU3Eli3k2Gd8Vu/m9xvK/OzW97s3pNpQr4UErMBflQlOnVfYGclGB6
3VG3BUY24l4mPWgIlZmMgsLY9zCOBmbi88vnJlNOKH8evCkGrCdp4Wo3He03xK/yPVjPBv7YceKt
GV68dTcBRsbcr+3i6ZScIF7Pysp6bZL4Wny+wN5LDphvjhGYBrFIVMCtpxDPxdZ0Wqz5a+aODaPb
k23hczkQfNSq0/UyUaEKVOdWrYqAMqhU6E9NUldh2Q5ynRbMhh67dg74PKTtHtYb2fDgNUPcSfwP
WlEz28fd6pwHqvpyes1I9BpmNpd07SxnbOIB21F0LY1NEv8xVtxTF9pLJLNLymH9v7phxMTnF7ny
iOxMYT1c4ZeQ4kcqJ/9qKS0pjuKhOdJy9TGoyLZZtt3tYvCDQF+Jl5YYOHou2ynN+v8WWGhtYJGQ
0UlowM7i4+EUibQXpsvm/YH55Hw9IbTU0wXkbxNNfP+yYmfOwumRXczrN4My6LloZiwsgr/a3pcg
us3YXmi2N0IAzMEZO17VkOHylR5t36PkjzNT+vHRn2MoQFo9OOQZ6jndv4Gb00JGR4bzsGXgF5Py
p/qryQ3LF8gm8FTnkG+L6Ws8UxowHZGrDpUbLiAdihD5e81Um6daELpBAT5tzbjm0q/Y/kUF+gUQ
MH6AWz8zdVINMsj3dfBbaoPjUkyeUloQBBdz3Nl41ltCHpLDmwk/EWBlGpd1pIj1H6OG2aU0iB6E
Bizxi7j7+GfVvg+nDEY6ZGCxOGEwJOsiDhbcyhONV1lDlj+r2CoSZqP2uSF/kIDBLCPJKonc3C2N
vD7Dd4J5hot1hG8OQG2HIOJctSKLQVERnvhxURMvnzuB0FuGAUbhJChWJiZlsbUBeLuBvSytXySF
vtL1sfUdPh6NEpLCMjZrhFSoYIDnsfY+rO+nm9zFNADbhnbFh4/tZAn3XnA+lEKyj9en6pV4UGYb
OyshToKAIsaroU34MEecB+guwUpyY3ms16AgJhZKzd9KcKH0zx+6QvVBYPOULFO1pnmHy25ik4zb
2NwWpW9TTO5RydVWDbRtqElNBTfomhdqGivXO+lAvw0YDcICebm4ESyNeP7snhOrA3DyfpQYUxfE
eOVx7AGMyCfM08L/CjbT3kb01m3R0fcjQwWmxgX5FitlW/Lg1ocwxRruD9OSoUbywXa/7FIrntz7
AYWZyNahvRHNDsn9dQApaOosiO8EUMYQLxH8j9UcYpSfG0rsAIQYGfN/xaBJjEwc5UwDf+U8mYIo
vLy1BRmUn0xdcuvkYRNm7Gm5Q1fSDsFBmrcfnUw/U9evqJvO+js9q+Hf8QDQ1MTrr9di8nnhgmMV
osAN2jhS/lgsqhMLOr6PWlNklP7EhMzF5mTGfg7eHEUgy1pEucrkx+3uSX694eEE++P6+eZgxM9j
qBvBj81NBdMGbnKapxx6zxg99uj2/Re1/VmG+CuGfmnNfv4UQIgNfLAdMWi7yIfAzq6GdzAOWhfC
fD4URJW7jtMbnoGKQ1qb7e959oiTbmh9MKHcxVDgC61He/yNGUYf/R1odTk3yZ4dDEVep1r75y8A
CK6gNcfnFLZKhl8bYjT8HfU7wMKu98Fb3JINZY89x5FujBrMLbz3jUhK9VkQWoQbXOwU31iJ35Vf
FIbn9aWCEyrnCKxqS/xF6tBVDic8nXlg2t9NsqSJK2mj242MMrA4qc/dw/PkciVZfNOt/8hfSqbP
X08FVxjc1t2nVLz9QpbLliNA5RkeBGEfSp+qUbuC+XLHXnVxHH2NDPEAScXKcfPwYnjcywkrsvt7
3WjJfAg9sJkAVE3B99bWoQxtKBCI3ZdjpDcFPxOHOBiZD+tHm4W+sOudX1j6gGQrF1lAzzrtzJQ/
Yre1SnMnaiTmKZyOoaBxxskJuyxGmwg7Zb9CY/wxnjnuzdnuKE6vXtLF9nmnTMn5jqMHYBydE5xe
CzZKr9JXlDKpiW5dexePpl8AswEXGBzWISsvSwAzXAaqHJVj1eGRZAiEFVIfBuZB1eX9PwzuPyBJ
y3QeVoWgXRNZxTsDgi15/xynFICIRjpS0GW5OplKSQy+nrNFZ/Q9/K4vCcAr0bJRqOIkC72HReCH
DK0esJNHx4fqKjMphEY2Fzvq1SRHkgdAuiY7LgU+kkOPUiiRVkyrK7yaEWO6N9ene3DWa5bXlkgt
gQ4nekXpJjrySawR89L/bywbjnf4ycL0VK6DUgf4eekNCv4IvN3bfOITmCUjXE2jVzqv9QpXxnYm
sTyC5CPhhC0qqZ3pKusi0W3cdGaay0YHAAw2tlKfws4tfuJumTY03DpeLIuU03EPjFHRxdMebkJy
pqVlq/crkNRcRggCjKb41Bfw6bIaKaD8FrNem0rQwRDFinejVatxu6ASt2zE3vU22/qwvhKnvSoH
nHNvKLOXU0CT0hatMppCPqnkba8ZoU7lyok4zYUl3Z9czxPmx3FFyWq6uymnyes7VFJFQ60D31d9
MOd/ZGUATIATyEoS1ku/ltqrEvjlSobIvqCTkfw0Fbeay3K43CpjXCenK2L5TbB7ZJ2Ri44oIYND
n8SB29mhKS4Tc6f5+8wsGs7CS8P74BArFSvH6jqf3VQnjCRwGc/2wjSYJCcAfh9ksWrUJyE+Iewi
usRb5YK5/Oekt37u8E5QddrwVjpfds+V0KFwWe+mlUG/Me6SxaMblPDofD8SnjlrbcJEmYCGFB4X
F1XWCakmenyZywj9HPsLygxmpTVlNNPw73GcwrHVu0+jw2qN049QPbLeM/60pHPvWliiaqkS4QYk
Q62gGN/fAI/Sx2ftFNx4glnNUccAjcesX036jBz0bgK7Xn/HNJtkD+j5M8xem8FDL5h88fpfjgnu
Oprz0fSrzmwNpa2HIpPkAXgQwbt2ydRXg6ZXNaX8wlXAdezTqDiRGRi5intYBvEb/PkUOmHV7Skd
jlnJqu3Ou+muRLwTGihMNMxw0fcj84Oyxmk/D/DPZrBRipxLcP/0HsEYE8WXwSJhoTbwzgYvSDHG
DNGU2zivbRyg8h5CSLNUfQddDr0mmIyJEMaMwVvXdyvG3aSMweRWxwCf7nL8o7+Gq2c5+qI4sOKE
9uIpILwc/SAH1hQxL3Yy7ccgxcifZU5GkZoyRfazAUCT4mAPSBU/5WsTuZUFq0w3KtLYuQJD3DQ4
HXi9PoIsaTYBDIakXXlwuT8SYPj3D4nopL7uSU4+peniO8ViENf1EnJ2E9VR9bB2PMUZo3e33qqs
uWWwgZ2AGh1ool2xyQ662CwR2nr8VcNV6S4fchn1AlF0Y4aYHeaA+ezWWXhnnCauUFczyyJeLyHF
qeuaTcplyBnUa5Wl7iHX0ZYXWhN5Qki2wfOZfFGvPDhzq0c+VTu6yVqlQQhCQ+HZUcHV+DXgf3VG
V9fByWtRmH1Fae8KPTYrYcP/BoEIXqcXcJzzSMc8blqTnYnndhS5bAAkLB6jEy4LSWqt7WE7nGwT
xSNf29HsPeTINs9aqYIpSkwaLXR+ZPjtTUiLyMxwf7IUHc2pMolR4c3yoZU/4T6SP/VbhHkiueQj
w8YJcVEbHwx+oR93CI80mYhkGXGHGzlQLsILWTO0+6iB7WbAloww4LBXec6euimR4hC2x+KMbcS/
P0OQRuxkwd2fGZrTzPSlh/bsXvw15zLU5ca+YNWueDebljqMIVMDCqfZCiKLICWMwQN+9YzL4TJ/
2xFQ+iPaHtMRBcYtXd26xQOLsWL5S0PyF5QSwlOqMOCbDWDsTUimPzcKHJsDY5Ce7MYHDc0RaJqD
bKWAnsQdun9rl4LkgCxxbN/2qZQW9AXCTOO4ZQJrG7TF+GmP8t7TPaG2WX4iK9say3Q2s+5SF1kt
GAVVInicWmwFcG2e3P1g7qLWUSRJ+L8H00AWT8xbGO++Iy8iu8bhv121yFw2kOzGFuIOHOox7uo4
j59dYfMktOI9OMBcNmDa4Nmu7H5lLeqnBlBb65yRqMI551FO1cTbcdfUhoNJxI6ZzwZTkcgQ0xjx
UghYfAoEeNxWmvRgZAfZmHDJ5kijp1Hq5wByNg/Sk7sT6yiGyJc4CfYwRE+FqCw1Ikti1v/VM0o7
rCXk+xxdw0HGOo/ba5enfCWiimaomewM8zT2nH1WcCmnOrEJ632XLo2b10aGHI4z3Ieee3oeRmtP
MiK9oaCprqBOeycI3i7PvNUyB6p8uEMIKgw9fM9SHT1RuEpG5JUPwFjcsZv3ABjW8JV68x28Jesc
NfTlxd0DAYaIZRF35iqBPTcr35mwkD1rf2qqviFrNsT2u+KRdIlnqwO/cQFbp6sP8ZMea6lUV2St
w4gTZV63UL6wsBvycSfAK6ygkQ3VJYBTdeUmhHaipzvA2gIHGNwVngz2kMfH2UOfsJB19PZx6il2
DSzUZyI7lBUQ4TYwpqZB3VVRmPbJj7VBoKCksvA59Tsure45wATmIgv102EXWA2T7V4bVVKcyo4Z
y0uDpzb2g0s1sJQmug+H6HLkvZxMLWvQee2scWC0B9xt1QNcUPPw/+OkTdhdRvHiCctKri7oZ4wB
2cmgQh3iTs4zXmDIuBNaPt67dslDVG0u6YRyMSnPzAzhqkne9i6GqASL1qiyN5usYMJwwMcS4pNk
b+TncXmCXxVgzaKnW3dBL/xf0FFUnoKugvAbm4QOGir39wVVRGUwtF6V/nh1ieWAdytX/i4Vl3v9
g+wydVYu9t7kmZpi3MP/eN3IFTi9YL0LxKMwOBGdd8N7uVJZPu9Fok+rN9pbt9n21t5xOJ3v1Uyt
g549s5H/4ePS6k6WMQgs/Pto0rvg3a3bt0TDOLRP+Bq/RqnOpStjfJ062/4ADOmpKge8UxLFlcJS
BYeEPjv45ernv4csM8HXZGKA4yCrcNPBPaaBBDVlcYI7fYQArK4fFIzTlF/iEmP4igCBwTYXrXxw
8sYWyH8JPGCMo/UQxEaMgTcrMmPvsERGk5VjPOAcXbzk1lx17DtZA7HEnLyZGQTY1JbtEuz9FMBg
wgW+jv+wX59J2zG6a1RJ8k0bpYxO8+2eL4H9curP0o4jl1OyCgvOZTJq+blbEOCvKHL28B5SIobZ
vCJmnmIYea+eM1afo8a1XP71CYSmTAneLuvKAsG4yeauDikEzjvd5VKYaBgsoyxCMAmLPKrakdMo
moOYvT6ae1prrcVEfE/RLsMSrYXgzpOF78HzAculHPXOonCKoUm+5A9uZvC7vurkbr8nGIEXQnv8
wuanmxFDwR5EZQYmjGpP9zkURooV5WP3nbSVIrXfBXuq/tg9EJi7LVROV1eLyNc5ADJtaFrh8dOU
zEoE07Y3yVbrdJB7/qw/tain8BICw1nSt2EctyWowwnUWn793VEkW5o2bRcPpZSefdC4Xpmj1JA4
1fWsfoKczjl5t6vNj8r7QADgI49hnUaqsgpPHD2a/Zbf73dctLNz0sR+VdFvqXLe9bNRnFfPRzgK
/FsdymgaBOLYTOr29ZTMuL/LGhC/500OEJOmyfryyFHDbgh6QPNK5yzJOydZGAkXmF2mqR8dHDeg
T8q5NAYiZGiwu2lMsdYTIG71gPgk8oesDSheWEDkRicCk2DnjrGOdYLNU1UKI53owAw/2W7FTz7c
xmp37qWneSb+WQ7w16dTS0kcuNrs2cRl77UZxx2J+f9kAgyfo0s19TYYvAZwT9F7UBohWhcEbeCr
5e5LDgnAUUjAJVhtk7kUuCy4dIq656ma9+ptJg3Ios2NCtmHaay3ScWJQ28aOk3UFSZc6CoVKcT7
NVGrzPmFjU3ktrZQ6hY+L0FKe7z+EQKG16c885ihM0UIou2W65jCS1cOz9Cp4ZWOTWVFmiT/sKFQ
wmAMzJ6vlyfC9zdu15s70PSrACo9ieWuHIHHP2WfuFwOiG25L2cCSWQhiwmPQAGNIZ0WVDnlUwnH
rjBxxUkZ8TroBpFgVUqzu2lsp0dh5y5O0a0BcZk4254Vf8HdaR/LUl6VtmyGbwU61b2jg3BVkvOU
KUz4wP9LO3C1EdXo0ThKoWYdBb6aPgJJ1iAk5Mav3XWFy3sdkgBcrOWHJQlqy/YebBzt7RTjYFGL
jgp/nroFhLwLZO7RSZk9rSbTGTWSKb0bgZzOrRHu/8YhT0RbW4nqhlvZ/Cgdc1uskmcObS99PrXC
t9bG84jJZy8VzbAmggpbpUirXCK3dusQfnh64OwldlIE2HnokjZzTFWN9CkJizZ/QKTxk9LPfxzd
XyYyoHjIa4ehchgCqWUWnptVddw7HIQrT7bRpNxXVGDi7OiHiPpFU2bR2k3NEJFZjPzkAa8VjsLD
pG4se5ZYhkdURFIBCfZK/VFRUgd6vLrxENSgQ6HPd/fcQzja2UwLBLmMeA1CcMyBmJTyi0U9k4QH
jYC7eB2pWhGbWUpAGnNWY2hOWhiVPnZ2dsvxLhCoK7BBDbwrRrju7TqVOrsP7mrs/inO+CzFbahP
1yqoA51ri3pmu45lfwD9ys3+5MM0j4r/b1NCivL6ulqCccz2o2hoyRlvSR84LHdAfMsqfeYM3Zrn
OcGknsABeVDKr+X1FVTwTuzpWb3fmXte+CHPBV8zC8SyRmGsqt5cBKyk+T01E8bJcdaxN/tbmoo8
CgzqRbOili/KqVsoaaB6Y/KA+dcxVsKE2RU482UBndI4uIxV5ZE2cTcenxVaeb416zTRNV+CgWn2
DYaW17NICOgVP1QGUnR63jI+F/0loRZA/rCWwScreJhmxbAvqQA/7tU3ABTaHBBJAGgDW/SOXkxF
koQ2763MiggbnRBmmAaRiHJ+PbvS/5+rvTYBEo3u44d2y+JvabhfNHOW9ThWeiCWqFPlhXumlwXK
0EJsM/DmXxPb1tK3JPoqfQciJvT6dFA4jtW/QAgr71bdVPd5hc08cla3NXLqZXZrTpthxFS5UubM
G34/8jG/374vzOTGoWngc9iruWzyW387gGmOBtMXe9rhbkfyFSGRmolO5xm0mUMgYVZv1NNXSxHt
O7PVxIU++ZlNGalDQnEZ6bmnochpsarozzTkcDADZ6ZMnwMsH57zWYyKse0lb95/LdXXVOth0C7p
h7XbUB9ZOroVKJkum/YyQE9oW3VOii/ujetbHW9oOWPl5InUkQGPmD/oBGi1DSWyxEuCZt/43d63
r7aP7LqM65nqSLHmVQ54aRehS5B97B0NGf2pfMx+UyK/RL8WsZgCVYulwmpYRCw82geJEz8jdrIX
J7Zwfu4NfEsNRDTlXWDbtQ0C/J9i2HYiR0AL1hbj4OqfrHyM7od2CYDsLCuJptH657/ekuWzizCL
Z27jE6oUFM9x21qC/AZ5snAi1CM3ifg3Q6SRMkPA5Ed2GVE9FZ0Tj1EOOD1slxiJUoEiamKdoQSE
9X6xtSl5eHszIFPNOE9csk4luA+1F4+kXxn/lU58dJYk8TMesxa3uDQA4k33qkz4/aHzTJJnJpgU
bk6id3BvoeWSDpouO0WaMmIaMpZ7jsm/awY1lBtUBMUTvUbaLiXCpgUkizbMQ9+jROvjSKQm9S29
dUt1umQo7mUpBiFqLp0a8fKZNvlnVqWiZNRnA++sSy7atCdpYAqmGO3I9cenqaKI3cDVHpOckjpT
qeBCrfYriB/dJlQptEKs/X+kAeGzCzfyCMRWM67lmxTQh57PZwHG/jMVNPYvocuUItnMRswaIOIC
n4+Ql3Axz38/HV4dM4uL2CFLxTvHji2WsB3qePt3kn4sFg/TTkvfL+eQnBjDIfNd0DWCDFsvxy0T
6SsytVfE/LJr/Dv2a+GzwQBUImsQuvHeJsZshOF5srsUDPzVThBEfHEBtpd7O1oiwo5xHF+kmmij
9fJo14X8fEKkXUyGaQuWj4uQgr/EEjqqImUH8jaJ8BP9IkyO4F0qXQFK8n10ghe5/QXq34wgAjp9
wWdsodog5o22VTWusdYSJu2RMaqZywGvcvRcgN8g54G7/gt7ooLMP4Kqtbx7R4j7cuatiBrQi45N
nJP+h6iUZk7Fmec9QWKSvl8j3Ul9x9a2yl5CAQylnbuCQaEI4R5Bcml+TzdjoRVNkCck55Cpp3GX
E6ubK4s2j81cxJmgFSS2LNXNLBp1clU+RvbZGGlmHmcipdVS+JwLPwssIcXyZc0go6NrmRncfqzx
0MXGHxOFyl0bSoIKAALI9vr2lb2aEKz1+rpAdYUimcHGZI4CwE/jYRm8ZfwYnAvrCvmdwQk3hAG+
D7kobtejSpYoCnN3OSl6K4VI0E3kjqQsSqAlKlRHm+R6aA0H/WlxuPDViaijxAKw78qHguhBjUmb
5BR+nF9Ix7VNNoW14CLCf13y0X/3ktgfg8M1+IHrTZgAI3x8xtZNkG9Fta0VVcUAZbq0jsdUM9Er
vMbbEEb/go8mI9/hItIrIY8bopxQW8F+bVHYcWPoGPosEWUo9HTiSZAlXKS7P8kmkX/CrAiFmTJp
4CYHH5p1ellfYswghDP0YOH0zR3Y6ZQq/ZK/tajSvpQlq9pOG2mBUm75PINiDxsmZjqBgxmIMD0o
AcF4sZb+Agzi/34iDBfXIlN2N+QFFAqXhgIZi3kmtXm+8MNwOp81Ti/Lw7rS0flc7+pfSaPDBr/9
gK4ULCfjPfeEsIfsMnGY02Gw4Uzr4Ia6KdmMllmN5LLSticOJnqvSpTkYbJnqRsDkAKtRhT7aQOw
prtxyrii+p14AlQYA9btUzeJHbpnTbUjAoXrJjMQj7XAQli6cdckyH2KeMlzx7s8x9JZ7drmUTw2
2JVSrotzn4khzHk7Li71ak5WQ1E5cOCvlpQikRqa1Qg08Yf1wL14OpeXsZZ78LT9lxzJtfMazmJz
y8TX3LOU4MJzUYgeZjDkaNiBc/C1grm+eDFa9yglgnihsmgUQycR1OMqRmBDcx8ps0hEltdDLc8e
5C6WsQt+IyBcp4ljkA29gmue1gYnVWLMn3dkV7NtB1S1xXeNx2toM6ouUSl2ZR/xB0p3IBqjdga8
8svJN7D3YGplYgFuo6jDwgaF1H9v0R/bwgoWwCpNohNt6au//62iYYVnNEzpN2uoIZmFmIktt2Dl
aVSZq3kRYPlZNr7rZGpBXCP4phrspbvdIJzQhL8bd6wBtkGmzGqfSBQsQ3LkhELtCfS+HGvy9fNT
5o4AXO2B4odkf3b47LbIq98WgFJUGNboyqTlQkpo9xTsQxDesXuSeaMiVPkT5IY7/POq4VyAxITb
IPluiJ4zaJX0f3s6AEnLySgzrelvBTqB8FzgHbnRdyA7kmi7MRNVKY/x93S5xKYBPClJWIWfnHIG
7pgryCpmJYX6alGSkChig13CpUOmo2f93uxW4bxKeFLKdHuHS7wmhk0sFHqeBdVrnO6eCAEBrbkr
KeoF1zCh8s8xgNUgW+JBpNAIPWyY9TS7bk92hWZWDtkhvVp9yokWPjaicqRsyNrHXDNWEzBO7keS
HBjsVUp4n0lr3De/iFp2RCeal1XdU5WebQXjVhxI7wlpZC9yHo1Q5ZpZ7KX8WGbJbLCYQemmaOtO
9bI616SXvvUW6y/6s3mDcVSSxlTEGXxBGXM2h5jcFpyah8AaOhWo7oJ8D8c52rdpfX6Ok+GnG7Ej
SAsEiIq5Imx1Uka55ohjgB1NKkwugB0WMx1QNncInSklzG+oYq8mWku+OKZQX2MkOXOJ6+zNgu5E
86yj+tltkh1DI8VaWLiRc/02oiNscKzK3k8vjqT52lJjM2vzzTqVxFiZYzAsAA23a9LmuDv+gkfD
AI8QUaHMpmCYTo/NUYUUFpO5JgO5JkSkb59CcyQ1FMWe3YVA63MZr/odLuxgtR3XOHwZxim3Lrdy
d56jw9GyOwDKn8fJEybjYcj7tFQtVwZelfK5WHMk4WEUbAfZkFj15Ru7RUHV1CWaD7BckQiLT67O
BXsXcomqNUKn688qZ1WU/0uwnql9yud4PkXna6NB8u61t/EZrgGjXwVuOzuKksK9lMRh6vy+H9BO
8MoPgDX2PebNjZqiIeymYjCDX/HmVWm3uZhSr8xcRv7LG0pG+zqTCGpYLg6fXXHpL+qwdxG4+bP1
pleb86xuBWmRS2uSCbbxSP4SM2d7b66HhdJ4zT4ChSKH7PBrtzulmmFTsBVFZ9EZbb3FELnRRuGm
lzqKHH1OUqO/acxd/TLyzRErbT8B9qe81ZXV+5Wiz0rW8EUXTqEh/0sfEmINy/ynV2h6rXcaqTId
atbIl3SP1aACV974id71sIYcBtaRWqYq4Qgrq0IN5RH2yWVXVYGVzFAoDUv1HvaieirXUOfteGru
UCwzg8AS63ZktMFoQh7tuZA+bdSG8+T+c0dPsmnB8jaCcvEkwbBTBLqxoVHbmr9W7Oij3OiHFJoT
insbAD9ku6E4FCNr45ltsNxUBL9YbwbZz2W24oEustlQ+ILmmAEcMb6yM2aaiXS4nOIP2Bd1hhJ2
hA+GUkhKUN5+ewmj/GplUC111Wk3DiW0L3FgQZ3/NSI/5NaGBhg1ZKYz8/8+TEIB/5Hx7xtL1c7B
eEtELwA18YYJhFo6zBwM1hBD/sUWOty7ggnevnyDsY7Kh62xggGrQO4rXjfwfOZicdYWsP6vW/f0
k9muT0iqAOvgDiTZjisv0yuBOPtp4GGvVb/nkc/tPQAtPAsu1imkGsB+UIPS5cuMWRXURoPjB4TT
QZp/BfaLv5wGvDH5DDP137hN6bSqqE5Oldz2GpwzQjFETKBOU37rcl1XrzJNGzAVcRR8GJTV06Jk
dhanF19c2QtUpI6OmlW3YbPJISmwoKc4m64ftaH8X06HKH0QEUNT8tUvjgshaT9FchS3Cx04NI2j
9ogbzf+P3RHFkDVMZqfbqGb/u6MxWVL4Opgzm45pAeTiXGmPBxJFQfaPOrMpglmJPu65LRQljKnk
STcraTu/3EwCI90VRr5G6pySzkLf20wL5b3DFUD0xYld3zJGixBKLw3iAFiELjKer7bG2XYswkJr
Y03FcHCrvPAcrBccLoeu8cqQvLCnBdi5AMxfOtSP7w7xmJrs4h3kDwQL7slwmup777X3cD5qEEp2
XFgxvch35qFQwFVUEX3G610r322WC56qZTHaZKARqYiPLA0dlsVhuW+naLfsWjcKn9mVrkHqJ3vz
0HA+c6ayttt0tL6zJlbS5uUJmRJUrGKaXQytQ65Q93HSDccFrEvAGkF22FoJLLCtyHImnFCewRmA
7+Zsf96nnBmpP8z2P6EcboasprNGvxF5WjVksYTqe9MK9EiFOXCXNoq3o6HQGdS4gZcBbDaj6veB
1rX+xLWeYQBQ1UBgSanjmAwkE8JWa4GwQdJ6E+j6FLrX1oYmfeBqkcsGdGTvLWPqN8D7EtevR0Q4
k1he1IMGFUgaEZufse2ojie1Li6vIu6F/cbpclkAKNFu8eEpcAswB0dSI8I7Qu/a7iXQv68n9pfn
WNdQlOphpCbsozPG6SWeBCDm6xe+F0f5M7bijxA3HUHkvnbgmK38PlYuVm2KIOiqij6PvnVHYdeB
xsrZSchUbhVLHR2f5TmDUpapfGQt7y+LX2oeIq3ww+FIFQiAjdmDRTjbVpeBJc0r19/Kv6qhmLTh
b83jvScfEG/y0lyQ88s3gtSl/6VhnertotYpDrRbFowZN9W0qXBucNjp7nWFpQ0ytPLnR4YdMyAZ
3Scs9KNdLQYSgVbA3bk7V8b9Dc9C0ILxJcldDiVaEqwW9UOViqTUjRsnZTuPRhwfliANp1ImMwjG
jfjTiDDcvB8gCyZZ7OI4rylj8fI1lA0hFGSTIA0ObDo0BVCEXWl83aEqOxRYmH6WpxDynm0QjrLo
cUBlhPLN8ZbC4+jezUN1nRNJMm2Dvr/ia1N+rbDbxLfZSrirctcpl5reInLnVbrHR9lgvmhHCNJd
/dlEh8CeA2kFLp+aQPzz9bMvEr6zF8Ojc6ZzzKdso5nbi+j+qBpkVrSgNu/LrZE9515SaApufT//
6j8CTNnN38fQjyHs5Uc96QOdnad5Yk1O8tLGfgtmeEEHlQsFhL3yD2OOm4fEhGpb/U7+Vk76Q97R
D0f5IRe6Wmd0jBDFAXhaxDIqMMMy8bPUVou2IlpMwYsGf4PmSt5ltkaEC/aAtdQcctVV2zrNUe5c
UhNjDJ/I8c+jufcqkyRV9hJtSBiLSr//cwzGAOmEHxWQY7VpKPGWUC9gWVu2n7RZAWgvucegZ/kH
KGOihTXN95bO41M7tCLruQnuPLyx/AsWmFp9HJQjYVJ3T0pYmZSlhT05tdFpTGLcuNy8XkSPjrrk
7IzD1wVnVu1Jq/zqlR/WzJHPHp2dJl6ApANbPnVGDcbLXGGUx1r81kEm9mIishmAh1uoQ4H1MSsu
8yiQB5MJ8xgnNRxIGbjRTI4xlNSmIhDGfqljov6DFO0ixv6PPISfxMne1nnabMKYw3J22fdvovHm
6RtKqcwhmwOem/fzK5MmBYe0qNJVPVapv8ztUix3Dle9KkNYb8f7nvAJ6zxXo2y65ffx0O+2DWW5
dWI9rVj/YSYIP3OUMUyrhO3r0OVD3sjgIKUe/UcsY9A+r4oXSvmneaBcv+EYCWhALYOeVwO5GXTc
SmXHwyaVJ1otQeXSZB7UEAlsJLwNmOpHh3Qs1uagxwTp8saPHd7YPdDnosnCoHKLQQLKXrRNZbwe
hlN+UZAMLFZ+boj3r9US4jOY2RqZbnPzhmZeR/RrC1cvRLcJ92g/Itai9SBItmE3GSbFPqyapExE
OVUKF+Va1+bdZGsku9iOtfIatS7yG4vlS47K6LG5SkSaxqMkpK9B07g3YVA3zN2L7IhDKgAKS3dl
t1T0gWVeIXYb3+1kIFujaqS/2vbSDCsNbWo5njuFLMx/poiL05RCs7tWYBcBjhPwtcHft1EebqxK
SAl/0MXg4ImXrvIOsEV+2WfJXj16spSLH4nfVHI+WlnqSTBqs0DVBu2tAGLU0HzCxIBStUmwJK6l
n0OcdSAkROLlCNT4qcPyYwz307bjVIyhX3C0N+XuvAIhA5UxG2qRoofXhzOseTeoRlECeHdSgahT
viZ7TNqz4WRKSfyARobRFy8uNzrmpXTdabukiu4KwgZ7CJV5oDFRThTFOw3a8T1EzpCFcqZbs49e
OFl6ZKnSZ0jlZzKstCpAfk8evuuMjDxIxXC+stzPQfoqNSdAnavrdH7zx0w1P/LfFMjA5HDWoAcA
ZW7zvwQ1g/9qY3OiTcWaGkSi90UAzDMqaarVRCs5+gulomTMIDlyyLH9AYHWcQzxa+P99oHO26cI
p4JHiizDToAca4y/Xy2ifCeHiy3Tm/UT8k98hSnZPy7jBXFskYfAefEMS3eT33gRo7qJRRC9LdDk
dB0Q4j9GY9N2vtk47AZyXJDnDVZU5PI9v0qrw6BEKwGzd566PuEWTgNCOwiCTG+CQledcL4KCI59
WKh0kcg017JIkz+3KTbammvX7yNFO5D53BuYWXTQaxtiqQKduMEjLjDv9gC0skvMB4ZmlFmMuDZ/
fBEORaXSfkx0N9abT0FQmG9tD31sxHOo0xeava9i3vdKEQ+nTr9EcEuRGBJKKWVnSlrBdHc1XJw8
rf9ST8Lgf3fDGMAEYOZF7x3lRVQiu1EoA9YwD4ByvFVqc6PHz96AYgwUUmrv7ZI2p7JJzDScBUKp
Y96EJYUlqh0aQRxdNHbrjlTMnrkVU2UG9XbpsZV4Ef4MUN/4OblskTYPq/5CUyPHblFFsfDqs3xV
wrXSGjUwknVA+29TEQ27R5qkuaWM2Zu1OjHpvcqYCUQNT2p/UgKaDn9EoVpxcrsXMmCPYcSQzfE+
tHfW/XwW02BrEMKXu3NW0R4W/888EMr2z5pdeRctDdpeinKhQ7QeuNyQelwVUKgIROsqi1DLwAOb
zDXPnLw3mc8MdHmcShELOvk6fTO9ORvt+oJY/KhJ9ZaR1qpG9x6IY5piUWL0cYou39HnB++aXdIn
GBdb1Ee/rqdmyDRAR5MjBiOMFzZ/ARdq+J8EXO9T8Zj98Ir9E8DBeXleCIPP2VFYt69DknLZ6GpD
lmelPJFZkiLJgpLinN3AwkMNBRpGHEgnkCHG4ejsrct24K6/QUCQw5dE7HwSYjPALr9k3F2fhxwD
2+og3bXKxVLv6FI3YAV/ZG9DepD7y7wnyHsvqvZqYyxnIFEMC1HKjlwHSsIpF3yPB5oUrK3oZYVv
v1oVA0ecWMhp12V/x89+vARUSSr4dDQTYYRfZKY+KypuHpS79STI3LGQZgpwnb7/A6twcs6YeYlG
GmWX3NtG3Qw2SFnuuLiyUFjYdYw/wjsyz6D5xREgOsy6Y8pv7zwSctHLEZQIm2Pg9ZgyYIN4EoFb
or9bpJwoosIQzcobVw8O643gTf4MhJwZDMA3B2w0yeMeopLig6K9zPQC+Y6CctRDB+P2LUjNJQBw
E+U0P0nMsLylLZF68N9hgiaSf6LkG5ELp28Yx09apiV+N1zHkVHXfYAPlVxtklciZKTXd46n6o7O
4NnWshLjwWsSi8RkhWUNIBB+dv28CH21+E5NMoKdwPXJIctJRtaGz1/vfpMNpRrdAldNJTNZwo0a
xtQoNAvVic7wEdBUXHxjCpE7zhuV7thpDXQI9GShgXLGOfwPgeLX7LMRYHD+F8svlOPprrei74eJ
oDCSuHT6a04RvC8qVwWTNargqRwi/MPcAQdXfWgm4Nx+w3UapAIkzgT/T+BdX6NkMhXN4ELGlTyB
qwQnHnxfMfD+ggeOZJp0+B24xQ4tZPIagRGqBA38HQZZjBIFkyHM8dXNvSRdCbQBt1C/vPgOf1Zs
1dMxKDCaljzovY6QL7eQZK+P/Nnd1bwzA1efYNenTqsMCMs2dgKOQMJIr32oSCGdIaX3/ajA3W27
eGInvBRJ85LVRJoH8jfF4wtYhebAEuuD7LZHQL0MYhK4Cb2ILyOTE+e0r8l0/xdTg3MIj+96HqTM
BWgygxhM6t9zCWwX2hwPHe4TtlgOmJO7UTqa/8mhfpfFyzqukvOvme/jgEDARB4izoGtWoKPXZhU
C75Yv11YJg2kOTob9l57SzEh5k8M4qVtWvUwCN0GUfLAtpX6VzYCzZ+1uc3zvPcsxVOf2+0qehd1
F6AKz8N+1EVFoYFF01oazuXuteAWfnOb+0t5Ycscipc8J1bgO5aJUYlW8qwP1WI/rPiij3cW0RVi
TiXUa/YKxRE8YUxhbj7IF2cr70Pui+QK/AD0XZg98RNixqTsD3cXBeXkUazose01u4DVFSdWkepz
xKZk2WKeLs+8HTC7IiVqkelqQcCcfqrKvfz98c/fhavOONiWeZRVnp0QyOZZ7g/f34nyEKD/hFJE
36vg+kKNwE4Z6FoFrH2vDVegB4hiH8z42j3EfK2COUltIGCEP1IqWo3iLNL9cNtW/QdU4DEC8uJZ
3fK/SJeezMHK+YAjZlNhyeHnN5gEVVPLb+GtT7VKsGiQtDnsbBR5TzBz3jEj3A/6bLFw8lN3IdnJ
dxz1sNIso2KH0a8MFFLxfDVPrMI4asQchqYl9ct7LOfgz9EW6kpV/VNP/8wlqedzaOMzsMyaMFiu
pPzP05bbN+cD/1B5yxTlP0oZdXaOoRS5iiXjFpDLTRRlxqxFkvxT9MzSIbCu+IXssP5jlP25ILm+
Igx2sN9jIjG9KxN/gVao+M9B+U+qV6jfIMyfVtlmG9xohnQJEdbPcmQdbPe3qF/6relb13Ib7xCB
41tkhU6cEqLepc0Ha0XU0ceyvAa5QIF1fAbBqZ4PAXiQczvYbMPdXCifG4e1VN/rsfD8ePxR47zh
Xaq1cstDjBiB7KAGaT2GQv8gKN2IqDvSF7Y5KWjgTo3WVlBom6ArcFW0cTF4smKKg1yuNn70P3ER
bXbdRq4pQkWly0B8BK41LmFQC2LmqBIKMcoV6ByUNdYF7BqN25/4nJ/CsJIVDqoFcIxc7b1rsQNb
rkVHh6/Cyl0CMYhtTBzy89EjEF97fuVD4QXqihTv9pY93gGcKT16u/l8WV0E6UKm9Kjbg5kHTsBl
5/AU2BJwM1ocGy4b1e/0fBXE3tuKAj+CCueKYJoR7VosuptcWtc6sbC2Y96oM89QhcDh4MEJx03R
WVYLr+wZeZDUu8+2nHQIFfkd98V9h/U97wMwksI3eJwIN/22gKKKTMTfwu8cTpd017V76rOsq84V
Ls9vpdbhjtXvwUhttIIPEVeeJ1aRQj2g3GsA5kmVDe3+3jqBTIh9NCZtIivDRx0yO+j3wHG+iN4e
23Qlp0PyvYvvNiy/meA3HZynP6sd4EibuSwrUM4zaxtTA5OzHwcAaswbAQuiKg6p8faUrwDonmdI
UiJW2kMlUN2Xxc01KqTDw66W3hgCwJm6rtymT6QEVyelmsCarODpjz8dHiNxJdAmsi7R8Es/fKBE
O3qxPhcn1fq1kWa1eK9IFFSMw+H2dqQobkveJhUlaubuMBvhKVyIKvgKItrPJQ2Qbpze8HrKlRu5
d6trMZUYkYHxHceLBe2S1udA+GFNmf1EqcAjZUlaat7NV5zOkfJeE70ZfJN1UEBBLD+kEgi9hlrQ
tuDGf7dprgiYmtRBe1Gxe3h3veXWJoImnsHH20SjjEG0S2JkuZTSAkenM+t45le2RuI7ACKLYY7g
6U1SWdbpNUKz9vP8fNQIpFW24CskP90Q84SLnw4h/0sW6ikFDftHehaQj3hmxQib9qwJJFZW4Zfy
eU2Ox9UtQiyuclmgJU49ue2V/5fb4N9O9ZthDKl+OI+lReL7aW4dB7fIbLbJ0O+BVVTXWdEeW11z
ojpibw3uVt1fOFLK11keuDf4Z17r/5kTN38mArpvtRy3+EiuQ4E74neRSeHXJCcVAS0Yzu0Cwvdk
ilvb3JdccPHNbQk6pYLqalyNoa1og4gQ95WSaA6oFGdNBwD62f2bujbDb15+ZUhbmiG41cmDHgdF
Uo/E/zaZCzLAaSCT19116IIzVPqXyuAFS7wuAYZ6dqdkvnvZbkXGVWSIfF/FmQzV8hVQAvafyGSr
iCbI8bOBF5Ydf0/Lkahie6rAzYuppgkmgtoI7SudgkjK10A6qvKTKa/+h7J9aUmDPwWriLROyYHc
4QM81XsMKKlSDMWfM+Vukk8fEzYMCuGmscpzSZPnqLdjJ89QFkbWaMzDdPYOtY1IhsWjbBgd2Z0g
e293ekTKx+awIyyUGD08sBoNLdsQy3lsda/aZ5viHuNTK+zWUVtEmNGWe1M9cnr8EbRUBomt8hmM
Uxmr5VLOO3h8E9uoIX1P2xlIa810i65F+xbtqJ36N8sB6+3kB/kQv1r4/b74YnRYowWawI6m5aB/
hsQIlWJU3m2/3k/DNE1PxN/Lrh0cMssZYz431FSQ5aqR3Btit5NfQPyti2ticWSh8Pkgd2GZsnE7
mbUf0SutSx79CLep9v9oApCQnb97t5payxzDduSLSHYxOrHDG59nO3mSb3bUO5foadYBVJ8fIbJM
6o3rSJe1MxlfCEAGO9qODXHswUEmg0ts9qgHnBiKZTUWTeA8JowfU61SrnQWJnB72frZ//yQu1qQ
vrBBTLcAnxyBYG78HSIFElWlAmyz+4e0JByYT0Jh6bzM0M9Ha9rCmscIF1USNX4E4/pVjCA6UT0F
aPEniTPhlpgNXD1I18TeVDtkeA9jqVSLw2/lNbwoUFuxIPLWjEjlcnGp0YblxcE8cJ8A+cTjyMFa
r6DOIDWwCsHIAdKbeR2CiRhBGfIpYyP0Hzb3WIbWVMKazYT00G3seaj2nsJUyGBh3/aEOPKCpz+H
5j9aPgSILdrnwPavtGm7oZEG+3pIVDmS/UEYyw2RB8NchCooL4fsFOYm4JXwB68Co9l2WWt2ewW+
sLveheJR4Z4hgLONm+kBDBm0DJidhNftHyWI0WUuFAmu47uOP0RhYtzDSoamLI2WqtIomrVKGB3H
zSYMqgACaiI6CtAmDwRrduE2o19ybEteSP1HNXEtOjRhk78BdkL7mQio9G3kp1XxWf44GL9Tjsub
0QZhKUckID31RTK02haXTSX0C/j3MmuXj47G38NT1RL3cORYqR1ujrUWjPC82cVGRyjAE2ps30Ic
8PUa07x0NuMFX1O7B1O+Klh7EBVVH6pXpkEZM5n2ENkZMOD/yg1bEAuzfVMNd+S1YEQKfpJbL9PU
MEbinXtvnoLtwMzryt3aKro05UI9CSJ+EgZsJEYy4jH5L+fIAYF6PJStB9Ew9Hj+j4SEB5a1bZTr
3L2G2BDgy21D8j147rIZdGO5lzjukMCFGOMo5xM7BothFzbFMLd7VBzXLGHRGOL95vFmi/ab0aTE
2sgghumWAtFa9MHiyk51sWNyoRPUd9gjyay7Gqn4nkweWTV0MdiRQBg/ghqDDlONSAhD3BbvV1w/
GM9+e2DIslwT5X9hrj1b+s7e6sLAbgoMsFCTKgJr7MHiiB61JMTntUiPctNIsEpQNY5u5lbGk0AJ
kisX+TL6hxK/WEvuG+nZBb6GGIk4BTtAlJkamLGYvegbhhK7ZMyr46EOlLZ+zmdtKNfWLkrEXtFz
YPfEle9lwjVL3O6iUYU2+LGuPEaCCH2sM/eUNKpYKPTP7ePeKvx3k9OhtDKLWx1h8STCezMS0FSs
9wbpBbxeWm4hZ6a2UlMXfLN05f56UumzSv7I6Ab0kAAh/r6HoqSMXgoELX0PGxBaGqKVoDKKZ5WO
SGoJXAfCRzd97/Axf7vX3emaVffHL6PMXd80W2IyNyn6EStvlAinhds3QxPWJXvUC8Lc4ob+cmZF
yft63JBg7lotQQJ4r9a1R+JfMYDzQArsnbjSgYHLjOgCK0LmkXCmRj5K9lcOUR0tIq4saMbe6l42
gPS8tQIml+9x1JGIUqR5+HCXtyMP/FuFnL2UYaKnpXbBLBwClKTsewDjrHUDsy4RnEP7Et43mffG
t2fwgGh9cXrpVMdpCZ7D9B4um/mnrnxT/gKemxllKiJZMgEOxos4A+x+4GiCIpw+pMAiw1GJnYXs
Z/9QL05nezfuuEnF2/PrI7xVvJctCQk75LXdwrlbh05nFaliRPN61crqqdC618oW1vbJ1bNnwVUg
xypKyZ9e5cp2gE7pRW1PjJrpN864aK0I7MLS5M0wMNg9zZXoUZ06qr68NFTc26YPR8gZsWVHDbgS
YCXpI2thJr/DrnSp3LXGpJ9e2wAEMAHUe/s0oLHUZcObop5QQQyEbxphdAPC34K39ybXnl/hNCVU
qJETa+mpLjMpPTZPPakLyNiqg1bIVEB2izr6kdmIqWeBGHvd8KlRXdsf/9WdKSxWvqhMd1znEGnR
dCHjm12UqqvY7wJlw3CgG93B68wk+p1A1BWGLP7FVTRMlCp5S3rOGtwXABHfAmbThItHzqB3x1pn
Fy8h5IFuDrYHyBsDj/IXzgXyDByHLUtd0peAtscFMBGOKLQ/meTa4qY43BIaKvzIeBJR8A1TmpBI
0fovYYFglY1ee22ga8vgVuUtNvQwER0CBsAc9+EBEpBQ9Qk/p2PYxRglTEgQeg5KlGf9vO06ymov
ErffSK565jj+L02/spniUoJcxWM8b0MmRh4rAIez9Q0S2BiMuNHXUvWaIXoWGWs7iODEyKRMoT9C
lOtquazZa8JC0HGdz/o5yymXnyzm8rytg8uijoVabHGGcEtO+1Eo0lfBRVwxXDZXqpMskEsq7Gfw
5Fkv25cl55LrR3bOvNBKrpYGq1n3i1a7Hy2NZg3d3dcKTF5EBARWSY/NIUpzZ0VFa/1Vyc9zvvk2
dQcTjPOucHvoW/i16STelW1bRM2qGtvVn7ga/09LNpdaYHya8w2Ujf7WMnc9JAVUll3Fk8uGjKAe
w4NwSrF2rEGmyiQ7NJGObNX8dvvQ67h5eBABPe6I7tQjUez5joQVgoc2OqPELE/1D2vwEhqWJNf6
+Jtxxe+BdNi5ZCXLOe7YAO5Z3/mtCBly2eDdKSOpPBzIca6k4ByVoQHsQdnhPwRyGTiFAT5KqRcM
x1LdoxK52wG4p29GFGGZntJtT2G8n2Rhoe1erHopLs2e0T2oeha01cQO+RwdozdcmQzBkUHtBgM2
6ObZ5UN1RmqRNAzvtdd5RVx2u+m5c89k2hwAhTwoEPAvuYUigi4EsjRR2a58LIic8+27R0MMbfXB
cXf0IA92MrNe7e3ShxYXCg+EPIFz5HVBPRenwALmb3/3v2djsHAbuEAgXF7XRpOBQa9WiR6rkirw
H6wFlSap86/q9b5+ykZgM41xYRDMd8dnJ7t/HZiaL1/G1JG1cCU7kTJUQGEpWKpAZoUfOFwZDiNB
8ldnZ5NtmfBZbRFTX4zx5UjXSj13N4MIw4nP6ktV5ajayNCchp6evPeJKOX/RV2NibTQa40L2AHR
o7hMnx9Tp67mzg/4m9SbOsol/G2i0JpogQrMOXuuW+JKhrdNiVxTz6Fn8durvCad8Z+r4SzXIbsO
gzhvD78w7ARsllfyM5F21ePDxPzEzh/ilGTMi+45Gy9inVkb8R2p5pzcaBS4NRA2zaHGNoIqLkCI
4iGQwS0snSJm5C8cYHiVd/CMW+4wUwvY96pxjJP/eB+nc8NXu2WodNEzdlc3ps/1AdD8n+VdIznC
oO+dYxfI2fmBAf8qmVLerzdJJqLFU3RkY3TTdz/dgCXijgt0CiLyew1XxqT1WgCDoAoQMdoowxjM
5KaQOHpIriPgPvF1ZTs2vdsGPaG2MNt4HgCB7Ii90OGu7wjgeITxOl9lbbKhWxo85BWRyxseJk6p
0F9sDcoGTw6PZeXEaU7eC3o4TqDBXP6w3INi39FHFurAh9a/ch4md652fAn8nh5i82f+FFkv4T9V
qdSFAHk6SedozItbrtyhLEA1pvVC6spnKpwDfvcjMgqRreJvKkoHPap+sERgjPqTTWOR0CRxHMYI
cORtjp5F/Gyqa2O5mElTxoNk73RAlhYeIiV0iazFmROgOgCgW2bAYaO718nJTylk7sby/cPRQalY
prwjLHXFw41gpWPnxuvFdgiQh3nUNS0P55pb2ZLd+IEzVMgP2+e6FzKXAdFay89WSEKQFX9GNc6Z
zozvUYMOLs1QeJ4C/sqa0Za/q2WeoXvv3vH68OtFMyHNqgF+jOHhJkTG3PWCoozsMooHMwacPPmZ
VOHx56kxlaIAoKHAdsZbvNacgZwKneKlGesFx1Ct3xSNMLa5mhLUzmwwBu96/FmssFtQHLINwFuT
4BbHBVbTPpLXYYGWQn7NEvUy2mPNIJtYjVB3cAceJz9I+Va4fRVZW2J87AAgmecGB64gqHcDKDw6
t3qMZTu1jWV/wFnL3pWhn6gbAArMcSxd5wwbDwBcQ2mdAAQNpzAAZ74Pqw2l3MyTmNvaZbWHOyIm
KnzmhDci1AAPcLb2GQ5NPVJ3INb/BcnLAX+Iy4AEYuNFrr+xPSVIjr3SIJ3nuTsizw05DkTiiFeu
Yi3kL7yea9qYfo4Opv23O4YUfokTe88unocbhY62sXNE5lqWKquWSMovK+9NU3fDpPt+Y96rzBp7
j0UZYhSbPcrGxUtS5r0lhIEI432QuFRQ5ZOmZ9spVHGN6RsIjjYpMh1E6d/M9vvATvbx7X5riAif
Y3DAyX6rc90qbybJH4ge1KZk2324o5n5lJpPT7tLCG79dpDB8EBZsZ3jSzxuoLx8ot/pXOkeLcas
duJk7ZIByR4/l9yeo0LS+r+R3lpzeuTiF86fDjYEL+AknD6O8MB9Mp8JUhz9JxfqBA73ojNM/AU7
zESkE9jcoHBC/1QVnIAYPKtopPaex+SFxSH00Ym+PZC0NLRQQOTpMLHuc/oHo1YSn7MeDzL0JO7V
s0UKP336W6LVpd3wBVGW5TXmwktb25jZetdIqJUF989tARK0rV38nZSA5XqQ/lgi6CGCmMWHKlH6
V3i/ymSkm74noOroHKhGOjIl/MQdXEW7vtK8K5QQ52YWVzLyrBx3EemAQJbyoJL/v7Wi75+39wzd
Bl2gcMZeniQpuvqeBFcdOB9aFvAZsl+3w2RvBej8ohpG08X3t0Ssrnopc2MApRvMD4z2FQEVroP3
QUcFWr4k/40m6G+OmbbO9p3b0GYxqM+FmCC56XmVT61qABFm1I0JcTz6MJvkZ82LWrhUK43LH6Vt
UbkG3xe1maNLBTkRyWbccA8q/urx9Q21SQykG2en76dBVv9xWukyroXnNQwsoSA85JhdPriwS/Sq
WnrI2BGHU/SgnMWObIchZN/Nybpfpjkrlh0VESK+iI2IeH7PIt9FTsveZmMeJZeTLlVP5HKkxS1c
tfoKFOiVrZsVl9np8ryQHzXbVrpiX9U1cJDqp1+hnPdwmPNoywyDWTiHpoGs2635E8KqQQrDMmD6
x1FJf4E2QQXAnER1nGknf+al5AXM8GD5/y1/kg0JFjEb3icYaLLQTL+P37gpkGJTKsK/9BbpIe3r
81SVWN5n95HEf2VBSNea7605YaINkp8e8zPGwS7BHHBzCsz8bdPKoM5wCiW2raL+W0ihm+4pMyy0
AK46cj5/CclqNXYIwnn8ccATfE+Ks3jiWOXWQfjH9sdvZxufgwAUEtJe6VTrm85Qgo2BqLzKvZ1I
S4kCf4UMBF/U1mX7U1wNd/Wbc3XB3FmLwqK9rk0jG3rN4CPzMgDlZWUp/CZf1PDu7nvMpW59Kr35
RTMJjmGJyRFueAckdytUiiCstcO2NjwVWClHEQSX6Z3CRSvl1vWq4kzl6xA+mtgZuSc2lXe6bbEW
voETrfYyxSXfwXPyMXAGDlVT6bxFt8r0i3MXQwkXUHBZ8Ft57r6kBRTxx/d7NB1EKMgSE/dFANXE
gkVhMRKKhQAibjOmEf/TCLM6ZAfgpmFOqbQRcmsTGRNrsSQSmFmNst8pnlV3id7yESVloMeaKbS0
DJUK/t3RztmH5SH8bz/+j3Mkb99NSTXX173+p3fMj2S5hnDIr89IP4Zx1A662+7MNnOV6bzvYnV2
lfyxo+WcNS8V7KIdFD3FuKmvFgM3P7tgdLUsOp+J0SceG+NeJWTjHdqmVorI3olIlIU9s2dOsN8M
8fNvHn/uAEai19vPnseGbbAt/x+ZQ6iCMvmxtB7+nbRH86wKmQxM5H/T9QCzn5iOs6iWc4S3g8y8
+naPYNvSM6eThUpkHmkhrTrBRceAZlcHGd3oA02Ov8MH3VXG8qP+p7dQB+O/IUSBIfGXv88zHYe2
PVfH8skxNjZa6zBfhfTA8oqOcvDuqCc0efPilImA9VXa5SuB74DKl+PwW0uPT62g0vHzef/WjLR4
ifqeaVzDb6UAoiRRXUCXwXGPvo9u7HgI42NQreAwvU84Ds0f+WCPeQD0whjTHLgdt3YwUKFySmdo
hZOYqfYsyix6uClxZtS5xoooU1s284nxUeN7mjWLQ7ZFq3KF0w94VV51vpPqsTzCflBqK5t5BlWr
T5jYZARTlgkcqDPXUecnn5TPCQeCoT0+dnutgmzkQu5A5uoc+ZaWFq8J/jI8sLuHdmmLJe7A3in4
13f6wTOX3sI+XSgLypp3EYbBydrQmn0oPmI7ZEhsqDy/4OlTZHmfMfyhIYc61BebnjDEh+ykaWge
8BcJqsc1hUj/O76fyLRwKSM62hBwJVkwDNQQG8B7g8/J30SIvFtFUvPTVsnv8nGysZAiGqjFUdep
hub7so4HAo9Kdmh3OKbo9ejJkmUyFHOlK6G4ziYj78W1VL52oDRfX/n/sg+4hk/9wK+ZPKub4h+e
QXjUbqSJMmpsmGUmQG4ndbi+N9v8t6QcKg+EwCzP8kyx2R9cVkJk5S/z5lcJVRXUFO3Lv5rvSPsj
atE4mBUaWakFICrteEys22ifiegbliyW2574oYere+F5mHO6V4iYq8nju32t9Fq/jM0AcaKVcjv7
8gH2QZQ7agye7qe6Cgkwc/D3fhP2RIBK5PHf/Iof8msNEkRoNpZViWT+4v1Z/zRD1IqorhwoMXfy
Opa8tzmCzl0Fb8U3/JaR15kIfxjXkaDO6wauFDB7GQT5OKwu3XP8RohPbxqxnu249RaKkL8V00BF
/w2DZKr5QKfA8mk768k/+UUwS5/sd+R+Z11U5ZTHJOAbaCSlHYXyWuxRh8RxiwGvaw6GsZWuJkXU
pk9K+vEjlBfym3OW6tOXT3/dEREdn0rQgnxX+jYQsMEef1VMQTaeE1xbkoQpgUHn5ordX7YBEIFD
yDoRv4Q1O68I5aN4UMu6gcxHnC/srGtVFR33sUj2nzd2JYofahK1RlLf0twCE/bgYWeO/VkMo8N3
KFowN1mr2kGl/NRX+nco7rs0g8ARMBiZXmVS6q524xmj3i2OyDUhRMRMxeAd8RDTi2Y6EX99dxvw
OYzayKpSwgSKAIAbJx++vQGyVJmWqYrY7keXKV7nCBL3w6hKEeKksDy2sCta/I9MvNtqn9JxO7n/
6o/ep9FYXTTKJ77gpqIw3Aheqx3FU6glgUTF8aSIGQDlWsceXbFD2sGwvsa/8iwqFcZanT7YCL8u
G+0eU1FTJ1LvsAc7dLvcNtD71a72PAzRj6ayjBU9Nzq/FWQZSJgwHCurW0E0mfG9kjkpEDKX+IPG
XS93zsOYzKUeJZJ850hof7iRce2EGIOxIB6LRR0r/KxHlkypQcnpMobulHqiVPvnswvvIIjb/7hT
WyroBWURTGdoPhBOtdvMNNVxVhwjDWDQ8tIqWQV9Rgczaf1Rs/oqyrbPCbVB1LHurtMY0fMzugnM
VriSxIwM8MIrtwgtl1fxHZy/nxb10tSilr21c7RUQEFfkXyJZTNiBBEPd91nWQJUUheYaG8ymajn
GrWzoJZebk7CrAVsLFbBcYycUEgk1Sb1uT0JMFWpmKO1g3UYwkDV4wBuGRTLOF02NZDv9wWQQgmp
MW63Uz1YlXEbN+8n8QfwKJ3aVhlwqy3P2vQA3w9HQEqy7NJ3hiOCS8LTW1VWKE1dz7PtyPay11ML
1fgJEwEukT8QuOgh0EvW5RzMcaILYBG/wAZiCNKmbq2zPGDDiiF8p+dElAyDiwxcPc4KNo6W5bm7
lvqqTzFKVR1njPq8+QEA3mh7PAnf5AnM9M4eo1BZoSo3tPg1excDSH5dtmdm3kDk1vuL+9xlt/yd
eCQ19y7WEQPcb9vRggBUMB3d/Ik41AalFftjq9DT3rO/m7+Ar2gP3dEpRRNHqhcaA2SadC6i+sTZ
9N+4Rru6UyCnpQ+EAnVjFsQMIBJ0+MLd52jzhtVT4afZ+DtHLTZ25hw2loQHNpigZ4M+M5Pj+Mce
aCfjrGVEvXNgObi13edTfkbKK+UOG8B3C5ATnYdo0qHc1c7eKX87KV668TrW7txPKO/gOWAwSqFr
eu6YelGPbFYcodGqD4cDixV1W3Hqx4c+wsU5DriKwFI8WuGHbYjfWJO/TZx+44++l2ucQXY9Q0ex
HJZxT06QMOHqgghVo2qWPnK7iA6ICxfNYbhBa8rETF4wHtpFoTopa7wt7G7mb12iyvegC6B9MuZM
IcFpiBkDdo5qN6604S3YhdBVj39y0Gm4f1wJPV0rzxNOnTGCJ+ylAp487b1jHt8hwPAzmoyoZZz3
5jaT19kQMZvwW3YXC4I5wAAsh/rt100EtoShxhUVKZcHGN64foJr1Yx5T8QepuzWtEnFtQyAKMUY
vkvSUmp1Fe0uHd3utAabDj9eRTTFdr6vic5QWLkqF8gzSoWQlZaW6ImZLdqHBhQFNLfCQDXC+YJ2
e9yXsoKHX7O8s0ImYznRPRjX9LwkpknbSVu4szNH+trK++Pa1QBwbG3QdITRspkS48BTL7MvraWS
xBxE5UOrF76vk476T7YLNgDHHlBzSc//QWXh4Np4XQRMiLzHTj+w8C3r++prq91o+7kmDDljra7T
l95juFAP2nukVH2SBzPqfm3OxyO0yzsdb7xiZ/QxQ9SqJkAvGsr1rwFEZA2Unv+tlrtXwh23XAvK
Ho68GtKjUGCik3Ood9S9Kg6NNqUtI+i+aGfP1FlrU+4sJuF099tJboQ7/qFtaHMbyBvfnwObuX5Z
BdAcValS3z+tTlTe6e2i89dWR6vHQ0gwg15Pn6z0Ha0vV+TLXInkTlTY2+UzhmH6FiRYaTmYhgvz
SgvXsEK74R73gfj+Bq645NKKoYIJNgtpq5upm+x6uMV9fAiB+8qGUCR2KO7tBtekOf6fdUAVZeqf
O8gP8Z4DVPWLPgawzeJ9+cVFKd9jd5CBCtphRj9RZn2Aynb3Q7XjYU2vGqy419cYJ3Cm67RWfOc0
0o3Bem7PnuyqHeNcLiH6hT6o2ptTK9KwIfT1M9+jvf9qb6Rsz1bT+BxI2Ngp6q4k/rOJ/gOBmT9K
2DDnD1W49+G+WmLJ83o+OfRtjdpJkG8UbDAcdlqzKShyY4VtRSRGrxG6WN/ynKRBHyMabawWjA79
wG4n4LR0i92KzKjtQkylZmqn6Szy6wGWFNaNOmoJKIjqGghRPia0GlJNSHPi5xbleGSs4Xtsi94Q
trUU5fBVUBwI7+b4sdOipof6b/1BWsi62utfyb3qYE5hSwyubq8UIQ2Uw8N+D61fWTrc78wK9TsN
SJwwgQjf7Pr7f+GujT83UtRp6aymLGTz5O7gsv0JtQ47hV98M8hKlc7ThYh0Dmr0TSSpqXWcsPO0
AmDXeHwWR/meJAKN+uDrSvNyZlnoDH9pWPrMqpsw5rdgZTZvbXTM+iY+FHPPQN+ADgNLbA5zmTyf
ruw8fe7oi8UBrAcyvftXm9Bd2Z6ngw2/XeOernhUGGzdE2xIf62RKjfNSGvC+B0DloDh04827Mwn
tVC6yWPNUBAPjIALn5rC7f9a0hkz7GBhwKH6grBsZuczpXPqn2dlGnPfQH8jXaG0NPAUH7ESJNw/
M9ZjZsWvLM8hpfvQZsyTU1qHOHlaAcyb2jmVT1h0+KoYqRH4RK8nVV34MJjNFZZxG0j9Srmc1Xoh
x37yJFiwZgZuExSxWTQB49YB5wZtSh/kAwEJFa13niRNS4ieli7UrzxY9R/Kj0uJ7Sp8NX4Jk9fA
HWo9YsqUm7VpZifvt1QIgoFC7Qwi/pgUsVAdl41TsbJKopmhVFJC3+AskqRN3S4oDpLiV3MkWl28
0HpOTyFeGRMYzyqMn9A6FB4as2/1XWXu1Rb55YyPEG3fIc8gmyAJDvttI3F83mscnPE2UqLmsRUR
GWrqal/XxYb9ULSi2rUfbQJm3yZRB0Cy5xBZR9P/iYM6T3QY+jXC7C5XBaAwqsSi2jzB/Wk69gqE
jqbvgkSFunJO/xOccYLlMSnknmCNV1mfaZXpDFJZdw9wtIW+67uLO5NZujclj0oVy6tuli2BXOet
TmzJGHa6aOUZlJWofO7NknN4VGVS3294MuFQkmZQfRX7DSKoojDqk/tNyGFi3M6kQ5si/eQWoEl+
jRR0Pk5qXoI6blebMDUUo9IlJtSH/9FXGYUF7MOpFpEMLbl7QySP76Cdv/wmel/4omiB3cAFresE
JfnwAt5JHWWe5oZPYPQCtudRjupigHHBeaBRaftos5LhxLRfayDodpZ49PWHvbJR/t6sgY0OAD9g
wIDh+AxFpaOCPnKSbwqiRAihNQoJSsRw1O+W1NsqQrNsrgLuM7AIa/H48pA/igc6zZ4pp4dxf+Au
j32N0MioX7YiZHU2TgUdQUO0dGC974IRyI3wWOU9IIPDR2I+EO7Cyc14BuoJ29JxROzGFmzaIGFC
5tJX+vB/stZLr0+RjRj/oUfV/nAQ0Zwqw/foFqw0ZD7cE3ctpe7vBQzamzH0nMROxy6DdD0u2O8D
+vk91wDWXN7trkYxRClXNGK6g4Rn0nfKOiaosby8DouIblZ0KwCW7Jjl4+rkDpcIKZwL8G88jU5r
m4uH8Wg8W2rdo7zbULuVXDzD6zFBjG9AUb6kVG719fw712FyNOtBcG6LtTY3xaFjS9OURHY8YiOw
EgjKldVnHPDevj9U3l/AVyyw5WtF93NFWm4mup1mnZdfWEm9jx6u8b2ZrTM3oIGeBfLNRqKK5ful
gYg122Fec3wjo2T0m3NMrfjiduhhm7CUBy51z6fmkr2GSKqeod0+V/ZX4f21R6ZLVGpyvE4Weqm9
WtXjlqC5CLTYAK2PbOH+yolfLF56BHVX55U677EPFDpWp5kN7Vxb4ya4XKjdfK08DpFwW4sxlZuC
7oSK5hMkwWm6OgGfiJYjVDXTO0aVaS4f5y5LsOydmQbcaCmzXBFjmdqJ8gFit9EgYtqitFmWDqeh
eePpBuSQFkpWUMNQ6TP1kKNth7lwVK903zLswziel/0bfDC5XEKCiVBLKw+3tajJMNcwPb4cSmHU
iuQzlWtI6B3zRP8k0o2p61DoAd92yTQb8OsKrBUA5AbzZWntPjlGvbY8UDstiHPn6f0ghdQL3YDN
H50q8O37zooHvTWfaHCZ38Rit7BzYqEY9L1vbDzsFXeRd040WTmPqbJZxkswKR0IjIRIexieiIw6
Js1X0/q4HmuUxLZdYhSbzLq2rgrtXpmUJL/eVsUHHT7dRmuShyiiVAL7H8GKWMm3+4FJc3zNq37j
IxB1kDIYRUFmDqoXaWEfkGPlx6nDs1vxAiQgRo8lZyJGPhUnYvMB0AeaXW354alLL5jM3CjABGVB
98p9cxB7TCaZx1cRSb5yUze4LKvMa6MymkGmTnHdKswza8cZvMKJJoQKgvEvqaM6Y3FBKfsd25hO
BqhBvBfgJZplK/VSSjm0yk2L1H9hVk165pnEZnBWJCmQQ1zPR1Lk5DOCheUUEu+9fyL7dl0jkvYb
82V9wSPT/Sdp+UnvMz1OOsvNaZfPmf6d8dQhHOsV0Uu+5dRlLsuLXBrQtzIr03ZH9PMFQEy1Bm9V
oKBLE7mGnGpaCI1NIg5nDoVlHXRexlMD336z1+m20ybE1kgZg6yboFd2ER1wUc8MORsONtgERt8M
yjzXHgaV9Ldqk2bjPNKAyqnNTxCGZvEKKf+WfwWrc6UJpHWQdfmu1BIrT/sNSr6dgVvvHQZ2X/eA
GPfx0r5IxGjCi4mr63wHbELIEu49SoRsqas5titvhvM3KPa8ezE2LUrfCwoXqP98bx2KgMjJE+u+
a11K95QhzYJ61hsZ6p5uJQegK08asz7+WWZsc1GLqw78qSoYVVgrar22ZSEsxiDGlSX16L1grSpz
xBtPL4QxuL8B5B44kAVgPAU9rzoQ9xZURPnhXPDKWpEKnsi8vwqkI8YXSHdGxTON4SWJl6GdaAYX
XxBluW6zWtfyxynbfXlVDEy6Yig/WbzYG15BXjiOY2vcomPOHyInBpl6f+V61WoHUVjTzztSAGYb
mHMCRm3lkiWpbEHcvsc/G+s1Er9uCAQ7GYPrp0kYGLxjkXx1UqWbFCvFrBbIjAa5OE0AJpNEIMVf
wF1up3iR2UGizbLnkQ3SgI1zDSascbSw6rZP+F4HV/Ax591e0+BfPF6hHk2BmnMQnq2opPDLFbsq
Ob1RFlkseBK0ZxriQ+AUMzwwwevSG2gLJWVwyXERbXa9Vqz2nTmEGuOK5hJdGMfqzsB2QNEytB+/
cKF1v7fGyFKRQuHPOCPvZfYDQwclB5eshbhIu0W2VTT2e38KQxiRrY+n0nodNJSgKBX9/Th+8ARF
LwwI5rABgCdSCXkLtnCaBStyg0HPaFKECik8rrq1nlmGgXT+4kKY9hdE41V4ELrTlIcwPqPK8g0O
AW6gEF0e41Yh8pLXyGgRU607bk01qx9GcygTcNBTj58OiSuGDXuANtk1PQdwedSs9zTYmQKBGoO2
ITW9RpIhPtR5Hnai9ID/hyGK5jtihQeCu9bAg8bva55LkTzrL2PPPufecdJ/9ChsqLmNhB7NF9+o
lK5I9GsB2zFISeNAwabZptR9NGKnSq6rVEyim3PDRJBz/76H3qzqO+T1KLlFTb0CrglLyQU+1jRE
lgsG8cDt85JfH/kKYuWWMBnkEBF3LkNxGFYPL6V8J60hOKluSwJvxHNA2jszfNUWzyvA3SloHhpY
GlYJOaKROGzi93zA4wfGVWMjHnVsK6IrYlSbfpiYDDmyjG9c5afgN5AVN0u8FTdlFPQEGEs/8Pbz
wG531WB9FwD6yCIJx5Xl0vVAFPOmFign0EjQ+LweqZST6Y/d9jIoDGW+V9nxMKCKtMnyEUXtLSJf
C4r4MnUFu+8L4fPUv/rFpx1fxCUG11w4C34Mn3Hti0vJAEO+7SQwDsvo3JyCkR14ISWN7UFAdU/f
E5Ma2GB19VqWTzEisx56ThaWyyjd6Ctct9PZzi7ulpNR2jxUYsAiVr7+OXKsVLcBWRrnb9hcz5V0
19j95ll0S1t+LPWLz88hJEoMqI05uF+ZtAeDoUS5BYOm3wx4I25WLySw4rYU3yC4nrRFpJg4pPUd
9O05KqsaRgT10NT4da6wnEyYEiMO+OKfSH0czu/br9SPgcdCIklwjnYvCegkwmHx4CTJulkhzeKC
JmMgR1QxZvB1SPWs4y4qQ608J9yHmQCw3MvYvKi0fS43iPxM8zGX25pj0Ree7ICFh9HAwU5RLF69
Oxu4jGI2NyfwircMdK6saRBsRJW8skkLLOLcEVg5bLqs0mC3mJM7205zbPsOacUbgIVtNJ3Yox5p
AZrDubWFq9Cruc0QpVM2qfDjwo02wAHsqMd/YqueXcuvp3DtcVUHp73xwIT+WfiCl26f1phVSyF7
82vwbc5txsC9qyLdTllnG1JJ7mBN7yR0gBTOIuuJwry5U4oBDACqlQ5byQy5pucwyQXqgnYdUOw5
VXz771HizT0iOoJVpxxfMqsHNYeZuTsuTvPKWXrwtYjmuxH2sDAWnhlAQNaR8/biBXUOGjLSFgKp
eVZk15AFsgosoKH/LTVlWgKXj3M+Nc0RXw1N83hKObtNUrks/tZwHV94J0ZdJx/0RJNIiqil9UP/
zDjanShQcHdEYJEw46WS3drGmST1t1T2xnerAREHOem15naPYZUcO/u9umWsw557V7BgKPd3mb6T
9X70DSw1Ea2/mXRiv8oMOe/G5ZpvvJlMiz/0jn4wpmJL0kKvocTQlUqkkXAZD22ZWcrii5w4MaKu
vjhrwlx+sWNPw0f8IscoeAmKx6q96b5wqTvpiYG602ROR8jjIFHYUpxXnAoShCdaAlsHIjjGqK5J
jGCa4kn0mRmbkOc2U9AKs9MOvYu3qPVhRlwGJCyViqWGawILBl1z8y4eHv/c2yydGbIB7IQlwG3H
TukKNzz+sS0HiC9OwUu7AzBgy7iiA94PU0iZuPi1ZkdziVsMBA6PY8iF9L1g3WVTKPyrf1EBTnb+
6s49IHbE3r5G3NkXbapklU2xqNFLRIG0S3//rJpyOd2n9O4Gh/5ic2ygxXny7Umb3KgFT7BKJnqh
MDCy6i+WtEXhxkh/BJAv1jmP8XMuw+myPS3Pnn1+Dd2z8LSFtigrIKoIGIVAU+087npDi5FJPP2G
RRzhHgCnC2MW8yw6EW4YgQbuLksof4ha/rryt5lUjVm8hdttk060q451D8KR8ONvhOON6OXDq/5i
uOlDWrGmSA5fmwOasP55cCzblJNg6d80ZIvDHOGnJP5Zii+j45N+MP9bBGugurPJg1U1CuLBwR5z
OXPGVDYMguHYwB3KSQh4eqJB+JnhEBHSQ4q0ZGd6zZWuybjP5otmqPpZXzGObu9VaZx3kjIgTTIy
8mgkttaX2mogjCzAFvHP+BXxT8rtrjCvC1E+qp0TY92YaWWSRRrXGr+KSTacIPkWWQmOtmAuo5c9
AiOBVpP5TVtvBcq1DNN8XL0DIF/2gfsQkdDPDBUTvMiF9dbnyDqnUjxTj5gzRt+XuP9puf4ktouJ
46XvuZ4rFUo34Q6hCsnPIsXATj4aU+NCYZVB+9x5D6IfowOfzV3hIzmohUb4ZhUusmf2+WWWcCOs
basqMXWPJAywq9EzAw0ENBVzQgXLPJsD+d/ZpK0EfqCs4gOE40T8aWvYVue9kWtARKEaED2Y3ctO
4mZoP5Ah+B4Wz4G/T5NVSMkAOiBNfII2K3rDCY2G9m/U03UXlXfmYStZkRdni4dOvADXz0T8SoEd
UQtIdtFKkz7BLOG4Hi4FOSiJNjVk0aK9+laTgGdcHm+gBbAd9Nc4rDKvccWjN6AOB5ZxfLTCag7w
Wp/3Iqllki0DGQtYrIsoVbKwOpcHiIcfhMYBH3eiYShEJR6/MJBuKzUzRQeYeym4nTxm4RF1YKQx
9OAloswXm9txjf0YMeHgMYq5iFZneprON8yyJ4rwhDfUZxErsGC06/mlOiEnp/FuofeugZdF9Xw2
sYMzLLm5NsMd7BLXOoeEL6NiLI3K6FolNiOWB39l/EdX0zlOw5iGstoxenM0yb65fB6yz6cWL2r2
pEP/43FeUDjAhUtUTbVhLljl2tJiCvIZP1TW2k7uTfdODYuU6KDG1PH85E8XuCx3nMU+Kg6XrIDs
WhY0H+zwecUZkfRtmQnKeinvbz+1VVdac4Y/RjDc6SRdln8XbakFVV4hALIEVoCfmV7osUwtJMzu
9alIhoFIqE4vbJPYCVEXf5mFXPHxX7Vvmouyqt18h/skWqt0BJwvNKf7j45J+v/UIvNVS+5jrjYW
rVMcpfSip+xyCatw5rnpsZVkC7Ef8rjXZEFa9VFftXhg40FEddIDXQlbaD4vOnML296ZsBTge4bW
yc9zVPjcqxZehCjLrdL9t0izH0Fru9PRaLLvwT4fUzpNVTkkhNLAIuWBR9ZkVhfz3wP7q4EWQfDl
TTJqrEQdAMmwpByCydTmoT/6iJDPsuJ3H/qfvPe+b+i7cmScjOmHYpzG2TUczXvK5cW8y6NkKEal
hzke0JASHYUnC+yGlSkEfcrphYudhTNXu4xV87iZZUnEEDOu3e4Tj4aKPNzxPbJEiBbhG7o/Qd2E
HVKMlCWmLrD3HTtgkvuViWys2wSCuQe5qgViuq5kI0GxLFXRTb25xyiCy3wmin0ePbQzo452kN2O
NI4TTPo/wEfzMFUD+cPouyCfvy3f7myu9ayPoZChQ1tfdlN7SL9Wn+Ri3IkXhLzl8oacZQqrns9x
e51ekTHO5vgNjNAyRgcDhQhEeCrUNWEs01LM0dacKYWHFTaIXiSiPUO3A2bF1vAZgq9p9MDfzgGJ
B6z7+/+6xtruGTU/Vr7KF7o/yEJgVfAzNpnjOXcBC44zFrIA2WYtJVhIic/HoHzSV2tJLQesp9St
Vg2RL/bwJPpKX5ygFjoDAVriGCE5xQqBQKUENwB/7pYAnGEwg0I7m+d5llazNaz8dt0b5u6Rgp/1
lN8O9CCRxai518nHdhT77ffh5C7wGjwZ0VcOpxX/RKfw0XWNPLZ10Zt9ksPKbHqi6U0Z5hEGRX6c
+JDc2Vt0dfP6BDNkDkyc0osUmHn1CIq0Q2TtKGL/8b5OKNhbW/BSfflyy2eBur1W9EDUX07yCInG
pRSiDJeLCCej2z3L1LblzTin74MgGDPtU+aDYetDRoOKtHuOVLGl7FBxOmF5YvEv0KZuGjA4lIVD
RCGJGNZ4131jiJzPdOLT3vysF2Ux8qAi1c6J26zE8GLrxXOcuqVYs34LoardmPhvzni4m8S+jRaX
SMF9VW1FA5OZoFZ499raoaUjtIZMl62pEQ+Z48hvLYK0p/xX/OgHjxTwLiICi/fJupIHzyfsJuDl
oalNa5SWTFjFttGoeNk7d4j3+N4/7Z6A3eiyaVWb38XpYdL4My03eFkMY+EWSNpISc1N2aCPqAfr
RDFn7fqbOLwajEqfyQff8oKv6PLjYyDmn5UyCNM1G4d6X8s4zIESbLhfh/VoSLlXT62PJDehJvUH
zpbBmS4fsqdyysGoxrojnTgkcy8f51fjdFO8baDxKaZ9xw9pxmdV5tTebZu2l+OixAD0eUtpfzkU
YdFXMJ1tsJsdmDnc/66sPr+ksEuERQy4bnOrGI7F1w82UaXU6uW0W2yina9POza77qiJMYfQ3vWo
cEQy812buwjwQCLbGnVzMwlRuGwzKO9K2pdZ9S8WD/90svTeVdglnm8MZ7trg2G0fK9XSv3k7taO
AC0JwAm4zaNsqkICkiaaBN7AowlEh8HyqEE/gjC5J/IENlw9A3gElAjtwMM5aic4ewEBU7Gyttle
4CqF9GUepMYS52lVjAw6hHsL81fmUyJX+lYmnrJKLPzbUIndEPI6PMUdawCE3TAsa89f3VjMNpqO
hhb5Py5qXaRHeYo2r2T/kCnlnTzY1Wc8W2AbDmGzwTkmc5TgaSFyF5fIx650ha7/X91S8ptWcNPQ
1n2a2fHW+VJdt406gyIWnKUF8U9w3YwvLY7SQH3NjS9RvE1EAoSoM0mGQoO0t8Vyt9B0mMTaPPmg
pSNAI4cuKFVBmGmtLOalcVNg9SKIS29LwpseU0YXq+YiN1i3KKcGFCJeJUKvpkwKcuFzneO0sYrx
l6FL4Ot6krv8p98YVFfc6ihlGG4khQFXCFD/NXNlRglLrbjg9bqeDRA89cEmiQDDi9AeSJ8ByhbP
Xo9AuZhxakO5G+WM53t4zykPBDYKXENiLGOL4VfS8K1WggzvufY6SpBUr1RAVmB4bJfCujeHzIMV
4UIZ5VvWl2OJKVniKnhPE9EHQKAvyx3v2NzuunfB5FjeRtoEMoRC4KlW+zud2zYoLqn3GK/TYqCW
niOXX6Lgcre+vQ7zPJvorOoJaSXzQucZIIOZpJnOTP52TC746+IB1Wc3s/A3yqvzNcCnif9SLPvC
zDqYOQJ8qu3KOtSIlF1FGtHn/2wHSYzF3vKuwNcb2EyIQTjfplJxcxVM72bXk4LyUTCLW5LDIhAB
VpZvnxvdF+utAeFgSNka6Kgx4YeGk2NGSrJNUVOq4fqz3gTTZMsK8LTgIUXM59ZY7PfJTRGHIqGB
2b9LriVjN1RbGi01ol3aotZ+Dx8LRBM/FhPJdLkP+GmxEvE7bvTGfJgrsLamqwqTyHnXCCR0/xgM
buFkjbxpzP0OReDmF7CKQ5gebR2CejpvdmY1D3X7eaqspTpRxRgKRZqHbTzRWuyej2X7R3vFiRG/
PH50kmSTajNMntpsA2/93s6eA2SPMvINrEpx3D/BHlwALUZZWAQTFsYG2/abTSkWZ17aIl8IsgjZ
JBBUqg74RI/THKzVFXIhNsynpXJ7rIWRRxWFWoedf/1y+KCiWUtC1Y9g/XQMpmuxhpu/mP3+RJ79
ePDufgCSuSKvtzr8parvHp7TRC8lwKA1tnPvJDFAHSk2Vt5rpsAbaeWopVq3titA9fO5iQpLHEJV
yOUqBcT1aIA3yqGHxFlMPVECe/mwf3WWMleTW+rIHNRNBJ3A+BkIzH+QYMx4YSPnPCbkK6Fzrlyk
St24SRunV8PO86tF0RQouXJeYyXhyi3JwGDL5Qo2zMADU2m+mFAdrq3zSdpOOtcxtEIHBaPQTdcE
W+v56N9yaIUb05qX6ia0hscmXCy9Sc3LiIAqcxwNIBrh6yPL9ZqzzMrFbcLblv+Lkr9sweNdkEPj
d9lNAxZ/nWD1MKrHjpzHKLY6G3SVm8Gppu873mCKrsheKTaLi1sYBE4bSXtuD5l0twfrYJdrokvs
/Hya0X+Ar52D45Wbjw9yNM0v4NSpu/7PcVnuvD3E5nA7PnvvdK0DAEM3rwte/y9UA4o1HHqk4VzG
d0a8aPRuE4xHvNNeiZqIud7LUC0F3uzlGaCu502SE5wkV6gvemiTwpB3AZFVmqLy3VAB3G1queft
4qeRD5EC2PQWRU0P0qUdZ7DMA8AD+oqlEVA65VqUC9AYxQD9/lP2FFBRzUlBM+fMn7iHX0qoPPv9
FqM9vObvwh/BuFzClPkFCilrnLMx1mIHkfZclsrfVmw7aXuFWD1IasYoiigijLOgWP6/5aGD/bLl
M4v76bfE8rrE/QY69ac9AeumeuwY2d5ooiyEn55iDZZ5aihAOOho16eCkkV8y0wkf2yBia1slG/6
IFSyPo4Ya8WBOQ00WwkR5Lkfvhhow1w3vo/md331T/wLnZf4qgJnSRGZx/YPNEl8BOgmUi9gJe8U
8pGTmun09G+9mvbyakD1hoPd5CywywHqtT6Ggo21UNEivVJmjDV+y0WSZLiIDKkuJC3i7UKBLZ8m
FIWMxSv85BvtDrsUutuFVXzLHFgtxzhv4+j53WRHEGtEwCnWTFuJaTA6ITKe6cfRhfRpR0OKjT95
mwfs12WwDiweTZayceW2nkEVcZCOckNuC24HIt6DBF/KSj3BVfEa8JHYusu5HEGqPlvbD+SxcLf1
WwoHlIcaY4iwTX0S0CcRX0JEjVCtiFftftUJYuaD7sdgSaxNDn9wzaVBSvwA56hupLBKw36OzqEh
/2ckrW2rAEj3CHp4INChQVedd+5uPBB2I49eZY9tS21YSISLCzPtWjoPkkcu1hFSOtVnkYBd3LvQ
HHozj6v6miSE98YnMsy6Bxsaj7wgIh5m8+yv5vdNS4J2tGW8PgT5DEYI2OQiCT5U/pbOwwVDyYPg
Ydx2D2xUbO+VHqRAXPN84icVr2dDtAFPTU9EKQxh2CARruh4znTqEKqMd6OM1j27Uk3E51FDzwfj
dy3vmSW+Ek0odLNSnc5eiVdFK75kRC7DeXUH3YomOXoIxEBhzkOKd3hvJuQAVQ06JYW+AtUdxWCx
jBtWKhOwg29S5AgZmTFGg+1qtpa4csJy5TM6mdYyL/NAnPoa71QJ4cMJbwSHufsqAKUZyOUZmp2N
A2DJIRcJO9IQ/4oKf0GdRrsiGpEhatYeAVoPlySdbIB70ek4IseQjQet3BsDP3d7u3QqiGdBDhPm
vdMyGHMzKN36hV+HTTYWvhjVm/RrV7sJ2McCj/SH9RBcMkSChZNKelL12Pg91oT5qNeYoU4t99Iz
XfWk2Y+O/IQtNMtyU9tuMYPiPZsQGUpzN5bsN245LI27AtQ5Pv9ttCyM5lVL3+JBEQwQzsSU+M5J
RWNA2qDS5nopZ39tWq/FEO0ebIiS0bJrH8GHCOdt810wycDBK6uXuVOZRHUlyw2yZeaPAEykYu26
W0v34WTjCXD6tZuGvR18+I6wxxhzxQMQdozo2alirbk3qijeqk1xbWd22h6Pl+ucoSr5HhY0ODV+
RGGxRfukb+SGcv5n7/9wDNy+e7PDzUJ+Ma19Jli+mKM1jS35tWtfjtH7CaEpejjKG8tYWsythJSo
OhhZlAXxk2TFQEx15+3FhkxCn8nctnuCK4/gMhMIyCX49JCXs2io/pAr2mEGJFsjPKVem84tqdEc
f62HoVu+3Rsae8GXpRXRLSQLoh+r6ufxJuFnzcroFQ/GG+LGGQpEF4St6Beeki2gWsbjkInxHtZe
YFLOcb/lZvCosKP2cS2nRIw2vO/w/u+sZyL+8s6DuLbRbSAzKiq4RmGcxIqqsEBiofiBe4v98Emd
RWCwBN4Oc1sq9zAXP4DMyejamheac5zy0j+wom3kJS0QlcePtrvr5jr5leWUgTbj47rpaTzTqgfS
vzBqDJI8Jo/otG7a3ch0VsGfPHB0XjkQByG5lpFakYOCa9cXMRBa1uG/4B9xxkewtug27FfVZfgR
L+VI9PEeRktjzgpnX+V/+AESp1sxF9lIjCDGGtMjWLdGHtdDAkcef907a+18/8zO71sMNgEU02Ha
Q7Hy4R8MSPNwrFiu5QlPJXSF+fMlmH9RCi6z00Wun2MsiWOQNyt2hQnRkIDLZeO+vqAeFkoI0x90
SeWJSJYanf45ppL0s+8+bZkB2SvV419+cjRyd9/HQxOp9V9vu3tyyinR7xVEomdjMo78rX+x+FZ1
KPJ8PO8YaRX23NMOaMMyVOLawv01lyOKDCS3BNYt+9ahiNisiM95JKQ7Ce38pX1AOSete4Li45L6
8lg4AZxiCv8wXad36wm4SUpW0qKOWUOA105bQx4m6cMN2A/GPFNGckOZju6FkT/urFK8B+SUkA6v
KNN3vS0zgCTwdc5ZZqc9LZv/1cWG6ISDsVE4qipYmHgvXvxydA/d9z1KQntCEOzOtnirf8l0pY/N
z3u8msu7W1BT5XqgCzgnfrbBZJm2FdpZEgXLy3qTO3cdf40OInthGwpydmpYP74X+k1svJx1PrVU
g/Ft7tD3BfCOOQUv+ctiKwH5B5FtAqV5ESTNpAB06SCVPSNesNLsY3R4VqEUh/cWKMhLTqq4QoXI
uhau8nRW7uJ/dWRS1Rht79AGv4tilm2Luye0zaYD4qt2BsSLi+YPaT1VKW80qY55APxQGQVm0iId
sMdDGG4L82oJYbzAsaWweVE0dOrvCVAQpp6Bq9zC+S6NAK1nW4yHC/UrEBJV8+DGhVieZMnfzmDY
v6yb5GecIQC8ZIfM4wefPuGuDUx9/OL4S+wZApTlTvgoB4VnbpIfiBPcBbuvoBaxLBdjvOqf08Ve
0hKIJQ7INx8XPCOlsT87tpPqdhlkFbZZ0b2H8FBzlfz1dYXyk1pErgCwCrW4YRJpP5JAXGHf3lK1
rnP+2sBvjmjgNwPZK+Wqf+jQ0+5/xzDoMV4ZE3CFNo7oXEnjDZxHFu6eT2eGIJkiwzXuuoSI1T3t
PWvLqP1AycvgH7XWW+6sTz+ezuuJCXdRLovjGoGfVUgmKgDWISvXM0sb5LPpLWiOtghkjsD9IpRI
yaolaIhXEEfVo2V5WhxKL3HO9JC8fANDANAIvaggCRowB0GEtIkYQ2DEUBtlooB7uwEjXsdOmZw8
P9CczfUv0fNthKwZJJlYhu87Buhd+baNfCxM12433LnY5EJfSj/xQw1/N0Cf1CWIe7R7Xau42V1I
VQYn7Bhkm/BF2sWxM4+0Fk+FPEZE5PrNsDarnMpfsOoKXcIgaCPdu9o7mLAAoyJh5rQShwX57Y/S
67Cv3idNOeQIAgM19E1V1QzU6IBZtGunagArdLOQyf1h5dTqtqwqjn2q00R1MtRpcr5GAyuJnaXI
OmROStVnzz8Fb3KMWdl3zLh99MsvTjMz/JlVfKsRNCiD2lybfxxcbcSpQDy/iMhIQXKZ+6Z0x4HL
VHu1RKxKlUHZurpSSd0EXjaYasROK61VMbRmv4SDXbrctOD2roUmPJS3VYEHN8OyNuknMP8fF6x0
D6AubiQf8jU9hj1qruH1uMe25G1DjyPzZcYysGlEMDMsj1K1AFggAtyY+K7aa7+DDJiLjaVhLnDM
EL5zy8QnpYE8onpwTCa3rk+ITS8x5sdcDj5xiIeAjIEF7lyfjT4godLWD8S/DgDeZwpTpkF3JYUF
l2XTtpAP1XAjAgIl/70i48WqEp4ye2HVqlJB3osHemuwCqqS+4PrZXHqzcYLIpIY/3b/CKx9JkqZ
53aDt/jjxHlG8HH5Z7kEeFiA1jy5/zLoQ1/UYOwIftqmB99VdeanzaBQ7S6GhHW79wXgYCkgETNp
GyDy7yn1dtTCDxS3HzAtne2MSIa0zn5imGUlGvucRV6HofUyZPsPJAC5lqrpyIbb2eRfNEkz7ucU
jtRV6hvNlygO0YYNiUDte9VzfN0GQilFvX2wY2nDv/w1roV9E7S+OkCjEsOaolAPuorCmjsG4N+c
M5D/WQJuHat8SSdQDWhJemfgeYDC1v7F0Hmv2I3RqFdxwYq5VfH3AYhXNgKmSG8hMV450/WHuya8
+vFHqnp44NH387xSsjDvu2EUk8sji7OjTeuCbVJkvzyTF2bxBiakl7yTfbcznHXllJb0IV4IimJg
duRUIm+9nqCrXgiQ2O5BCdO/OnkdZU9W13UFcFHx3Ti9mu/6x6/8M7EwiV9KmfJe1hj0YkFAYMgt
qFO52wpWZA/0B90mi3UE2tbtb5gNAZYIegGOmfhlHir9aYAcv7PUIFte5TNpitUUfgSxLRmckKns
SRfmySRoJFHyw9I+bvXDrnB+zLwKkyqT0jW7yot5J5QJjckOd2/0HuEumr0IgND0WMzT7vU+RGAr
r6QZflST2//98ZvS+IaCR6fh4L8Hal00LnNzlqqe+t071D+oGmwY4IHWpyrYMUg/Zg9tIR3dXafV
7TuZXt9sNEVV4xb7myY2BhhiycwemKaso30uynzKmPQ+SgrAeXZfLVeeue+tE+lIN346BdHYNEeV
gmQfcR7rDCp7kRbVv+W5ySGndeKxvnaYbG3b6Ft0RelZbYJQZsQt8ENggsL20fdoO2nHtNvvmdvz
olBJLuu//Qd9X36T+7ghLhU3lb6V4QLBSn0xbCi2/IgOskbRdb1G2mViN+n8j0wn9/YgvNEsUEXU
8D1CIQqRRQBFCS9gqEUgGdtWZ2HzsVqmBKleatQPYHu77b8fNhK+v6shk2TF8LmkaxkKkfd5VPjh
q7Xlc5ls8Ae3xitFWG1YsGIz8/mbAIJ+eV4fzp8sz+VyuxXdlJ7oMrEnlvI2WxyW0MZ6LQ/pkJmA
D+ztaPyEdZD3Q2w/4bFIs5zS+jQ7iT+GC8nz/C9SubKEhzbSNaD+iVLRliAPhg2mtwM0We1La46V
CQf4LrjJ6NoEumn6uCl4uZEhzUMaO9dwXP9pKU0iml+5TjbohY1GIa7AwNDIWWzYVoEpiQD3Pr1N
XupQgVUN4KnccFX0wlqUtRQx9jEKEeDcXfAeqP+bmrey4azSh/FCWyZ83dTEmdHIExNyXt34a487
gECdyXn4rWzXaTiOjROqF/uX8/9uBXshWnMIs+pXZVohPCC3DgNdECAMqdeLSu5mUw7rvlN60ZvL
JysWSHHTPiPQsMuzKg/6HlDxczBsPgWj+uO/twzFmms0DPwIRiBOLXAsy4uMw6/vb90zEG9iJ+Y0
eT/gezGr6WorQbJJYM0fdQqxWIwNhp/LSIMt5qjZIpaDRhV6VoxMF6wKo+dpx/SzwV4kp20+fVFS
r9VBn2eA6sXTXSwdj1U4k7h5rnF0X68hsX2bIzxPdHiM4uZXS6q4ke/Bf6meWPIfeSxhy4mEanHC
zdjAer/w4CKt+yXLPZp7j/WuFIWnKmmOXKJOF3+yelQ4jOzuMAI2os/IgPjrs6PEnZhp5AzMUrjz
qRphLvkGTobOvMAPoWHfEY28HmBsJBKRS/cTuqWIwBttml/KtkZQKVuR7FhG8rZdRG1sL8wNimzS
6MDrqdaNJHC23ls507pjJLIR0OYTwbgYhpObtUGS6V+8yhZPIuyGEArsa6Tp//UCEOtjMm4umpGD
RDMF7ON5S07n4KKVaDB4M0AiK2/sX6QtUr9gyJdk/O8OStw9uNfwexA+qybPC5ifryJ5qJzM2HAM
CY4r84lYKEy3vfx7O6R27G2L7kqaGqurCzMZEiPHWg6rdBXILB7vJreFV0YjxD5yeetoPik7Gmn4
CqLAuVrT6kQh100R6d2/cj68+zAWuy360LJwWJX6wims0rSxUih7J1M/EzMsr1i34ZpQ78nqpmni
1HowsjdAv1Vdtc8S80OWhQd8xaIP8kSb+AcM52/wHWi8c8p+esYsqW6HmOWPFccfCxDsHmmLLCPl
9t+gUWeaXMhC/jAKqj2xOVmLSlupNPIF+5lHFSEZM2WYAsqH8xiR5LuZEdokZbHoemxC8PIOR6Ds
tCK9OiQMZLrJp+AwR2JKnuo4ERBvRM7pLxKDea46Gq9LEvIDhEfDMo5vNEYX5f018AtBbX4NdzET
1vNDT/bGfYaXouWJws6FXENYf1kk6dEJhMFoLbH1JRVWk0tZbt5//JkRidBGA6yB3cs6FHy7KcwX
TMu5A+ItRmf8jJLCMQOIF+ISh5bp5pplnKobmWOiMZcq+rBSZDF6K2zWvvxxIxumS44I0wc0ICzn
LDzsE11XEDs+qD9HmZaYBsFRj+VOPEAxIJlSK2tbQtYw0nxn74lFSfD0+hTZrXq4VDzUg5j/3ZDN
UUC0IezWcdzILr4CBQ4ozwmTIT/PEtpvyooIGL1+rNEPAG6OWuL5KGQG4XMSpsBum8cRRA8lGAIv
Xp1MPPHMQfkJ6Y7saUyYOI0MoAMS9N3ENtKbCXV3TbhUjvl33LfkSeJeop50uhe0n31kTmtmnVXY
5eWysrSDHqMy0lAFc3aGs5Uyz490XZIQmR+zQC2eIb2I10mPB6qxLLv/bOVpfz4gmPYCEzrXmSr0
rJYb4H2fAPr1CVI4xMqHPWsCOxx/0PdVJQRtfUROTO7PBtoJ1qJYWx9bHU2At5Vo9PbQjfF/Llod
DUt2iJYSSmgNZ3IPURgM5tnfUX3GZ14mt26vWputKbZmecDRFhGkHo+vt0XAK/AeDLLJdN8Foxfx
igjD9XuA35w3qsEgtbo3AHR0ud9Jy5O4oxPAiKw070f2z8j+Y5y8jwD/hGwrB1e8ojnBWZGVcB+B
La22DSUl5R+F/nQu+GnC01QHJksEeauN8YXFKgy+LdNUzwIROH/OY5/+sK0rA5SaRoVAxLjzxGAq
N55+dY5dV/QlEW9th8hZQQBepnUqcwx3D2LbTD4jjbVZZ67YMbR34mUJrtiryj7Bfcssk0fQqdIc
uB3mrwxXQ8mmqzCFvBiFOJKefJ4OhkoqJnYT6KOBhYUO8Ni1Ouf0ZQozYD/vOFAageq6wsDcw6Q8
UFwpKLfac2O31borj/GFF3jg3UFb+mnjNQjhSpt+B6yOylZM+9Qg3YJrTPhGiee0mknlrg2lE/Tc
ATxrwNSjwcZ184X+IJxU5/MX7aULKygYxJibFEmD18ahxmuxBU1WJY3zKvYH7EDV6UrSWZxept8f
jslFgIkdMnZ0akCy9HQudCrYMbU6YudkgoLW3/F7QYfKKZ0P0nJlG3YMSynz8osf6nHTZeuldUOz
29Hzwjx7HOClolEVLRhhfe46aB6yQIoFpSddRe/xOSjmTUoxShZRHkGXy+phpe33NZwUYbnFstrH
S1DJFpkqARbFJq32HlnaLVZMOorEQ9yudSVNoUDyNgaDHqyvah/oPZINhLI5okbP6rl/OvaKAfQF
lFeBodxf14FnzHmBMguktIJIy/0qi+1JcB+AZGAGY7aHUBbaBHVfoZwNYkxLGstaIcru47edHVdz
KpV3zqsa8SLvYsW+3WTCl1rGEe83y2ZjhC8Bek7I5E+FhuR6b/GOjeKk6XeWpO1uXocZ/ma/CLXx
3zTX26bHJsY5p2X5/uM6Bch6IdwVMICtW1J94uTnzjG0M23rXscAFGG46zSgbh0rOjaRwYu3/SwZ
mYgjvCQkn0vT0SWAGMjsHOBNQt5Br/GIjr9bYPLV0iMytEBmLSom7FMjK/tWDJJcUu5it8RqHO8z
TK0SdGIegEt9kIgTZ2DNIJdSxkE3OvR7g6NNgPb8stRftML3vL0vTqX/VwA2Qcna1T1A/vJCHd9V
QNRiLeX3erqR0MvZ1YHemglGrEkxhgbnk6oi00uh8+/bgdBf0tYwgMZdTYIfCZYQ0sCzouVIAgRL
dwZ1lyJNYY5cJ9ruWkibj0i8EGiDavLdRkxslKWm3i6Gz0lpiGiIDei3nD7zAk8OJmzZdO6NcbVJ
FIWQUhNM5zdlRFHK/i+k7tCuQxcOD18e/yB7IMggRN8o3Q0bQbC8C62O2wBGL6A9PM25sV+Okend
Wf+u3ho2puBRy/eaI46E4k4UaqUgloOzJv0JfpZKZaq4662hH7a1fv1ySNmIZYA6eTSQbwjPV0qQ
2pUO0VFW4m/S3ewDvNrXkNJb5T2v1GYo/N4yo67b0gSZOFM0YYezefhXx9uMoTi38QEw4TM2W3LS
yCgkz8XH9FVDccIMa6MEuLopyOxA8eO3fu8jrTFTecwmajo8GpNwK84cGmykOg+s3VSRu27zur/7
PIAsBHxToDibOFRgZK4Ue8bfQ2UaVZYBR8B2aVJTNA3IVfFQoGRFaEjGupSP+3XIX+2j2ApDI1Pt
Q2yEDoPUJJBSwkk7IGvr1/QmddQFDkinTsG+erJJpHFPNRXU+sCR4msTQ/OQyEEWMnJrMFGUTnLj
8zg/hJFuWUuNQB2V1SFyYM1isS2EnArWnBVDTyjS5HNVMGDh19+g9l054vxb1Le1/fibsv9U4EXt
oSv9wUAYa4S3wrAbU90XC0H8dblykN+89BGdyaAYWT3Tr9JMHxiQr0ISwZlhPU5RBvINE3v5gd+Q
Tekfp1pcDswUkfw2PUmSHgM7JRTf4koMJP4FaSJwXBE/T0yow0JuGqeWlJ+95ntij4biajDfUEvS
TFC0pzC8vaqesBpMi9lTfbxcr2vW+Rkn0abO0Va9uee/M1iX0f1CWxXSvQSHm7vQwrSFKkqxfly0
iR2bG3BGmS0lL9ffcMjQIcfxvUa0+bRfRLfe4nu14LVm59UvTzaQDIomDkQaBY9t5ZZuXgW2HbIb
lSKZJWyQm+kYdsJBhHR/fphCtW5f/tRIA7hEUfDLcT/Wc+lS1scA3xoN97zPxp611nURm+FdIaWX
ZUc2YvHO97IhEupdypTLlj30UrrEGNByXptG23mnWOxfhhmdro0t+sFm3K9cr3YG9Iq9tfFh0VZG
N76ipPp2nknOqqu1adsjJqYgBAMxVfi2O41uZ3YRf0vGHydAxzXokdZz3CE19gsSgCcMVA+h20Zm
McHdKpzaH1iJHaDyRxMpSM6TZvby5naRFBEhS7zpWjTSGEDCfpIkulYT/tIv5f4pH/6RcRxunBgL
fvHh7Znsih0IBNE0Shg7zOE3bc5gbONeky0GIQ2fUnBFb8yao8YH6gEdsSbLy/a/8XrvnML6pDjO
Zxo0oJx/xb/jVJNeVMu0m9Od2nxD6W/o1grl10Me6+TcpZMLJBteRbO1YqAWulWH4tYQ2Kb14QyZ
kBfjkjqwz/KM36rqJBybrZU76HSNHE2Pao6pehAdRpFDHZkCZjVknp4hcHWmwUWHl7VHKIY72oO1
ILgXDdzFY7fXul9akGLLNNEY10g/DuWmitIYRTikqTgU+7EwjCtZnOgmdJnQ079tw00gp621MEVp
ZyPTMMQnG3IUBChdWcRAvg6uHhyt6dfgLnfjt/iXF5XR1fqY8USqYCPnaoecHHBkQcCQOXCdZnke
ivQ8oah3bgMLMZmpHI43SMXRU0Fmcu5EOvaANFcGZETVwdGeyO1fa3bbKCcsahMTFd5RlYf18FuC
uynuKaXBXKitzOxptcYu3IH4h3jJTPM7ZuLr1NxydAKRq3JUPXKNn6ih/dbFHFBRJoalkQFu0Q3o
CV9lafb97Rert1wieMSJ8dsybTP4xhvdpVgb4v97nqBeS5bdenn9CzM1lV6hCIoA4kviE/kFl6wk
NT1e1g+ojEgGdT1yPp0y0uTrMkCV3sSPMg2/BRoOv37NTVLDkhIATh+Thwhp7R2TymgPolu4J3Fo
QziBDYySFhLrwN9ps1hbHRt8TUYdEYj7Fz3Kgb0RSBO1qFEJ10gnjfAMcnDTicPigETdoCEOJU17
PBPgP8umMhGSzxZhij2Y4SjkqovVjqVKCIgdMKQfSOt7BFL7cQyJSxupOQs4WAzg4xDbUWCfCeC0
X4owMhJYvgDTTkIjMB4+Ow16oP+D1lGTn/odvvs6pMPg1X/7fB24mbwPQ+luVrId2m487eVjRJbR
oZxZuIdNLiYEAYDb2nI5S+WeK1YHLjGDlPvYXJ293qkSk2I0VTZdMR5PIk7PsM8lL3HuSZAB9F1Z
sbDulD9vBrrH4KpxKDoJ1+52LfzEfdaoMC6dc8Jxp/au0zGi/XiH/QjdhecGGueICNqfWL8a/hZ5
IKvBCGWYOzXw508GxxgH0sQTuZqbWW85zuBbd1h3LrE+RRVUW6BV0CxYjZak1w/Pw+eNnw17ZdFe
F3KVsdnZhKkKbKXhJXt/8TJrlpKOebyevaPSWnaBWAXRPG7kTQpb0BoFVSP8SJt/CnlkhGAEdc1s
e/cUmYFGyiwy7HEyFQczhC52+qzZSrrZ3us9I8SuFSeKSc7oWUUKVPqEWtAs5i6JjdjoawlITFL7
+GshDAPRJTxbyibcKJF0yqvGGeCrkVSXwt1wyb1kEvEEJ0l9EG5xSpdlrzmBjWGK0o7AvgSNqKfE
+Pdv9AUiF+Wcx7wods6+cNOzIKFnthDjKT1Sp1TdHo7AN59k3n2pMQz7LzAQsjfyuO4Pes0sgcYJ
cH+ZIJ+M7/bPa2Bz4XKBI9D7nhE8G6qEsgRj6yTByr4Z0q3GrdDlLlETuaST9QN4u3c6mmlxk0KF
6ArthatKWxu6QADQ15U0PVOS7kVvhlcULb4Lsb+WYx6ve/i2iauLPuD+zIY7L+GTKBBkUtupZEjN
SecnoZe0KIzuUvHMm2LsVhyA7408XZIPjnZHi6tiU/3IdvosSEHSzZecAD05zLiti03p3ymm+O79
3f2nUWz9AZiNEkvojUcy0VIuW5D3FBWzdOV48oV+RFhZRQseqZD7bcBSSpLBK2Ia5XkaIw1ajWsS
FL+ONruvlLZEWBy4el3xmq75OtIBcBlzTYDnLX3sz0P08SbuwUR3HUgV511Pwp/ZzJ9PaUoXc5DF
hAzn2Ty3otBoGM/SISLz61lDVWdCqroLwYlCtnPaYJQuxow8+yhzJ/9Y4PsBdfSxeVYpVUh0/mDj
zv44H5+hZsIO1zOhABAnmJv7mtaZy7TyOP3Y3nuLJMSRJPunKCX4drwUrd38/b/FJKVslDtQUL22
2cq9wEOQA2sSWSpdvO7Wg/E4mNiiokGy7LCectvV4WUEHQ+Fp7f/+FcwVD0fpjGnJXEye4Jgohkt
o1Shwjg79LWyMo2qQEOtojPW6wa9izQOKBtL5Hrkw+dMudgf5JCyw5xEj9/sv9yEyBPLDLMFe/zJ
ALr/O5kJFPTP5YzLbl1nr560HQaQK0ZeCCLk9rY7dTrTYGIxxhSozU2aJnXpRxROvFDiWRaqUh0p
DrKfeVYcGRHki7eSktCD2SYDVMKd/79KAnEgOL/cHks39h2P+FrgkOGv/a2ItlVax8sXXZqZ/2se
g0kw++/5QRcOxmSo5XUL5OaVSOjQaWOUOm6URjTTVj0h0Md9JsO/7Ft7Uz61+V19S06Y+71BSJqG
8QnHCClSMmOg/nEfcxnP8q6iMnInVKnF1c7FTZw8aNg7Dox2GuxE3K1XzzxkdUAsTX6k3LP31ib4
8N+AhhFWbe0TDJr8R9fut55BW8q7oW5ubFJXHcNJ9lXHs7yp92cB/TZvtXpBZuf/SkYphBVFp8Zz
vgjOZEXXJPRIbwcskoS7/cB3M5HHjrvJ/cW92WjhgPfx77MPV/ETIpxuREEI0rGt/uqeUOWO60+T
E33Ywob9iQBTWLU/06Q0b63/5IwNdcIz3XGQ4j5tGKcnsyAlNG5VkXRwhhJd2++64JXaSQlSMSEh
nV+BCHcH6nVOzqRG7byle67K+rsKZtbmpuy4piM5E3wSEkXLcOIeurHMXet5u4qShm4cLO3FhyZq
os/w6SyzmRiCo2ziplxFDAjIv0x6dxXh5ih6cd1vcC8X51w3p4JjQHwOFUVI9dofxFzzVaadA+Nv
xd5LI8JREfQ5i05EIE6vPgIFiVcQx2mfHDP75Vx3esTIFq0IM5iGS+Q2QKmQoVYR1XcGPpoSMiAW
0OpW1zWxJPUo5JIythrjY1yUHtMFEnDEn8TKExQ7pEYwrxgzO9SFjvLDlRLKPpXjPzJZrbsflFIT
1E2YNKEm7HCzjFoTWaS96JOtBf1fhnrLruOrrVwz1ia6c/Tf6MczQCgrXabaPCnUuuLBgPsRTRzg
5WlZHMu7KXX801K2NuKDCoWldpgVZcz90zpHxRAu27R39qizRZcg9w+qDFq9SmPY+4kPRLB3wGrJ
IiO2xvxDkIIaXnGpLv36ukqYvQdBFeXIlQFqEtWUI99xFvieTDUl102RARqohqbWl2lDwWmQnlzK
Jd2mnDDyE6fOwbugIqF1JHOlycc8waENbs/ln7uJHS6H/oDuaqyua0kLHj/7ZUEXRZWv2yjMUHyu
96PvdZS8qWfqb/mHNRZqvwQ+4hHTIdfi/oq3WlXTm9ZvKlObNFyqau2JfmA0DfRde0cgi86n7HxM
aHyjS2Zvx7B/cCCofaaTQTyZXD7/MkkPXa6w5/3wjUUiznvNeRadTlPO5tkFlZVTAY/E1ulDguqh
16lJeiqdA/yiw1NbQEgYiE/tK850WOr/tqZyr0F5DZ/MqkwtCzpVeom3psaz3UPrVWU1SqMb8cdX
2Pg7MeMKWIHSn1Yt5fmDSN7/jDkuZhPLYC5TdZrz4b27o37GQmFFTCraCE9Wf/sGk6QYxXYV8STQ
CgRmgqIOWyWrgntfPxbfEBlNpQYQc24AcoVlJrEbnXBStn4WszXmN4mTHEvvGqbdNodavgYFZVWL
RBm8MXMOuWLe2WwPcwSnwdRLaNoBPKmbQxmR0qLCAj5MAZjBCBwCizvdGel+17VfBM7Rx9lwrDSn
pr1qzzjOVLAiVuXyF0599JBtg7uXS5pwNXhKfMKC5duhNMbU7GJWqYTxLoEazvjNDPJ6HIf+dr+5
qt12BKGKvPa5nGUQFa+3r0uClswwGMP5gRfKDr2c5JzqOhlmOIZSqzd3IjIKrqWCTIDY39bqvb+5
XUTCkvKp+gowtvmgm6wsD1dAqqdhVHbr+lhl7SkBICGJ5Vslypfs02ZfWL42ETbU4pmbDeDnDdaS
N5TDK4j0MwFXzgVjrng9yFnas6rGE5ECV3kTYkgXb0T8h9Y81C8uQAx/r4YXupOWfkBCKDH271lD
8AGrWbDdagX7uM/DA6TK2fBaTna+8KxMBHU14Hu97QlLSY+ctJ7yFszKoJuRVQmUxiViXzff+YYY
zMGDdMUT9U4cd5tWxLQbGcVt7GcrUloyMV/Lec1PuhTxy0s9DM6yvvRGxHH7nhxPzaBHf+QpFV6B
42Q/LIRi39MyF+cAdHtBDHUeAUgBzw2hj6xmyG7KoxDO2zJm9aeny80ANPj3vtLgHRjmp31v6SmL
sQeyTW+IsMDcivob242ijiAOV4M8JIu0Y/2celZOOj/tA25DisKZkCtyex2EeXvMkW+rxAJ0obTH
IzybxmpjxZUzP4hn/Ni7R3II2llyXv+GSarTR9XI7rgkMbCGmXPMYOi7Apt/GOy1svNX9yWMT8AM
znMcrM9L1Q42JB3H9F+P7p9NWPv0YGNw/7DUxMZzivJ6GIp2mXF8j51cgtjPeb9Ebyn5JykdyqSh
2ZVLiCrNTL82qHs6V5q0kNoAmnNl2wV3wyEK5je2g5SPrJRsyB4JoqKQRAnbE1LhRRwhwi1Ds5Hr
xcZBCpq3sTngEaLGyM7PM3RgPXEkFICLLBevhuT+yItqc65AXeZuLkInIW2POpCnRpr2ukPCkiQd
Ad3RoPSbuQF0nT+/+o7a7FYYc0kctGa+54V4driTHRtGX68wywv6ElCkBCHIeCv01iTUASb2y7tp
6H33d4gCBGJx8OzxO4WTPAzApzFZTIsAPMsdyLJkTio6rzWGZHCP5UoeAT9Hpz+O6xqkrjmPmrhr
AuIhvcTyWp6yfkYXcC0Wpp3nSQM1dpEJDGTKfIRb+sKzq1MNk92wgHy1iPNHBGYzeYai8fBlb/lN
NeSSOFKYTyOT+/x0xfChDqg83J6/J6RJcfegf1JKDSZLu/h2UY77/LLtmkcHPHmLjUa21eii44sk
dQoy82m1NGnMwGsz0RECnPiKAFU4wCKAU7YL1sGdn7VqmVp5AyXaVDUf1nlOvw5PIpQ0txwFC8nr
YWQSKHNkrq+ULK2jzPQ1vKS9WF4BX6CX8TP04B7eRw+kOmuiByWgF9gjTpkVl0NRzlsOT0Dfz8qw
gZ/jgNRxUf97IgGtc2DmyWEr4WTEQLqQAEZddMLVFPacTHhW6mJa2/eswZ6JceiKeBj7iFsD1vEP
MyPAhIJO2zUAi9FciBjIz2ojmp7y/AsFTyBk6nvLv/pi7n505v0dKlIav9cSJYyjNQfJb5Ga2eEC
UgWjacl4E8NQXAAY5dZQ57dulBIMRTUm4oOHhAEdjLOmyuEZNlxjw8hZOarTRPNewS6Q9LVBbPTk
c1aGz9vsP5ZZgLDMtuc7k1YixR1Vzuh37qlAIHLFj4oovvmDfGIYPj87jPMeBSmZfJwtMeHCYrso
3G4KjKC9gQXIU2xaMs+H7Uh6tBPiuMzF/MbIIdcaDPOTon+hqH6XyjgQ9FC2AsObyR3dRtYwFTc4
3FVJAJw+bPIY4Zrfq/IkD7v82tRwWDE14RrUlDQ5Jf6foD5VKNHgj4I1MWHkZs5321QkySuFRS2q
zTd6viZ5K+U4dgTtqdSVJkGHz3icpOVrioGBJC8YXur3TPNamN2oAsFMm6rFXT2M5rHGY7IZlrW9
HK7ZHnzrC0+FQ866cV7Yk3M7n7+gNLWl31SOQ6vVOzLzEHFSrqoloKPo3cfDQxnINMyVpuJD1+Gw
tLoM8zfKTp0avVJFVxU20NvzKapjbiGnQJl/CzDW334O03UsYO1Bv1aZNpC1mlPSiMLiHLCFHmuY
EfxuHq53UYNjcPDbUzqfxKC2ML/5zs252nZ4hy6N4ma3TvFFm5Suxrzu1ICHRpPxYRv8DEy1xjgq
/bm78T9eFtuqWj9oDqJlmgViG3tJKeYLUGStMfLloeUgL2wXfz0/HtTpibgyzw/qdgPs5YLJcjsl
xTSAW2VKhCS5SUVaX2IoSo1BvTMdieSZU1BvTO9A7TtoDOKXSMmTkrvRYyscCimk3uAA886kZKG3
YMqD450p6790knydd5a1earieUU94p5/clB8bRVO0MiT2zB68Wsw99j0D38v2dazjSt+euQ2tsxe
W5Ij7L1KTSM/w3k+2saiXitj9SkwH+drbLqYyxssjVeTxzK8X3E4jJ2A60jNapNZIr81bGvnviVo
+00pfklGxPlQD4Cx22KNYyGMRJ+19cL7EWZjdNFE/C8S3iF41B1F2/XRoMqdAehjXG6ecf4T+pBa
VIpcXO25PFLos/mqTa22qYvmXU4MhfEUzgyp9tPzj3vG7CZ+Hr848ItPrQbBuu01Xg43+k2NdHgJ
RMUONI4IpssxitFGMDqhtBwtG4lETitbUzg4vulArc04he3l+E+yRY4FHbZQTD/pNkxVqgBlkHYS
AAzwC+AANr081uxJ0b476uh225DLkwyBUxwVOERT1m1HFACj4iynES7/KVvQBXQ4Y/hpi17/PsFJ
gu11mZ5jvCb/wKvs+5xVdQymzIB+L6W7Waq19KlJDa/lGSRI5xaCV6taR5QgGHsyANtKm30yywC6
OhKgjciLhU5VyZd8G4b2ujaRvke2/LAz0sAYFc7SSp7y0V7oP6w0HYNBXUy/u5eFKYvh7wRO0tuo
Dr0Upn5MvkJtRuX5Bg3Lgtnwv+QzCxzoHGISrz58e3g5oC1GWzBs+wJN2uDDjWASPuucV3vT5+29
8yFQsttGTHcEbV16j0Lz0gMeqqxsGQ0aHZEa8UAxAAqQyUraXG5ZnlVJ9F3I61xlfh2lAa84V0YW
4lVnWCIkWIpXQTW9mBBjeJfcPJmWKF4pnpqEKs+1W+Ro8l29u4ZvV/2fzQruOxty7G3R/YpaF+sr
wONf6uzu7s8dTb8tW71Gf/WANOeVnN5I/brKFD30AiAsDGHcBJZ7lc9XvIkswC2s8O1aOattmuU4
WUhIAk3r1QF1U3y6CO784aCVhDEylU+m2EfAFNONG4BMQ1D13w6AjHj0ttszYI5nOx1dlL7ZUZu3
mco4C3uAKmKCH2FEBkLcoceBLA8J6EBZnxApMNjMk7KpGKrGNAXxia1630wn7TZua6D2cifuIsJC
sd+ch/CCsKpqKz1ee7qmy0jm7HWVvNShL5BhdVuFrjD3MQAu950fA0sSNR5dS88wyj+Z1Udf5bKG
HjOs0T1I4qPYlLBJufXckV/R+wOqVCH67JMXFgflN9Fk9ANwYlJRp1K8ZQtEBtsxS9oUm8Pn+DgV
ZhQLsl6ewo5ZAxPddBK5xau4NUiYQGf8tQ8+gZunxhZvUbA+yHoZ2YdTiJzd3FORsBgrFX2RXAcb
WeXmL+a/PF1ZOoj+/HAOD/2vFEAfMefZDQss48RLUdd0S4wIX7LRQjl1zCrekhlKrPowQx7J6nWh
jba7avqkjKBcdiDq7nBSO4CYhqN+ipThTV7FbcOcF2gGO+623xdERmaPxlWCZZ4e3NmiQdy3lIYw
RQWqDwMve++7j8B+MO0CWcKt+SfBzeQO+qveQMxf9fmcUXEblwHrqAgoybF8/nFW82Sk8ifbj4SA
vB0jbROyCuGgJJhzllqGYr7/NGwXYxQO5nkvnoPjp3EEOvKwl2pm8E2A+kgIoi9gSKP/98MY8G6C
oDnO6QRqE7pQhGkZjdR17otN7uKTwisufpmqFcuaDKig+kZKPQxXloJwBh4/h2fT17bnMN03ogk0
keAbIPRDYs7Z1J/5hIoP2fh7RQLCrHsYA/sl1drGtFM3jozKydEyqs6AJJKVsYnsMFEiSZd5Nc/u
b9BlYZ8c+5rPPV2dHmy9QNznuSJfKkyzOeTfsgBhLdieh9KqRlSyvyCgPagxs4UwhTz1yUqJDp6D
pp5gaGGMp/oNPt05lkXxMR6bLULYx+av0tPkvPs8UbntR8c5q0ZxUzLAWaz3icbl2+YXSv+SUexB
DTm6YrbigYmNiaC3XyyrTGyGWrzwUDZyQqNQcXnOvP2Qfi+qqlwmxFLUPn7wAJcAHODIXz8JigHi
R49B1RUEg+G7pw7b4jd4ts3W1rmvNHw7A5SbN02kM5ujzUfuGqwJNI9WUjdhBKAqqdpSpLbR4VaV
p7kTOu8tCyJ+zVIrj67W76CZMwu0ihLai3qDaHAd63IQfHkOr2LYoxmk0S1dyuTJICl0ouPzmoTL
9Eiwrqc3VRVlY8KSbor0TJq8Cr67mjcHHFAZDoCNMhDF1HB9RQ3go922ai/K3uQrc4lL7YQ25kU0
KtHuaFOFd5A3owGME9mzomTV4+PK8gjKLNPlXrPbn44YPQpSY4nH7h6DX7JG/VBK9wlvP+Rjw9w8
3I5Ar/w+e28gEF4pH8BrupCOCVJLDG3R9bHv9vdO8tsD85nashDLPm2ux0ZLLoDCrpzdHjg4WaS5
SVk0etH5tAgVYgMit4/c/YJtpXP7UWGDHhkokSX9PMDMImZvld96NMIZQKz1T3QcBVHP4htF5Qww
WUAc5d80EecLjztwbjtJFBq+95lUsSeDHgMkDYRFmJlQz1Igi3SWUlu6olfRo1tzCj2ngA4GoPm8
PP1yzVu/LTyCA4twNPEj2I54wfPdGmEpbIoeO4gwyY0zv36rP1T/BnIC6InW4Vq81uxKqSQJ8ET7
Al9XSpNkUxkJSoXSu5PSTzntL/MlCjpaN5X+7RUAhZl7pIx1FWHmpHVyRC2s/jS0YoxMjY5smlYr
jvhGbvfV2wzpP6127ZrQY5pcjLQqPyLd6hTknqxXVdBcLvUG85veyG7f7YKLVIJ2ypL0vGJhY3/1
mD6tX8tEBAcC+h5fLIoU3p5uO+qRFbszdFR5IWLoJd+DpaYpgRBQLyIKndfU+266asXgW589OqNY
E4se9v6+cGwall45beMMgferRb+A3aHwB3CptuVqb9iGR8x5ZVOPez0XqZ5ZJfLXsByvihbgiE1h
LwjlUUCdfXcW8urDU/WjMSnnshu/hah4+NXqWE0tKvFGlKloh7Bcma4C2i9Ff6Jlqvc/lh2ovlCt
Jrzw19KXNl37Ifqt5iViVWqEcjODAsT9nEcbMRQRh3xqHFhdjbTVFEUStCynB3GU4Epu3ycNDsp1
KmegSwOAmfl2dyp5geiA561VGYU6KYi0UPaZnjq0R28ZsIiuJyOvk19hOqU+59JiOVs7Aq6YQgPr
SttG+06rxElyvRf61x6dKiF5DqO2EsthE1ltnZA8rhPSiGjlX4a1T36535jOit1HKWAOfzaCYnPm
T/PMgk8aicY4I3iKc/b+sVTHP4+Et5+FyErfL1/lkw9jMzZ4dZA+XAsHOsNxvEXlSTYvrj1Qiojc
l6CRWNjLB+FKP4ZoL8e/nc5iKk0Bjlj9P00Yx7PP7/GBLkBfVS/6a6lbpjxD4VQeV3rEhCCIbIBE
PnjxJg64KeZGn/+aTZ+TBdHg574czCvFCbZteRFD+LHNcy6uQDe1Y/KQ+2bvL8xTybnRBKoR1Y9m
BxW+3UyI/N/EdnDJBK2QpnjEWU1rkee0ZYGnzyj/4dRpW9wg2dyuUqaalQF25M/aenkT4Or/4+Js
sfYd0VDEMF5gpX+71+GZVxAGZYfsFM+DTqvK3c1cAyYyNGfDaS7663hCwXi7tyDwxq6Ly+jZOklI
VyO5GLKYdCR0g+bRNq9Ft6lwn4tRdkG2bxftp+NKzoeFBj1rnYFibvK1O8LvXzSltujEAe+UxEcD
6LS92i143K5uMlakeJJ6Xou3HnrVYJAYqGIA2xn2xVoPHtgb0Lxz/kEMJmKFOW5KMakbDq5TrUVE
lJ5Wp9uj5pUHjZ48jYToJX6HpxxD//hvsKUl6H0QknhkbcUPJXn+E9wJfsFE6la0QasVpJGO6Vjv
i+hP2ba3BpYQqkEDIdqP/VsPRFeY4+7j+WeeydDsouq4EabmEMV/01fTSUABYmhbpm4K+nuyDKe9
H2FhAJeKyk+RvWVhedtSMY0OuszU+nAbx1W4YZg6wRoCRbBM6MRXz7XabaDb/FlENVVuBMeMsx6z
OQeDQhHAyJVNiAvrV8ec5mPsE6gQVzc441ATJPgUSI+vqdUHVKKxHtk8lm+oGkH3jxIYUljjBTr4
gLPws3y5HXbFPwoWGTY8gATyHko2UW4MAyv1wwc6BoEFN+BHt6VU6j/HX1WgOvo9hy3/F+kNDqjK
uVtdDm54sXFUoCoR9rcmI3NXs5bVZ7ilaK41ErvqtoVi87fh7tT+Rue5puIZwpqtB0tlsdS/m58w
UpQ9jDbyVZtasc3YIifilyt9RR2YKcmIMuxf5+EIWE0IrcVf8btSHnI0kIFHh81vT3U7hXyMXuCD
kVFn2w7a1c0Btdmz5j3Y1pt3TRn3QM7/A+XpUKspscvrZTaY0dlUlQBnXbJPfK7CxWJoBllcbyTx
DuDXPq2vzMkRnHVyFT3tMFnJqfsIV3S+g3+0nEfUKwPQjt2f77T/jCUdoK7/Z5sznQjgJqgznjep
wkCbapRooqVJWh9UEc1QAfMEHQfa5W0vjsTZCBAkcgo/mivexEoG6E7+udipaddeQc55zm9NnbHv
8KRGWpJ8TrObY5G3b5lKretertJwGn5BdxkW+pTMdo0nO5mNwAh0/0Gx9QvJHUokybMP94ir0PGW
Pr+ja8bFgLAnPPGyykUnuOjPrTOB9+o+Fmzxr7x+9djoe8GKtcw614jIG57jnUwvfybyxQ9KI60z
7u4/L4iqgFyI7sy9Sarwc6+orAJE/Ac471lVk66dir2jZcKrGHbs43QWqgju+MXIAVfb0ZPTO6U+
pYdvu+CxLa2zLrOkDuIXUQQ8hO21GzhKWQjEioosgObtgujAeGHLJts13vNLbaZDUvM4xe+ipoUu
SIPigBs4MtRWKY05MwrJoKsKfcAhk43AUifWUG/QrbCBMIIR5WNCuGwLgbizhj765vIXqsOoy4pg
0bf7orlwMOoSiQpzD19+suNgIx5355nKZeBn3/WxwMMUFzD8rSXZE/nwc3UJ3ffPg6HB1ggL6nmI
8nL8IeogdkhB5WJiec7OkQ7tYjYezgVZiMsFBbamWz89wTUK2/nneqvjQ8To1AkBxeViIjJlZqTO
t6Olc7ZcweB6j5wHWjkbnAXKl+OwCBXCxlNvDeW6jTqS+lJq2goso03tYdyxt9jJdvDWRHnc2h43
ugsRRWtalE3CbXPqqHRiq+7CED9X1+dDOlWE2frKpLDJe2BfdeD66dbbq9d1olSdPR8cL3KDHD/E
WKfpGakNjpHLrrlZDdCLImX3fk7pAV2OToMELm9bM8j7nCWKWNT6LsJ8m9B1Hw6DaXP9FLAyPXjV
yMYbiP3Q3hCbRtrwLZ+Yc10nvumFDTVmSUpz5kWzqyzA6zCZIVIF7MkQKw/KE36ZYq9VbC88WCHb
SxnYvOBnBiYHZ4NrOfw9wA1o8OB1awWrZ5FtZJeGCLNnPHCizWkqIgd3Wx+GJWi4t8woS118PaKn
c6AMOOlwIwB8mOAqAMCdEOqdxe8+VHAN5MTEy8nQn7SStpYNVpXdrRjUrqDQdpphSvAU/LdYlYxW
i4C/KY0tQBBOsrMfvPLyZkVIkpcHZAqpDjdJsjpMqp45An6ellQqzghLE7PCBoGx08lMlTeMwAk2
Q8VhMPTXAsx1RjK7beVb+sxdZ3xer/wWn15aSCYWOTjLelhaMPT3ckeON1hHcTZgLt0ndZNxwiTk
gNcarcH4inKY1tfA5v9jhe5dKbjSyYdzOF99Wv9+9xT1oJL1ZHQZndMbfntEUK7scozIexg1eqJo
LY7kLp1s6yZ2RveTfN8UowsdpcbgJpYNRR26r0ALKdeXSGiGqwzmug4EO+S6kjHATngNc1lQbqsg
j2uOedJ5Xr9kphsCKGLtLSbbFFV7BzaJf8sAO8RzdQSNnidJbFJP1GPK9Qe1QoFOrMs3iV0VK5nA
AHzc5PC3YpaIbvfUvnqjo+PMYfdnEG3xKQH+hPI0NM4D1kIh6znUO1Jv9hWMc7G45qSciQkmtooK
UFHVnuogt6O5Fj9d33fxbZnbr8pfaw6kUCpAOS71gC+jxpELVNg/bcji+TNVh9F8qI8ZpnhzYO6+
F+ciQ+Wu60jsrJsATSCcEUraM4Mxo4XrQxk3Ura/S6GeJ9jlz048uMAyOsaiAUKbeA2eY99TBuS7
9zs3LP+3owe6JnnNx0UI8W5NX3X9Y0t1NFQ7DRmB4xP9hunL1QYuAao6WckIUPF+tito01/lt79e
VrMv75icDNA4um4VPYW3UQHuMmLKyM472o2epBOAUil12CbRGmlC3WwF/uMcH6AnIaIv2QH+UaG8
khRWP+6HLeKFtFG2CTI4N+GMi2WwL3Bdw+JytHWv+FxSMq/abcOWf9E/ptGLxjT7oZDV+YtsjaD8
RxH1AYg8QMCvhrLlKWJIoGo5UxTJymBJekpxHsC9sseRFLDhQcqj9/r3D03elmcuTc/x8khviRS4
5velRvL0StL9KlT/SZeOnXt8doL6KJRnLg8lpGoXiukCjXWTHfcRI+wBhdVLpKWTPwXx/2E8o7Rr
QdyiHbYxs31vNR4DcBol45g/I4pOfxN8ci0wT+xfYb9J3+7AUpTQA6AB39UdkpvAW4YGGGzxe2QS
AG0oVpwT6pr/sK3vJZuTfCpWiN0isbfFGEJRLjbwr0f5EHNuiC72D5pMyTX/BzkUy1AVFZPkwQdW
HiNEryfp90uUcPcTUChA8NV7RCulrQJmW7D7sq3EXMp5dP2JBa1FJjc9DUuIx3zFLcH4Uqo0UZ7e
pypw8QieWkddUXpHecPBAoqgYpGSRztgRIVqHnEAGwT7tWOxh9JaOJj37nw1yy627NjiKdajhrEZ
w3Q+0iLLPZUPv3LOXBaWAbgxHALgege831kVy/RWxj70lAYaOVf5aVplu3K0PpWL5M5sxQ0QAD8M
I3zmUWMQ/Kg0EAyN9wLhACvqdzbdCF6v0GS0CizkRp1aqalHzE7iSmhankt8a/4a3Djd1qE8RVcL
rs2DOS02b50WMdhpUQ0a0H3iLUhCCN65+ciX1SoT1GVlRea+lr65IClm2xSb0r0tegrwMur6Hjv/
XB46HPrRV0aS91RAppGw3Lvw7328fplxPj6f4MoBaVlc2jP/Bd/SpbJQPIDHQS9Nburb9BY083Z0
pZby+SdSE7qUKZ8mGw/vUHyWW0/8By/g71hHOWbaldqrnRlfaVlf9qpBclYj31wQAcuNYc3tbjRY
NYd/cPf3Ff/g2fRPkOrexdbEaWDV4QMtpj3gNBj/VojVPOgeoiHxaqTQ+2SnEO0evz479Jtc9FzJ
rWZQ9d2hbGuiCmEi6ikPwZDRdl9EeY+RtXZByC1QWOQB6kBea1c+leyE67u7RP/g/VqodgIE1xOe
n3PMc8CN5bOCM+eGn2gJGzWwU+5K3FjaCUmZDkeiXmw1W4dYCNumHDrVkwoMqRU0wHgN2l2aDe1x
c6i9ZNp9mk2wiyjyxgDizAht1g+1Je5YZ991UPlXxcTsZmspsgX1T9KlkGBDkM8hAOy9Jp3Y1RLk
mh7LavRYrBOm7mSx7sFoaWgCMA/ljrwDXQUEepRRegy2YW6BxU770n4YHuq4AVDdrHQpDjZUtzeJ
yYtq5zhWsevTBF6WEoon19euM+gyNc/ZvijaSBDm1XN7Tq5G0a8K/JyJoi5Dor3q424kwVZ8lu3H
sr723lFg1H7bp2EFWstyz8i1izOP1d7jAWTs0YH+uRW0Yw/+m9LOcW2XjnXdseNqa30jp9mhLtG0
ucnpza2o0+2yHUNy6/7zKcnTgL+wfUK0Rl5KTy+J1d9wsPsIvNcvD/bLMK4as+74Pr3PHQKvfSXm
6+VljOpuIfhYCS/PEcK4uhIXTzaVU9WW1In4Ia0sRpBXJYLG1ofwvERslmkzkTgc/w9q4qLr2k6m
slxy1mLfb7KNX3yQ1hI7tNQd4PUHdELlnBcOqmxsh+vFSApbA4HRE5ohd9uK/JePyHBFff0plciL
Co7gxAAGBw0JndAr/cnNN7TPljVPW8w6FgGGcEUvYzqz3UzKFCGNC75/S4D8odAuaeNXEgtX95DN
0L2jJPJadW0L1MP4Unw2wlIshOf8LWUhj8PdAAt3gY3xBfssXDD6QJRZ8OJkbMP/b4kZZ8d8kwNt
X0Sg43dZOwpzNbDaVkL9sU8nahtleUQn+A1MiyeBdDv8MBwltSj20484Nkoh/XjEAV7IqD5PvjAw
iy0mSw7dKdsvW416DlhyN40IlVMZZMSzymqqJZ8AfjccY/p2SjIllGaelgtVjeULBF7A4KJ7GvjN
Ehvr4YihrvkIiVPgqamvVu4Rb+UbUV6B2+gv0X6T3v93ROp3K3ggTW799wGW8X7HHJyc9oGQmrBg
iUoQdE+4ITFxskOU66nMGBAOluWslUmqJULSx9jtAjlgb5JwfbAwmoO6rKdbM9bBbBHYMLkVvsXH
6mqfh+qRNwI9gNQFgEZwXkQFp0K9E414BQhBg4dILg+9cSW8HTreBU8wnifSIzJxR6FFAvWaJjTg
mgpKBRkuhZZWMa8ZMsMvVgBzMMUmIRgGBqxhdJd/miQkLmK1fjLZB0IUR/CfCEMX2HRu4YSvaEgR
vmhfilwZmqpCXym/onengp8dQ1t253/Klm5zvCBTnfbxsLZrvqxKKbRqj1ANZT13hiGbS0h0Qz9b
5PLLA0YUuhJPNm8e676PLj1YgOuzqtcVdMXloG8MtHxUoW1vG5l/2LRx0tnJoKxGhmlTZ3FSZKIq
mtwjfLEW5mAiBzkq2d5Vz9rgd5KS2QOKpXSB0MrL3qDmohfLkxSSdSzdSN4yhefYTLAkgPvjnmvn
G6i1F7q2C4sLYlYXqHym9L1XbHWeeCi7c9myiLFfcOG+1BqgOc4yO1NDNwqyWFfCYT2+gze1AApo
GCCjZZ69D9QRPb0nNd8+rpVhwzX4dFtWOngnqJyfR8lumDZCUyBsIpjsljItgQXtWFKT1A6fFO2s
/P9R1g9/eGpn56xPV8gwnrdAVfU+t6NcZw4quVOYr8TPLpSqohFqKcG0QBPS+DGJJOsQqY6jw/Ly
rc7FVtEy6gH6SUTgfz3dj3hgnm37QhyTHlLDmhYNQtEaYmEgRoVoXVgvUwi/p3KTS68bMMmDM3lT
s3Kd75Eor5d6Uicc3YjPZAqTcAIr9SL57QyXSXWQbwRbQP/Ogkzx4qu7yRfLp5gPayaF4bqivH66
lxvAdaJHfCbbYMY8SYsMKW/yozVal2Tw+3ah2bij6MZmOGmH9rS4ot4oTkFzDcpn016ZIf/O54Qx
xy2psSyMvvxwlJTw89dtUgusDd1+4b7/PieY6drkdCO47mXH3r3XVIgbgDrax23OQs6FL7+wKMw0
jr6O/XzKz8sCYxKi6f6aq3t4dYv6cJ2Ko4H7UyVELMr4N/mPMTWDZke013HCIlGmbNeqEjyXwkv3
z53rCsSVb0E2ahrUUuVDCWOvQ1nT0OMX7iQbOwEQBsxHk3nkjaTKq2UWGJuQDatuEdtNcwqwvwO6
pmW9Hz5VQmigd/y/oHVY7O7shxy/HKExN0jP/DSig8TqUvqolpPZ/a6eV5x1TZ4gO+Mw/sl0UPw8
tpVU+gW7nDZXtN/dQoymjS5pNyYIoBMQv48SlUlzxFc6YYA6fziNweE6QBb2NIIdh82pYNRlEqdY
VRwjtEILO6ZRaheeaLDztFJ0EUMPKIt7bYwRgrsVivonQwHyNVCaBpqQVnrvfdRyyxcCLElCaCXr
V5wfk0LthQG9UeHv5h4/t/bAoKqjOEdo1fqDg9LR6yBGi9Exo3aQQDOCni16EYzt54U0qqjHXjB0
fmdCJEdrbKhzAScFf3FDuYe6VTmqmYyFHX9cU8LaLUAPNaUL9TOb5u79Lu1mkj/aHFBHApVM+SO1
65R23USIxepZJOuCFOA8H/K7YjgUidyXksF3gurUCi920zI66Q2TBU8zeiFUG8GpdoAxCSCbu9Cr
0lq+k4bdrL/tVL9bmeYcav2gvs4h2PYe1AuJP8A4LcNug2z1BWK+nvfw/VNmOekNdcDe1jc2KHSM
XzW1KHeeFwe+f4NvxVqY8QHW7esSBYnCCWAi5qHQBpd+z8jCKg1FWw4zSu2RTJ6FlsN4dIxRjEf5
uqWCVqmcWzKcbM62FP9UgYCJFN9S9veUIn3mEGx2AbxjE9eeF5NZvidU3b7uRqWFKOkDxKUfmvq8
y3ddHF4FZ6qQygUn6e5iNqBv8pPbjJlsbfgKTnUyFaGYrPYp0Zeo5/K+bTkqr64bq6PbrTOOdk9D
1fq2Z74OJySKAXDsm/Q7IVsaIqLBrBpbosaAVfVXD31KWrOvYaNbFaJczB85KM1psGk0qOtPQfRf
HSwU83g4NhfZmk+jysUHLJ6H+g93cDsdSx9v68Nz5nHmEqby+8eLrKzDCj2wLCsVefM8TsXQastM
/7QUkDCKk1vc0TKau9inhVXJB1VGooRPLKO9Mw+7lYoTfSl2rXsq1E2gC6CLZKJBZ6QKAieyjPjo
f1SfPf062Ft1Zx57MQ3MVz4HgzesSfxIRWt7/Q5JSU4fUvPU1YyHEIoZ3Gy0620Du0sO4LNGgNnK
oH63F04Fsswy2s/qBINSvFPOx1ztywuN+pUVinqLejzWxl4UPwACHygMV3b+5CVxW00Q8nlsByCY
Nl6i2COXmKDS+I2MOYlfm8x8/xNFQ8SQCzHQcKOxFflazK6YoVpvbiD9UspXMiLbuXT9vwNDODLs
IJUryNN6jDTM5GbphI3HGuhR+ZiXIMkKZNZOrdkzsG+vnuGD6nl5QewlX8lsvSsFHySZnJE170P0
ZQh36Kg6L2vU7deqy6vqXpc0t3yK2BBrKOFgEiaRyBgtqyBZIzSCEEbMF6rhlJDCO2C9KuV7b0WR
OEu6gvXUQ05XAzdVGK0+hL7FBowPyuwmv4uWWCqbxv+RKijKtlowAVRtRQMbgR37tL3WigL4EQZv
VpvumM9XW1thEi8SvP4LvUPcysRdBd6JGhi8FQKGvmUlBkOnbyQ8yrPp7tgWPskg0vgtzNYSY9kL
AMS7AOev9CbpUfnk+GRx6MJauQsfm2Ap0/xG/hmoZpDCaByfZIH2mdtJY91o/1dBK5/x0llrgtRr
Cs9UDZGLM9saIWzIj5DwvjEzG76DTcBQ85oktp7ZT5FHTpCUNxTxpk8dItsvT7bcRZwFHTHDsPVY
amMzvEP8fz6qjfGlxoMdxFIvG0zMTiiRx0YOJLpb0E967Gu+VOIjdEByLWB0N+KdOe1kjUj5jxfe
lAa47MbJtAuG6LllAyOYsbdG4lJBXaVpr5XJ4jFifnLXQ0P3EdbtblbJRoGs9tzJEYe9j4kh51F4
Xs4P4A8sHz7p5s5NhWm8EQ4vjiYMatJLCKQt8m3aFCXVzQKINI6dlBha9v8BGncDugOcT4VExrTO
Bk1YgRNXHv/6iI5NjY1edCU6AHiiCELaHDw1zkbxeCF9B6VD7UahbU+2B8FbLZWN4SdGex7VSsIa
p0iCvflqhaYehOo3FQd8ew/9IR247HsJ9kgmX/dM8KAUNPqkB3RJykmV2Xu3hhvtiME3I1R6QINm
F7bzqSshEcFrctfGLisqf478Ycn+6anFurweuh71jBG2UKEhk23Sd+Y19k7CAJ3EXrBQO8fR/BA0
IOw2K2PN3equ/6oazIWD1vaAmsLHDmJViDhznyTm0KmXbHzZKPnEU4zU8LgBp/RknWifYqop9tD6
++Is34uzx38yrwqDBWYEpbTU3eq6//GVSgw2oHmDZ5/8nphP1mURIPmJKI+pbR81xGZaAbFkcxYt
lphh4E7nz48ZA+uhMJe4rxDj/lR8MQw0i2TrR819yBoAJYSHbvPSg0JGc0spfbI8YprvWQRN7zwQ
L3NVBBtjsJYjVX5ep0g8kjdx175Uq4Lj2eU8dekGP6OjjnFGeqrxrvwAJ/QmkCtCthRMYUIDfuP6
WwZzkUyOeJCvOnZIwnCvZMzUvsosrKNv99St7xap6kP54UZ9jAYfnz5FGI67HfZt+GpRFm07Zlgh
o3ea5HTLdbH8iltbf5cSotuyLFaRQTWL1Nia7ObKyCytJGcpbl0qbTC+YNJ4bsifiWPTyuVyReG5
T/kXcbNqE7H7QVzaOFXzt0HTlPvEqcDgaONOOu333RrpZ+0V/LtHqFqYMrnjHd2vN+CYoQI7E/Pu
+mOEOEPumqHrYgn1VsW4WO/ZOeDx4iQGG8YU07nbe1mRSn16YkYepiVtnc1sqXOtRBn6Wa/W703e
xkTMzmbWPvdKLIAFrI4WQVF9BiwqVl6PJdgIBnIWwoKQFsTFhtQC2ABA+fq8RT5fw3AfoUProZtW
b6KkV85PWd1X+iE/NFHkRbMmpbpapCM9crHEC5iY9pxG7xB0d2QTiBnp8XRz7VR0s99cfr0cmkbl
sY01Ruq29PSpERWicUcP9XFEa1UvO13IK6/NABSvZbWBmOsMVFHddzi2LL8RgbXlUS6vYEEXdVZm
0hsnyNDdAzFGflSwOxTxhnQ6pqOA4ArNb3wWN8WpKkzQUnTNOcq6xZu5U/B94sXV/g5fPzDCC+pU
TmfjYfvqZwdqoyVz/mv9q+ig0hEX+s1xQuuAzN6JHjB+c1GrktPo66bjQdX6yzLD3x2y8bAUomeZ
jOT6F8nF4ioB6O36wXzeNhhY6LYxhqTQmJM4Hb03VYrcFvKu5+DcYnwtV8ggVP+FmEuFfVzdhOje
fUeRLlnJ57pX8PVl2nwTdC/VG6/8TXphEEkPLV4msyxdM5+nQA0sDHBj2v5ej8rVAwRwJcOBpNzn
YFfph8v1Rm9nreZwwMx0WuQPu4rtcwfuypz/XipK4ANJNXXugOkXGm41FmjAImBNMuOlp6BAfILj
K8/9XoAzVlSZZg7sFgRDKyAFdkJ3J4IoG72SifT0rDne8TgYctaqyI+aMIWxCZuWZN/wYwzWYBSH
JUjSlDMfFxP6HhVoYaeSbAhTvWpqRDfAUUUEoQIFNxX+9ZC9zXWj3DEctvP1gz+Wh/GJpmGANERw
MqAVevIgCXUNSJuZkcuDzGYGtyxgLYsVa1E8GZkW4hE8h0CLnfD834xu0hU9rNvJxs0/uf7QYNP+
CqII1S2+u7018ycETJFLd/bCFzSDMmgBlzNg8Z++BFOkIkkmXVaozYxiv57/n5kXVgfAhACGJi1O
F6au+oL5a4L/n5OGvTWO4B/LPh9lXa+2wY65+jYrcijOOlpe5cjilyf2oQevEpk3ptRvN0wfNc1s
bEhSrRO+M63rWYTQCY3q9kGssjfyV5vhq2yMHLUwZo6mPhAVIErhTo/wDti2CVaH3ZEnNWIJlJWR
6wfJyUE9qfoIISdN0eP/H3/STQwBftXi/+msGe7wqB+VkPbRFY0S7bG2YKlmvpnH8k4BqM4usHS6
L0M/5Qb+jVl185XhInqUbew8KM+W0ZDW2CEhDn8h/3FwnJyny6LKvLjyZvoRI5cNzSRywgaORnsm
soLG+UaHmYmLH5JOAOYMofFfusR37/TACh5ds7a4WDZzq0/TO92t18m+ZELmlBJqFfJyDJF4YwRp
AtUD3K8ICNfDbeSvAGF6wSEqVUoO+qO1iN2K0MCpID3f0MWU8MMSttPeibWVj1od2o902T/ySFUt
4t3xtwqCatM+/FFF0GJjhA6qoPBmtUbSD/TJlqOI0LNn44+EOXGjAbkVi+qLZi/YjBUDkJBHkBJd
TFzG+eMC56nj8K0zgEU4iYQAAYnJZ5c8NqvBsLp7PzYYCb7W0j3c/YoFyVBAYIQIrFYKwVpC5UiL
hCz7952PxyZ+Ts/g+c+G9h1VQca7Ax78M2qa68JU5AyKpx80l0P1CLDAUvgIu7fe0V2NcZYFJocf
BiKWDZXNS+RRk2Ui7C3bpWuGgPYvJvZE53c4BC/K2ZdmWXMcx/J8vxQvcsIOJwrXL66NQdaL3m+X
BZcshPmXUQSbMyjMuNIrAB9sARqaJXkjnPGyW2uUebW7/WyB0v7bZTZlUkle0SX5O2OCcUIW6sLV
k4bsEY1Jxc1dKWgusyVSMP+eoP1CDFBamXQXXd938GednZiHNKPjsZWwciqmX69fYtVEyz10jDVw
qZLE2er5fAVP1rfoi6xrMU8i1fE4LupLXBeMI5Uxl8ALhqMpTNIPjAixYJ8ifn6f3MSqj6wpQake
LNxSyAy8Z4uVtFsO5sy/sb4eOR5E34npJ/QlBS9EsJ0mlWkpeQHpu4XuQx4q7TNibe5I700XMeYp
zkS5OT9MGiuh/PxASkMUYm57f26EUva8/Mmt4hhb0LHpvb0IFFUnEVoIu2Ln59PT3wGzmKloegMa
IDXp54/18ElHBHAv201MwhRXmY/ymcINTnZDTYFiqfvt/QKVTqXgGOk74WYpgpdKxppX/nuA/G8G
zOZqsyrKpU8S5DBoD1e5KGR8+LIJ2ePBE0MFbVKYX7dvf/zCKOrhkOF8fuAdBcSi1jpK3cwI3fTG
yMUAJmjE3pXY0VSRGfLj2s5I3AelWm3Kv/LLbYXx0YywTYTnl1q1kaEcmMhEaxnVTRyI/x+Qm6fj
R5XZ6imMOa5VbWXAlwZEbUxaDj8R23lMFgZCbY+rdhLj+ArwAWM/9+knwQyOQNcId4EKvrpz4dIY
EeepJCu7LCcNdqxHysSkmiXw8RgulvUyEM9yaHGpzx2h7/hvKmTESW6WIKdv4aL/Gtc6lK2aMtgG
dhmu/HlLvnjS7mbZu72PzAmc3tzPG0vDKGjxuAMNfq2H+Sai37/ibpZ87UTR9jYg7mSp+JdWIPQM
wawva7uMWMhqqEMRvu/stqjbtEn3vRMQVTguyK89im2lJ0uUDqTtugcph9eR0Bsair7Y3mfydRM6
qScw0NSG1wxcgfRa0stkGVUcyG0lDN1WPcqJ3ko1sW6j3pCZQW/2NTP3gHwOCJ+35PDpYHbQeNwj
64oP9Z9wNt2ibvj3Ac2Ly7jTlX7Yb3tx8MI6/WxwWlLC3T2tjLZsDFaaGJSIUDvKEs/NEMP6jLu7
utBBlMKs7l5AsIFEGSqrTly6+BlKd4aVxVme7C1ohmS59+JAGTlP1ILHaaRKANke/aOwyHQyH5wi
GUSfv6BUeFIAflzOGLoA3p/nNZiklR50G9rCox5EuJ0N5GRgn8ZuNKh5p/jhrh7rHOna65pLIrpi
FiWT/WeOw0/vhcSYhXAEB4KfOTCQoKg6T6EINGLjZtJtFnb5T+wCG6HCEzwSwCIDUdlnT6Cfdz1m
sMmyHl4aunyjzh6h0tjX3229qdopTP2DCJCjiyTpEiql+uKEACj2wDqUVkTyT/svh5g6ZIdqnBfH
G/wa53aRUKMmKvtxvbF3crdWWmWlTJrYTPnDFs7d9UU0Qo1p/Q8BQmawvWc8rbisCzi6A4Qf4nLe
/b44KCbRoVQ1zJAYd7PJSEbT8F+T48Os2lmrdxX3ZjSCmNvRgeWB17cIFimj0hkwZHAs0tzgtjrD
ss3UZkY0YYvleyAVmqk66YkrR2HIYTMNcawow2XDDNi91Qb3Q/0GdwwqjKtREJ/nLevpa4jgojgS
Nq/ZkCP/RLERO+cdLVpjmUEO0Fco9TuYTMU65v7zzST/WqO3PBt7DyrORNyBh8Mcf6F2d+mhv1yI
J4wF5VCgdmOFRilwe/dJ7tdamBhmc5Y+23Efao7PLRYu2/Tw8nsBTh41L1IoQ9DOlWfswT95oZ+j
+f2e/cxp/i8EAddBI95fy5jT6ZL69CLxus0RvpWF0jx4N9+KOhyNv0YXWkyxWR0klV+SfBaCemHI
sGKlRjLhN44yci3jUzaxi0mIVusVgUU7R4Pu7B55mBrpQ2bL/8k8Q0HBlFsIAyZjsDAXHM4oIF6j
ww18Eoa1Jh9dPuIFh13nhmQodDKr59SRPHP07c+CDPIlgJswYng8d7NynJnPMcEDWV2suVXZ6uti
QpwE3JtLKQvTiQyOElrdqtgG2l+4YaeS7bsewEEUCSXPLH6ErUhVGEUZaFr2CRGV3BWUobC4YNx4
YLLYbE6SWoBctVqsUyyC34b7FOY824+ZcS9o3DRh8Q+8LkMuQSDgs0nrBSjx8eLUOF10RLsaxCtU
5yaH4r7otQ2sLUD+dSZ56Vojzu1rtMDyqd5xq36U4FFXtITeut7UBuPOUEOCRscUZl9F9aC9NKOB
J8KW0/te1pygR6fGv41K8AAznJ9IXGu2lndQ401iO8f08N2X5dr/7SX9wgJKBb+aDK2zIy76c6Xl
1lPrrUpnhmXHIrVkKc8WzTQXOoiR/us8Dxog33clC3Eb2hk06Iy6swUJr/1RlXQXDN/YDe8tyKuX
DqDKvMPWIHQr3ib9x2f05T9SvArrXDyD+Uuo5DttWhOAXG/7eL//4nSbEHVzLVuyfYzUw+UVWpvk
3rcYO2RJw9rpc98Ft17NccC53oiwRmPDxL5Qqgp6Qa5ko0C+7zUKRpQjd30tzTi1zXlcztApQL0O
f2e8T7+wLcoiGherTIjtHDYULnYIezwQdbW65LSdp/FBlV9Y6a+fhliNMa0mgcQVrh4B8+2Sikn9
tN8lkfDZI5fCvuvbTF/DH3n2tLocWEwSNR/05Tb4MMVdYl+Cqw4KNSgVNSvCViZABx3ILS7+JSfP
PROvZ1+zBtsgdX2SkL/i6te5c3y42eNrRcXOCBGe2yQgvc7AGmmDghNzAXQFIKCXApDy1AM2m3cr
00lD0B6hYibQoUAtTIsrqNDuJR+3DP1J5vMO/Owu5m5/uI0KbJTs543FUtpsMxJ9rYLn2pvCBGKX
TN9JmeVq4lNmDpkpx1ktHQPXHvtvkZaauu9X5/l8fDjwH9yG8i2KncJLytfAG54bO6C0v/2igumO
alXVV3leQmCucr/XIJuVYr/WXSqKMg52jmw5miprWI8MJcMJo0xLmXj9HbzLemmMnbdLNU0glAvp
X8WPjOaj9JL+lhLKaDxG8nER7wTkaj1iN3y/Eze5Ec58kEZ9hL9c3XfI2BEPZVQ5UpAWlrGeguDn
SsTeHEYkSf7u1xxc1CaheEWYEF3SE+ZdDpSTIUWxc/QN5GSI0e1Q3ZLdoCm9TxiLSNtgOYKMaKNN
gZSE1CJufKdsZ10NdtKpIOwv9edmbiQBN5FPi8I3EbcirPEOBQWIL2/mQJif3JtjHYPYKSbamHLA
8ZKLJzR0M9/PcP0cH+P/3DOz+T7xbvxLh/4lM9iwOO5TMJt+tLwcUeruUm6anaQrR+nA4eFYHMeW
Z7qpQ2vwbcjjDFchno3i6csr+27XilKGJVw8zWYj8+mZ03n/wnNTP1LXMAd5s1AZsTathTEF3qP/
qTq8SVuZXuwGWkriasDYyKpYRjWrWSPn/akBVdjMe2yd9dupjZmuYiui+aoFcgz1HybxV50SDcqV
bxmQWPOiXTgkcp8TvpHAH83fJt7RYaylP/ja29RpiwDoOgvJiZxXAeNP9TQ+TZ2Kjk//ubpB/IFS
5sGC5uFtaXDrvIH4vGntY2IH3CAPkxaAjU92ELs8DRGrH9l364zQnyDF3XjNLpG6zDQO+ulnEWdJ
diSRjPrTqm/O2i5+XLcfX94e0p1nrcgueWd2JK6ppC29ijNua58Yb/hj3NBSCazlJEStm5TD4VOM
jndGksZJMnHHHtEXbWhEJ0oschJWDXwuf8w6neQ0Xq3D3Y0KSFSgQRA5/cwYgbELIKGG9IXiEx8I
4Owbq9svIF9Pi6OQ6ztlfQwhK/ESPvyPUbeTTWwwHgcqkiDiD5Ao/+14kxO5w4ma0YydSAbUAs+c
o37/YHJslQAKcXSComfdZXcKm9r8s9LTNYmfM6xGPVZM98TM6hKUugU/qzNvguhL433dUYHrd1Qa
138Pot/VaY47ADWhe9UpI8dk7LBI4SoK0SGs7uczxfxZY+pDef87NDaVFqJ5NQcAHFKVEEIQJagv
UEVYfKpVBRkPyhr1pqVFDaZXiszFs7rqKvdjvIvsLzZIDCyr85cebcgUeoDnJtDKsxoyqAX/fawh
kDkAkdEL831ARJe+Dd69Rx/TaOYQlSpm0vwYTwLRu9CGVpPw6Igqzogm89Bx2cDvDgWT2kNPXrxR
Zi8ughoGM+sdk1SHlKL4YsduC206uQdgslossxOS7PJDOrGcUZ5vFp+UHrDor4HmhMekw0ITQJ1y
1x3LBaVt2Cv0lVehPcr1U5vhXbWEd73ivmFdkEdOPVg+fZnMITpjKu7NL3VZdi/nVODb1FFTtHKm
OO2FPmlCY5wGDDgOciLFBfNSWPkP+QNf3RUVSYB3EVuxa88aKZWRiMBK1u18pzGha3AEYBZspOkp
8vslMxosVuzcmNHrQ2hfjc647rLNsOQMHzXlpwxj6diR369dkrDYHJ4w/C6S2C/p3AJte2TrDi+K
zK7MBrAXhEMa0mOI7yCodo7cJIj1+qF8wtFoeNx/Q87zvnF02MjKj7RHDJFQlrFrZE1G8/87+iwu
LBGeFG9LDpqUOclqBreGh2RO3zAxlKlLJvvUTSzVnqPe3zqk914YJM33QqVRSO7iv/MyXyAIybEE
YI2D2zT1xs0hgr/DAPxPHw7KVDZmvwtPg1JwrAE59RhsQ8iox5U3KPltDL40+hHUYC8X17n7NMqg
RRb3VAY8mVK1jbJr5tmQZJGe6Qc0Z4DwSUFI5fTWMq3+9YV2VEAXZJ1VkivfFkvaBUS+MNRyoPn+
P1dD+GhUoB/9Zz0lD9dXrEkfLi27m8d8KGjeD0tIat1nHv8gq7QySMuQZEwp/y4zi5gPlHkdAmAX
OwNKteCBdx0zqFV+ezzzRt5RcMqAUD97Ua+qkm+DEftEiQH6dM/JXb/kZaWRLfmOziSQV3YiepRc
FoY0d9B6wpEVR4umOyhHSbnd7rIWRlvyRpscYeYw+P+TC8gbvHYCyZfGYIy40vUVyQjJ1Vi8MOq/
G+PIMO+NcPgGFMG9LqNeGlK8icRMF4VIvO1GGtAI9KlkDlIioyWEwzKwlQ0cqtmsJNPDmDOzBEC+
KEox3XcPZ3IAlDOCyL28IAdDlyBrgF9mnlbD/KwXqYFziclW4I5pqtM+N52RLNTwgvNCCf8wG1XA
HCAwuvS7IWYhZgT328TjsmA+rCTNAQ0QuGVlbuQLrx22BXuPpDC7KvjMxm6rNxUjUV0P22GBGIk3
faVzmZxWQSJffFfAZko2iIpkp60LgYDPbH67NAZu3Qmos9iA6oQdPnSqvr7KkbHD/UlnNKq9ZJCh
e1TQ57atCL1ATzEv6uFuvMRKNayUUqGL3zn4TmovBVtsALnM5H2wNunN6PCCOixv+zQxG0fKxlWO
+3whQ9T7RWHraCyvzkFEMnut/tdpUNIzDj9JjfZmp006cmnWQcJ++w7HhIfHSdpS6p0naOfgOiHq
En5hwbLDebYeDJ5F4qiiGk4FpA3+i2CNILXycrnpiEiNR4NV02mqUtMOjWKGMV7mzGZBZbjH7xGA
wCjJq71hwzW2zXZcpUf+T3z3g/rH4htwZckaJz8zXlp7zkZa7XldquQAJ+7e+TElNLN4+Wwz36GG
NOXdS/pF3y1TGJ2idEOLYZOY0KCQMNcDHOKnLmsdL3vJrxjQACZJZMzCWWAisU/qcWfwB28bFRDP
6k1FgubHvEDSU5wNw+kpago/f8UphwFZSvPMsiM7o0ZdOKfULPOlJTiDV3UxuZIoTzXS8RHd44lv
VV2CXQ/cytPIYG2X1vqjvBnmBY0dpTXL5SCFpVnejQwb2kVWHbcGT5azRFdETPE0mj6myvU3urjy
+6W+Xjc5ymhXFJSQTmFKCPz0lhgv3NocwTuX19pmF/WAkLd/CAGWjKTq8uwEcULq6klAoa0ffUxf
SdUy3PSg+87s0fNQbqu/cwgsUZz2d6LXgoqbQFRwwCjPlJtvtzn32hmBr5awiwQQvx6oaA8b8iAx
5uXwO4lMDLVGU/Ti/5PcV7TzAgJmEUaj7VYoWwew/zVpJfpBehsEUhePa45AXPPrvV5wENMGkW27
k0Yk7V2ZxVzvLuwgkQcc/MLvA6gBJrvjAjVJzC9qAvpO/iaG+aS7WLQ0RmTCJg8GuYBYTztBtQUw
+kDitX4DFB8W9m4iU9W2vb+0qLftJDHKG8/i9hGg76usFqnGktPHIHPBZWKdz0/YWCN1XNLw3CGD
xSULjU4ScR325NGsF1rOf+PVvIBdyD7vp1aBdf8NiQ/2G0/zKwx4BbZltvpBM2+bFeQTxiUvWSGg
ELIfKzKD6xGo+ziaJRbHAwicDj5abfwqMXavz9TMRY1caqEx5fOVaMduCXfWJ+MvnXu+GEOPlM55
0eK9/5jGXBmYnDOcYG5Z1qGFhJQYLATE+euNKCTL/ILKaL2pfRab6gVe2QuGa82QZU8lcRzxb63Y
vR0ZoCqw4jM4wTGTk43uGcqdtMmss36l1QYtmyaB4E1ruYEGOESGQ8x/xMdjBcckHljaKDoRPgd0
4jankwwMeEmN9l6jT/1mb01cyAq26AwDd1DEqZ3Ng6SWXARq/MgOk1kd+dWJwbnFKDYK/BiFbuUF
2aKIzt9AO0TRXKBn8HwcE6WzbDP/D1iQ75MnP7JwZVXoS1/7T87RiKeuvLd4PjXXGR9SnMeOh0Fm
Y7FW/0cbrcKuTFwDuEnaVNOFuiMphIGa5ltkkGQMdVabDZ4ExNNKLHf1zuJkXL0HrxPVbngMbKVI
UiiSdEhuvgVcmMya1fPvQ0OuqGZi6wcmPJeo7iH7X8Ilu366R/onrZH6qn9IxTZxM8tF9ZwOf3P+
CnY0ln2d1RbSy1EHX0+0V9ETpacU4A/ar4zD3ubKEt33kQgox0uTpZoMbksxKUP3l9aV73ZcSl3t
4y329WOVMh8Nq7ANQrDXAKB+eeSb7rtrN4TiiIOrboPHzaUeVi4vJ4qxkS1+4d4NSLn2AV3l6b/F
ecS2inIhfOFaNOr4ioUCzDcQ0PvBTfK+IGxA4A+9GI3OIbekEmIUO1YpmqpZmdJwlDdif854KGmI
oQwp+Yr7LuAdCzZfPxeXjkM2qKDV8hVPYG+VaWOz9MUoQV2Nun4pEwieXDnRG7sOtmS8f7S9flqx
N5h0ZKaCpsSKS6z5DIcUcD/MgHjf2GpygdCApeTVhq9WGm+ZpUe8AAL5bmUI2SW26W9nJ87WZ/rA
u9OzUMoq4Nzkulhf1u3AYtwgwfiNe3taYZr4umPCDmn+FWu/z7k+RhnzdyJBnHzqgyo3I8lMfXxJ
VzXMpWV/bSkOndKIOrVkN+Ib8XeEBOlB2adIUcrxBPWnmPomUBdqc1P8nNbIr2N7FbhQG9BRnVWR
8O79as+hoUoHUmYIstwZJ4uoUCtITyxrdIJi2tKVvBE0zjygYut9r1N+zjcLRt2ZkKJYv9gwbtwg
Hc5mswCA+rnh/W47mJCNZDPpjJN+f3/qPsqwbVyaJyfqIGb69yKTj7jJ9J5h0ja9rKYOG8ggu+ZU
Hp+DvjDCnRu958GtmKSsncJ/FF2vkapzHjdhC6Te9/cTxrk+uNXAfK9wHiynUxq3nffOeiN+U7AI
W6EE1p8zCchpLMvUq7C6Atu2VMuRgTZP7Fhd8/51cxbqgDwZul3uR9BgGh33raaUolbySObo6uzn
/3DPVBqfXeATczROxOfMRs4Xmx+hK3c1qH5QNKXFsKRsdeNgzcPNaLLxL5j4WemwUg1QIbTxg2pU
WGc/DrvosY34EFZWmJhqDyRgKetB0oq/FVXZQCCcJmvRA5X7Nq6hs0jdhwq8B/LuyM/XLNfn8rib
ZQd1m2XRxDisnPHY+pXqOqkPb7F4y6UvnjRJJ0bvGGuP1D0HU4qntDOjsGbbd+Yy+7UKfsN4KBKs
JxjXnS/5CeY/XOXXIdvPRXBhXHGg3tpuiZXpxn9a1jx5SkFz7maD1xxbhhyR+LjE5uYCM1qsJ32j
DaDGuw3zJwu8YHrlELFsBEELHn7g7bOg17I9su4e6ORSglObUxM6SPRSfBdeoMfebes26fVjkLz4
Oz9nlcUS7szesESjsHBT3fj+G/2pidZA4eytIz2nvF8bSLzpomKOMiI2NIH3FYXZRgaNrdP6AhNe
wFz+gSvdvwHJP1EPFb3FFf3bPWFSkx77n4OyuFaqYRt7dVRcmViJx/wSleC7ci604WYgU8CGtF9U
agZ6gHqYptSYQmwgjjfcZIAxyKGhpAEgCbCkzQN3E/NRRY7Z0kdCWhgLHuaFo7ByoAItAqDt/teM
jTmd+BOfYpjVvXrLWPoc4UIdehsEyASMEGj6WQunBG+JNjrVdF36UF1v8gEI3Treb/PpDCmpdpZz
MgSOQH1zNjeBwEHQhnc86Lix0SckMvr5sPxdVpGBmAJiwC1pTmUFbfjGdDwVKliRbiNXYireqOas
za5+di6mk1zkM0l4eX8PYcyrclqW85KoMQiAKc2Lw4v2dhE8yQMjWK051GYk5ad4o7eFjDvvS1OM
aW/uky1q/lzHligMCKEYXCBUndMsgKhtom20/Q9fwRqmfeeZUO0zzay92fHykUSpPc8EFmO7z7O5
hP5DCdHjeycbhYfhCnPHeH1/tU/zPIqlEj2kQG/PrdLsrj1B8tfoUVejYCIcl9MMC4k+xpmCo/BD
kWO/CxjUcfY8InPJUdQGJdB4aAfKhL2lC9kRK9cIVVPXbhlnEmZ0FIOlHbZ3yqnh9qu4QVl/PcN6
rVZJRgQjF/t+kaaKiwkrtQDD1U4qASEiJQFoHzOHexRCw6E8y7kWqy0KQ18CR0GeGtf+OtQS5QhI
4AIvUlAHp6sUp/229JTSPskiwSk1sQqVSjLFcfr/U8dgAHBvQiNOpLWJiCTS6/b9Lh4khIyoJQKL
qJFz6N6DF0Z2ELx/1Z9Jyov2oqV9F1d4UgHHVbfE+YtvUK0nZ+NN0HtWY/YYHQtKSN3BnybTIk9A
DKhzdnCxnw8L1gakZX9EMkD++rYRE6EJrGrdJfzAGOnCzNt2Z5HY5SiGCVdTwj1jprS+2qT+4V3Y
ttDTjoumtydowvpcCOQkWnBMxYlMxsU+kim7oMqOdh+BaVrwXDkyMqtysrDnwqSiAAfE/FdaswoI
wmtgY0UFt0LMidVTcSb5k8QrjkTyknqvNOaSRv27u+NPGiKpZjmwBg+ZsruFHKJ9ZsqF20UoMQVW
Z2n3hH4Y51lTH0H8zlPAMmw/ZSo7bVE+rcV/QySFJ70P08z6KtZioqC2DoL6OkN6AYP7geBu25e3
qw8imuMveY1+BuUo/aWxwHzM7GeZCaKa8qN1mwXxtIvKSJHUN3ElhHdC6ALtbsT89slFEF8QYuOg
qF95rkyYtcuMgMcB5ffcMXFTtoav4tXbpBPo6zrjXClH2L6a8Cyg0fP9fTucCKded+B+uwW5tQnr
7oM6E9hMzdB0TDjVwR4IS7xPHNSWm6tewcYrZWCX90t8Uaf3dR5I/+PVu3EoYpRI4WDPaTPx4Qx+
RfCKMJ+BFc0boOpesO5/KW9Nf+htdyusBpE+iPy13nFP3kAObyDKsn6CJ9PVdUtrlxn5d8qh4leW
IrNgbuzJG9ucPgspZjb15VeN6uM2DYijJPyEVFtdEEbVH07Ct7FuPT12DU/qIcW73mPxy6bNyOwz
gJJErNE5xf+Po8L3PKLbXR+MqLWLVUwgYohzb4PoRqaFLnscuMUTAnTTxE5zpCbtuslFc29+4DGO
b9FO8wsMXDHK4y3sDf+O+0e3LdP0SJxsRF9nwNDLazsSZJtGsySUKaFOstLCD0cYa9+x40NT+b04
Uj7tdIIEpeJOpaRDMa87oaFdkJPiPXQGiDEWhdIrvVRYwa/sS1FWQ2V15yuVX2EgP/GzNNxW0ER5
lnzQk/lldcKeMA2qcYArDF87OYS5iPK+JdLV/cuyyuJ6SJSqP556BRQUMWD5gnTItdeF2AuJF/PS
WFMa/LBmKOMauRBBmKhNZKNrqJ2ma5wfzUlWwi47Cxs/vbt/snpwGoxtnu+gq8Qvn3T5KNwVNcCL
CHF8SQWdSZ4aenAv+xnfO8IL6/UCy18/5ipl558MIe6hP1YdFhonVtQU8YodsMmkd63u+ccXyvoE
QVXBPn9LBpmKYi/OKyGHBRz1Na0mpT2yvE6BTujCsMw1QNmreaXvSOkueIoBIXqMtNh3aKFgRXM3
SGYeFgAIzGXRumEDIbIMKP60BsUX7wYd/+Kack685wNxQf67EdgyaZO+fraDgZnEKEDDK0nc1K1c
0Qvf5S8Ax3t4FEw0Kypn+1/CtuwiOpTBMX4DBlCbEZw9N4nMaeq3LQZYYpl743x878hP36kV+HKm
07pKeEzI200ovn3NwBxgMJemSgRbjlyzW8XLK/gjWlr6AIptTdrD4juqQnbh3Gfeh36AWf1dUA+r
dFW4WJujFde6VqK06njDlcSkWMMGNXslaV+QbWK/epAXAnzzwE1YA18TPcvi5RhAHFZifAx11/jp
tin2Q1GvACp7PZvc8CDad0GmD7l4FEIqWJNqpPSm65ArFX8PEq+uSlYRRDWFwJQfBwnN0SKgE6LV
GSD8cKhi6MKnxNhfOVj8zYcANaaKyhJvzcGQKySbpKD6XR/Q8vfFqMw+4isqwOSsKQhs0GCRiJJg
/ggdgQqad8RZ+vAgO5L/FS3gvaZnKaw8k/rVZLWmIot/mhaSxVpLM9E4Wtuo8VAhKYSFx4FLnewj
oLAz+EMYIhjrY4NLjnnbnOzVHGmj6BFXDTr0noup2f1mzvAH4ocMCcp1917d58xKHQGS37s95jzt
zEcp4IAmUkPVw40Oks2G8Pl8rr9gLGczUE22mZSu8jLbFuBeDE9CM9CRhlC/vXWULCNP9RR7O2cH
g/12GOjTywA0RJeZGrNvjRFfsv5PDmYL8s4IaQrktQ3sEkBGfxFKxjl6v6MHQ3OCK5Vp6pNHLlP+
HYyqZQbi+wYGVfxiXKHntykG3cTk2eWdqBR0eY1I7FKxt2MGtX61xhFlH+Gk8ZX+HwD8jSyXlMXo
20BGK3EWbvA2ZI83R9kvrA9acS1ILG5kV1mqsuDAjesSB6bXxwzA/JTaE54HSvXrTeh9u4X4c4FT
OqvNJeXeIPfwvyt+93nalcudqzkrKHScLJuyezbZM0yogFlUPkR4yypJMZWiAEgqIsnG7nA0Z9vO
5DMQUHs9Zmap57s+gcKP2iD3wEP+xx0zabPDxfb7wHRMRWyloMbTb/njl9odawkGxrPorTFjPRVs
qgYwN1dPvxGK/myvtPbOiTHRpo03qlMYFkn9PPtjN5FX7mbWIQuuICwh+9bgA0HmLqekp0/F57gv
cnEImxY1FhBlWyt5RtZVrXcZl56dWU2WlFPvPNwXovkR7rchtrOvh+TgYYHcss+1Prdr0g9rDClg
a0ayX3PClrGwmss+8wXSJE781i+jVlNJAVoPzqkuUPpLQkgEB/5TAuOo6qK6c9XON8IhzupDf3Kc
Mz8cQjEEYlfg65hRuSdq/iEdj66gNH62/qrEu6YF74TMlWhjTvepiJrOIAVvbDkMJE48fTwENeAz
tLOZhZOx53n8qJFyxGmjfznhc7Y7SbYbhL4yrcdhhUxttVHcSZHYJ9s27O+Tht99mF8QMB1w61LS
3rU1Oj0tyFS8NnFS2V4W2c+djZhkhdntl91CkZh1TtxW6KW0YxBlm4/vqJ2pO7Md5qSeqkiSeHiz
BoRQ5gkQRixQiI0byH5M0Y0lNeM1kdYlAXBc829/lfwX7Dk9k3CY0pHBjjrfsIvmS5AjxvZ/OGYC
ZEeFUhQBq1Bg3CmR6uL3AJ2xGYUKtdzCzZKUP2LlAhYuvhYTBlDDPYw+OtQSAB7U8j9EA43vj5ww
CBhqEfzJiEVc21n6Kmg+6W3sFhJlQBeTxLHGfHBd/WVeUUYI3DLE8pZ3zHx2PX10ahlXysqn5xbX
5WqWlfFDvrINiCvxGV0L8JBBlovOpS8q+O2uy3iq9JbOVT/oOjWSzzeAziZQwnqm43sFtorDEvX/
WnDe4Kb4UOMceG/yp7LnnqTfIhU6YVeuU8YUgKQtSlSag7TSf44mkGL9bVPVcpKiqqZXeSUuS2gF
ez35DU4Qy1r5us8DBF1C9AqsX2NFEFAkhwTwmUHtJzwCY6KfgwmEpbdZZGPq0m2qz9aK1b2GDnv0
0Wn7Qpqn5rimn/zx+yLSsX8+D7fK0lSgReA0FWdn+6Zn/2ENRUnk9vs9DqZDk1Z59gbbXrqZm2+n
SHO+1EkqLHZUYuIEYIJD+3xnBJwXf7RAWnGEB6+oNf13Mf3UoKgy7Be25Oe6IgUJPeDZPaPiFKKN
Put2iVjRXKFYuEGKT6fK3Ni0i+pnM5JSwgTb53/P+D82ZT87iV9IqeXhuMLOlkMwY+9b4l44UwJp
QnVPztbwBOgdAQx9HO9XlfB94HZaqxxK0lUC28ol4rlWjVF8cVjJh3Vf8nbX8cVqKHkUXd29I5eO
3oZKiBY+o3LxO2+k/rZNX14Xrf2W00HNzcNpA2MwWkt+DZOV6cs0tbxxpSX2yuLEJiaVs78u5OVD
FjQ5Ew5fxSr1Wq8wO1RdS2lMv8ObW3I24xsdDvIbu+wm93wFOjSmzSTZm8d/xSGl7KYQ+BctE31R
/oAgwve41nHbj4Yn2fTMY9dCnS2MdCMfA9l2VM5qNgm150mMSoWIHnuVz4OQF501da2dct/UkPyH
+QiUhzlvb/3xDwtSgF5uLGi22We0oUWkAVAVLL0jtPL0GnnrN7N6+z8iHsJZwUt0MHOuToInDW7E
mpeSy5iZYBkijP9K+aQC63n2pKpKhCsPpFpVGBIOYM6Swmr9/ZvlkUjhK6lGkhSnV5tV1vuUWgnd
WsTEgMjidP6XOB2u/GHVRRsGxN8yjQbdP1x08E+pKl0FSbaZH4Xbhv1a2G5YBnQG1fEA6VW6Ok1B
81nWtI/a+tOLz6dCCKbfSYj2S1ERplTaOTdBpNYtyMAvfw4F3TWSHb/Ss2nvM6iWnTkooYsD7HnR
zm8rVNkM+3Q+sZf2PJsr9IIjbZfFq93GRlK5sJSL3AzoHhiSSGOHEH8qQozZ4UuT2LNCaV0OxVQe
zUxkKfRgjU/UcOFkhqAqhw4zgfpO84ahKjKL5eh2b3Yjqf1QuWPK9VNysCviYvFRMLn/j4EA4Xj8
b48WMPh9nJmaeoxH74vu6dowsDBVuoFAM9vDqxcMQ9wEQrg25oLzU2/MX5gqbUmliRoVMK8GSrF8
hj/DHc3nbsK54z8yhKkwca4rzzF/CP7Hdqe32fjer9rDOMHt2QV7+mAJ9eU2wX3fwbz6hPgMkSn/
+vtEy4vI/UT2hDOuRXTqTh3bYfPk19IScVsYm2ySRmjHOcqEi0wYMGFlry9Kxxg+0QyaNTO+GbD3
Wo6xIc87DmlKQxfTWru5rGfohWI4HwRDGoCFS+oUnTsNHNPcEBTdHFnPY0Kyb1eyS1rFlFYZoBpD
mzkRaTPbn5MYG0JOu0HIWRstGkrir4MDmlmeFsIhgFkB0kMS5UVd2yDfX4S7SaKdQeoyWfGP3Zss
M9z0QqFRs702flPVaLI7e08fDKzNSCp+ni/IiQYPXCWbxxwsmnin9xRqqR8KseMwxvlOR9jV2EmC
dTA7T5NFh2UdajCT4xl6b1Yete8/xDSRL7O7sAudHzOkKaIDloEhXYA7kvRNE5tyvQ6hcXNK96RE
GapcFeuteMoQ8FAW30md6ot9jB7Yvisf8y7ukqivBc9Z0ZqCu/QTm8p9kPy4j3KCccONc/S6RQoh
sADdg+9p2mvGEufJ+mAtmIfsNM//q/t77ARxCJHunssKT/vm2HKcQ5MSSDurZ2yHtCM+AqXYiBpv
wnvSOSqQuwKo8VPgXKd9CxzN975nndwB2mYCSPtvtanzxbFEl4gcinClMclM3Ct47ZzkP8gcem+K
okpXNoQREByO9PsxkDXOPZWpMeM58IeOKaB3c14un+mWd3uYHWKV2Ucy3saanmIcjjwlvbYboL8V
D1Pd/wc1265/Y2ET/KtWSRGfr9iaJ0/rPp3Z6Fvua5XboC/5DskMxGnwvOLkTCaL+2aR5gapFSFl
T3g8d1gIja6mnFhme3Xhw4cQ8UcgaOznzUG4fppr42o9IdWtnmdIp7XmcNBKi4cTe1j6jn2szVdl
vMKl4AT/Mt4EXWAYuIxt7vKSviJ6VcoMjtsUZKefz8H/jVNdQ5DFjwBNQTHhna2ykkCBFC1EvyY2
lsd7lgNn8MfUjiX2KPhluDeVa7SsdXmUwzZCMZazg9J18u4vvfM1KmueP8UzzeHs93SPrXfTuwT7
IR6lBMDlcszETXkbOzF+8iaJuQs6ke/aEXXyKyb382l9KW69cQD2gxhB65zmZUsVv4EZ2UnjGXvY
OMmDXI1SkvwpcHTFoXVom6FWS3HkJQ9by5gkxtrLYrYHH9GfnMW0SGtu4TPuHIuk1PLefdf5P/1T
xHGq2bBi4ibCSbYw7rTSWwwPR+CUDEI56E0ZihQUtLzxNv4t5aijUiUqg2I49SLodJfksoJbddX1
3zpNHJfBX73+7ppKy8OIArtIw6hctQxDIU48tTI62zNAgpR47isiQslkaP5Z5cubZNgFtVNqXOY8
hcH1LPHFHsEEeQnm5n6exCP1eXFwQ67uV/9hMY/ae/LENF8K9nHP8PrwAyod6hDEf2BpQmt5GWLM
YCs0jCB3GA12A44UG1LbeRH75AnUOP8W8KWFin19lEifMo11B0bT3/sfDN0DbgCHER8diyzNZqLO
BUVeonOdL2fE8zwr9TdRIvLs72eSSSkqWhq1osOrrNQeXZC4UFs2tLH8t/ruNlIywPqZ5i5Jd+Ez
RDMas7XXvrb/TQtQdu2EP3HfE+ZKvYNzARxshlhQiIvLsesl1Nk7m+S6kbRmz3w+rwGUfYuGyibE
qM+3m6/S4qLZPPu+JTx/kcir6S2gCgQrkbE0QKrknUO/+o1HWjgtG92xZ8F5w/Sis2ak44hSUJRA
Nmb2nTJ7CuXkdlafQfnsu+duC9TwJCxdweyW01nb4fSelo60S9b7VVMkA/4oY+8BYSwhd+efCJwW
Zwl5d/B/7rGDHSMqdVrVfjwjAozrDqbqlalIrNKhNRpnbbF6mPfwYlIAxGOG2FIj/urOMfkzpE8V
qGaAUt81Jj476tfqVj50HeIMIpZiCgYyVV4+vYT5B4qvNrasHhhPRNpQmfOmw3pHlQY1mzGb1FER
Ia1aSyffxGfuwna/M5iM3EuwrCZBviE/fBSoRqTtBv+z+8aW7dq0n5mrMqrWHMhLb+8wLZFRAtsp
QGQlzIXvDiY8Tg9pNm9jMvwPi8VoU+tz8qV7OrJJHQCTqmAxEUufbvMpcwgFweBuvUxKvQ9VLTQl
Nt5QSBrD66I9P41vwpeBxMxUESF9m6N0nZxhJXK3XJjukmpQRmVRXSQkTIJe0gT8G0s3CoiRBzGp
YWgBdrEnHISMZsSKiqgWzY46lo3tD6XYjuwdUGw8ni17513szleoF6O2JarWWXMYNbQnGg6nr3A5
8ESXYt4ONQdKf0Jf+vNQMPpmeEAFy8UMf2652YoDIOBhceNK4JOszb4v4ByqbnmZiBGRd2/p+hWl
ezBe1W3cTITS59rvaou2TW0N8EHf1uXtmle2lvk/Kcd0bME4SvEgzXRZZ6RTGJptmUcKDNx4bptN
WwE1a2bhvUVTEQW5nmnqq97uHH6RavFL4JQp1N7mvQvVXVRsbaIkMZecrKw25GzO/OskeJB4BDR+
FjpfJTC8mIL5Q8TjNkq5yYsNIDok1g1mbE82C09vOoUO1pHGuMqxnBFTHxhqHjhZUPcmu5vH/bJD
0SVE8KSg6T5WRfJCHYllYLs5x78MIe+QJCqTZTDzKzeOWYTF+CP3eqgKxWHibkqMHV9sLDLT/F3z
yzmp2/1CBKtgORVtocNoKfxQK+bNQaOQSkSEbP9bNS4LRbRT59j6xLP2HfkeE8WaU5HvDvEG3tce
90Jsg4hBSvk+8/XCd3jXIBGXlqMA4XSHMpIWcE+4hsHrniCmpbRhBIFWO9Q1YXunNeRZgo5peOuL
OqbLtg+P4XXbMCk7CBNBvZF0SFXaCMVNrc8o2c+lj3tUff0110yLzQngL7A2Ljt1N5RYvw4IJ0ab
92ukihZM6R9EHFZSpymOoVDPKT+g4s/7Jow+PJyUMilyg/I3Tup03weqqK3yLNsp1v1kqM6TadpG
3Okt5qwtcKfSnL+SmJiVAvOZEYrW74rwCV6hoOX3cYw5Ko7M8Fc/JiUiE1AsL3PWf1k94qiwO+Qj
Ucz99NyI41TxIDSJ4hBruVEsLF73PNDZ/uM3Pq1VubX5eoR6W12MoZa/3jgMpG+I3N0GFBk1dISF
en4CPu0UMIWSzPYly89IhrqCrqMEN2FBT9lXkfMVo5uyas1c0hjqwThZnvo8RkvhO0mDBQ/bfjNv
nwjKPPTygbIrHplYujVSOWqR1xVYvAWWaHAUflsdc8KSlTiIqxP7w5rdygEzawYael61prsCr545
ZNXwRNcSAOzIgAmcJnz92XxslZ3kg7xNkXicEtAtWavb/o1iE7/b2cMaF1VmIz3mBTatwQ9bu2e5
myiYCQjrWTjTGnMDb3Q52lLwqSYmJAsrWuB/Sdw24g2W1uoTt0XyS/8KUQSikuCyFBHW0P/RwOnr
UIO/JLt5kOHX0smiWpeUEz4iziDCQPLIU+zbynDpcVt61U3CBZbT6wr/geTvGFf2GTDMPwuibxqs
YelcxRJKa1FtqpxbOanDIvaBRT2ZeRmcA3oss2RRJfQrXHc9zAMdi1gPRE6SCVkSBZhIOKEQTnJv
fkIZkENvHLOn3a1R18vhSmekQ+iEx25tepWcsPKUiv4y5ct+kogYiiDxBqfBiA6mkw3HO3tYf5fZ
QgC6qL+IWYLVfVgjbUaw3n7q5ZVkU3qg0NV/4Vr2aexR27dyijH07AzLhXQ6QISH70KgZNW82dEV
2jpe1wlVpRLcoOkuC/wOD73zYirkoCtUb1bLU9imqC9/dwwpAvwf5+feZ1PEavP8DcC8HKFAtEAL
QPm4L3ScgNcHOnhjozyMZswQpJuV+y8GyfSp+7z7tC7jDhxUZg69oNxShVZRlRPjo3VHjE0JROVs
7We+PkbmJP0n7MWoqciGA3TmPS768kshjku6FhbF9Ln60/A8oJHWAYjfSfjGQMSLTF0HQwrymrV+
SPXsMw2FIylDuWfEJxUxDO/Hx07+IJgDRPaJrRnHPfpWNdv8TcnD3313T8aT7+3RksKej5sIy5oP
yB9LE5md+cCvKoODx1BR09VPncpPtAcyISgy3Es8nmKF5zxwPeLxTUaJcPopTIWgvR1iWG8vDbvF
FNC2nWK2u7496Dq15KIoulD6KaiVD53NzE1Rt8TxDF84a1C4YhaKxzaHjGkKFnb12T0QJyhCJeq7
vtgDNrmrO95cOrPrtkPpGD+44H6UCP3oCOclsYC0PcwD7Ixi+cMpoSYS+WwKpSjai+GE2TsiKE1X
s2bYH4gb6y0SU5Y3V7vKuiyaaQrFzEtffcOFeQHTtg8NW9DBvFwrDkFn9KA6ayg6yLazDvB35zxQ
vR4wcs+/NHLx23CJEI07dHKao6+bT7Tvncci665lFym93g8726qMGrGRE5a8iVTvX1WXw3V/WHFj
R2IPOi7j+OKjdWVycfwXLinPe3yATfLZ1NixFXsow/Mfzg/eAEmy5oLLD4UVwCVTRmufr5JWUq9n
MdFpYIF06NWwtmCf2LGvnRHyyviIpK0u11MyAGrXK2f8Jv78RuMsjqbNFHJoD1ZJDjIoV1pL/9gU
U7VmnoJ/p+OWIvt1NcO2id+nPV/tEHgTdyn2CkUWKfGvDC3xyqsrKy39Iq5pl7ZFOi5Mlt7yYbtp
TgbVfxqzL8QeFOVxSDGgnSGHFUyCkClRr+tmH6CqVY0XMWrq74RtfDsY+zD/Y9qCyuusk9lKLOGr
h2JvpFEePO3shIUVWrSU/h/y6z9vkZx31VT00+PGZCrvFFhjBiwR2BfO/4n8vMXuOBX+1giACANs
8wjn7MZmaTGZX62tKavsNnWv+rnGeJ30pLH0M5PXxoj3RW/YCgTYWJHuFo4RYXqoN29qzUiCdfTg
mcGJifA6IG22pBERFFi0JxqAWwbbZp+/9ROUF7LvA7Rf7AIQ3c9oWdqWGmvllep0yHufwpsSJVEg
CGeLDPsfcFNmaZFqwu4kEbgfww+puytEOAV8eylPvEzOgBANS33G5FgZNuHzsC5g+oiIyzjUz8cs
u/zOSAcVOArvZk1w/+lyhp76QRSDjS9WKkkG2cUCjxwjMnmwv/b8cqIqtHWWRiss+wdDPbGMLwGP
Y5f/8Gv+TCQ8HqCGuJUTAf0e2ogNlYvlXUbubZVE2RHvgz9k7TU1ANcgYskXpoCEEZTXjJqH0ENn
VJuMr3+29qQSt2qtrMtFZDqiZpRejHHb9a6pDESAQI4tyO/DERusKXZdW/9qIHVNVquEkaIizfM5
iPY5z73z0lSO/H2uCRN1Yy5bJ0i5zVzJh65HvMoteoWpesfQYn3a3NTrWyM+gThvxi1vvC+pOByr
LvYOhYSOXJtfrRwuOc6BKR/O9dwZ+ONSjTc4wyZHATDXtLjYPz2mU8uJhDGfkpxAW6g6verv0U81
6TAUuSmBkQIrxO3NC48iJLaDpteWRrSCP8l8JH5a7w+jRfwu5HEY4yhRK6PUAXpgp2sOXYXhNU/N
HwR1fKVYHh5znmz/g1oI0E8uIgpMU53PRXyjmKcc1MySuDbqugR09pte8/KZTNzgWsuwLGLUVChA
biuc7XSOgYIvJut1pL7bU3bTFvPio2e1yv0w+jAsFy444nuWuv7Ux1yKYF4azBhz1N2hi1J2QeEv
Zkts7lW9ibN5LbAjaFl9pcwAJkxKJj3g0x87Dad4TC+SN2x4JT/QEPsKMyiQzJuNkEvnjfbdUtti
x8B7MrosnbOu/Vyngp/8B2AT77QhSOh+vQ42xl6QpyuGOrJY2Mg2Lycfkzpxpgb328Pm6FMqUAn5
kcnEeUetsMOJp66i6zlNc20lNiw/hkKtYxzIEOxEZ6mT4MmPGfgXOUqihNrQpy1UIgHGCJmY/2nc
2rRVFnuU/tH8KzTQ5MQb3BzlLb0Cr304EDmWhWaw5+vp0Bn0KolYtuPB0o69anHu8PbU8H3Mt4ry
bqD5AQqKCOQrFI9siCPvC4Ti9JcJEp5BfLB0NLGYXMI1/Dwxc+PDrOA/z/Q64InQhChU/k6rRUuN
ZLsaJvYJYAB1CkPc9kT1PU+lhK+0MJSEMCXM/gKRfq+8CPsq/pjW6VsFDl8LXgOTLTwi74wrPv7B
FXhbYWf1Y9SvdpjJy1PKcr4rydB8P8zDqTK1+ok0vkUapUN1oZBeuYCGFXnAAECARIEm8MZm5X+u
0N7DyMxGCIoWERmN43AXYMcxeZd6VhOQvyOjVE1sOtSlkUr2fkXZeaib843OoKK7cOc1gH+z+XoY
VcbsmBOE0Zy/yZyjbDGFkej6wq2EYT6AsQ8jyYPcuIwiZbMf0QmU+kq50ErbJ/5NKhehnapcC++Y
l33QwifkQHVE9A51WYJza5842U1iq2Z9HnP3H4gCSifXaN4Nv9PrbsyEnsHeIgV7FqK5knSBv3Y+
iXb5Yp0A8bPBeTKWcizcSO6P3AzmG6CWwEiBtmmEICm0cpotqwyuyHKoJWafLhWd2pwjXLqBDxZt
yseTaTonHBZppvWOVeSNjtgJKfpD6/Jmt9oXgL1wk477WkYi/8h1heAughVsqPDGId3eXkm/vMAz
tLjA6DiTIkPlrePAKl5LGHcOaZ212NFIbd1wkizOXpBj+bbhN8RsBcPi79F9Wo6z2i/RPp1qA2tf
6kjkfbanvLKAgQXczXt/iYfIt1d3Jj5PzILzWmSoJq1uV+OyDZNdM0O3rjHoVFKORS54i6DySw7P
JFyPyJe7V5Y3XwOC7LWRsm8FSjQpNZ93+9jR87149Pp2KJgGLRy+N6w7yu1QQxymb+lGf/MToAUR
YY8ixliSrZ828IFIU+ajztiNT/6UVn4xK81z2pMtBnKkI03aK7i+NrlIMMR6Dqq7y4PjbiD1QoX1
rT0hEU3Lr0TjimTF68sEpcLFM/1fYVS5rmF/geUcXnDCjNZMH6/j5TQZIplLEcfi42Gkx6updWYE
G4mxx2hSIU34RH08VV0orSpR5Qj/A/oF/xuhHrGgu3T1MA48a5hhmAOov6Qbg7sU/WWH8etUou7p
oq7IuCJY5xarYIF3U0CQcuFl5pPgwXDUFJt/VqJeatmHAlf7hUriM6ShCar5jqarorS4SGWKeTOy
dXjXV168CV0jcRLEcr/l5JbNelqtR2dRncF9Hz+hdbAyWXQg2+VJpKSggUSTE45LpM8BhWv1EDEQ
jNFsVi/JXKYeS6a09v7HbnehgA9i+lC7APmh35pH9rv5eQOJGKKJ6m9t+jzutSc8s4QIDz7kaQFS
5GvXknihgBNwuwnHGCUFFHffaesyDT6EmpM8bfQb7CULjqtSdqOO7qjSjLYXgs3DIT1xgqHODVZA
C9/w3db+5BJ3Q9x1jrH8BkLe1oM/PL7+HmGKJf9GKys8R3y/oIszmTe4YqaO9ntqC/KDpbX1cTt+
mEwEg8E23F+SGrCPIUqnWT32D4kWDMyjwji1sX+wCHW/JCDzYQgztp2pyEpQXulJJUZcZTOdroGe
SEPeRJSzRfJZPYNcjerGvtf5XImkkkZzFoUeMqjTXzT8ZlEmG1gtKasT7S/5xJPvkLHj1HOoBaWM
jWJgK+mPOIWo82wYUDH2qTEb15ueIZ9MokG9uEh2GvZphJAeTneHQ410B76TaYD63TiHdBf6Koqo
2RvT2quFR5FplzkFoZolScEDUpUUt5L5uS9k3KJp0hYFSsSVa5PVqlToP71R/Vlf6+/XW3stP0dd
Pskj3TvuTv1l4nJlSd0psIGfQ+T86+gjGf0YBN5Ln/JTSXjDjXNCqHJPLB3Gnug6otC5ghL0ikzV
U0G7690U5CZmcdWGPETZEX9/rSMO8oo+sP4Hh2OVVYyzFH8H3iuRnEZDOSJ2zyeZN5HZqAbVHrf1
K47o39U0LEEiw6HV5w3oKdj+ICdhDA/ArDNG6ze0kFWJNIMEZIAcVyX2niuXTmTq8YCxGHl9ehQ1
xvAMOKvmFJt/EhURaAU3n+4PKnTGgU05ITFwL7xXtEmFFhwIV6V1e1/wPmopTw1vUeq88QpVu4Bp
36toi6YY3qQ7dKcI3uEDP0c6JMdefFx99vk2YLXb3OvKJTERBllCYKHPESM55iyRWHzrbrkGW2VK
agcRSMW50vTK3grVYzMY45NiEV7CYLT+9d5y+psCUe9e8Nuzcc6x05JQY6aZ3Tsz7L6SegpvQQgX
izhjsrvr/UOGENb5/aCImkyEvG33gkJEiKcEO25EJCTzxdhi+7f7EmwF+YgUdN29HWEDNuYtofQI
oedmuHaKBlnpug0mV8lQv4mtEeBqv8SLSRIMhr7hfLmRt9TWDmnHmyOEMK+sWEdoBfwtkCw7K0+O
ipxMjc9JqHDxS5TUKD8K7PcwkqBpPjl/IPRfgvBLpsnwwbEgKOgKZ0Jvfl6IEGkjXLxBrBSjWzG/
f8Xpm6J2YelMUGQifp2Wq/jUg7yy4YajSw5uPkpxAciuyPPsOSlEwTTkc2AFAeV8eK7WrTtU/aSM
Vn21t003R31LYG9fGNbSz2rhhOR4FXtGjkOaxelp/HuAIurF6BblRSkyN5gMwaR/8zABKlM9iP1D
maQtPtVWCh4oKHVi4TkBHumLJ2q0cgyn1+o3ei62BGmm9hxVM292NSJ9DWlPjDWtIsGbD5IsJ9ed
6ZZOrwHuwEVSq1xekdwVM7bZwYb/yf6AlNRP8Flr/SVI7PZGB7is1Twy2arRm18BBEm0gj51igTL
ONA8EQuhhchA0+3Ta06WGkxV1yolYovB8AyhiaVvYJqKMB/weSIaI6dC8M24+WwBwfiSzqOCvXLe
3Z8HKks936Np/2LheOK9mc6Ui+hMqu9p6Nu4n4kjngDsvvhM2NMFD3TneKmC50Jn2qOfjFWFJ3Qa
IQE6bYHqSr7CEvSTnOaSf5mutstSSD6hLsAhiJZx2SRxpLyblYAFgNqgUl+XHSxiuiFtxvJu9/el
vSOkBLQegBh/8ESE4UjFG4HFF1VcKIVBrs1eun7Yxd87EHzZQK69DMu5znkYCMZVxB37YD4OY8Sd
bKbxVXBANLJXH01Abwfozbob9Sz3GLjM+OB9zDU0F27AcTLb66pRPZLF/7aFOzHn+EiRsbkcDt9L
qAv00e1FddslrAytR2rzwtyKK9DxurUUJEaOGl/+XAXFPi99/NYfwHXzMJcJ2phVC1oDNIaKqVn0
VrJIBeVUvMk/gUyKHaDgyRgxbtgsrfYcbkSb+5EToF4lQC8dyiBzhOYjN5EXyju7q5aXS8qeUJFz
KZxCRgo/2tz+G/Jd/4e/YmFCUfsms6KvEVEcvrNOAGXZ+Gq1e5MD3e/WGkoOdEQl3ESHfkwzp0Bv
IDArxH0vkhurprzjGcxZ7CoCZYS4OiEoiD4xx6kf4EH3Se9AJZJEsuO39clSufJvBTUvoK3wArlk
f42EWK8uPOfpoPFlo9D/eKdznz2w1UbuIU8B3FPJNkNHslM69aHZdyoJjFp+ezSxkVSnhuZIvlHW
p8pkP19x8YJEi7yXlNMI5orSseEPwHb4ujA9jLd3zLMgqNlJOLxvd7Let+sAgzo92wNZfjXTwGEV
VzccXHJLMkMa9Rz5I7OrRNlzeZSbqQT/ZWIshIe3U5EDTEnNrJg1HEvPGEKtXUfuN1PB1/QognTO
XrTqWLSGU/lqS5FA9MNHurHrcuscymuIrvWkqnL8SyeWLRHTtTBZTdf586NWTTVd/MyRMruGV/Jv
Ch4JNx8+D8+y8o1wWnXe9nlmboEueHSBojRehs/StjIS12SmMBLG/A2tuCVHK+khG0zCoc9bDipL
rwC4+NXET5U7A/6H6nNz3qYI67y8laS1uPkWtN5379zKrVnB5plmXkbTbmLlFS74QCFBPRACEskM
/Azt3rvVDKPUWwzKlWCti9lAnk8Qtcyq+/+LHdul/KOJBh8ENs1R2JSvRS7UnAfZQx1YDHN0r5QL
4vg4co2mk7mXZf/XR7hzfsxG0JzuMvWcsc1YNGhlmun4HY06XIGLlXcz6/CtPnWPZMvq3cdZ/MD+
ihqlnDojtUX+GhPXA6kAA/sWrXD4JS/+4Uelf+YC2F8MmdNTvOJOPuy5yR/MtHU1AluAr8/Nxo2E
0oQJJQgbWrCZ1tBjRqgzthU8ImUhkB1nbY60Ei1wK/IlLE92Ottugbmg2ZSV9r8pNzYG68H+9nQQ
FCpfsfjKvxE4xL3f4pYHApCdalo8EdBhkPfHbGsf9ZqyBQLzEyNyDROfgkowHhhCeybacKEaHKos
J2iHVW7Rcf/ckb5B9gYg3UMT+WXO1d66t3GG2ys8sw1PYTjvftUKXLeyAPE0lCIZ8oThERXzAGrg
wEveKs+aqXcwMqQSj0vZdmHQsjQ41PP+zE5u+m0w/C2ZDWD1AfTgo1tnqXM2wyE43iwa6WZQMiDF
kCWwLNHZIf25HKTaiBI7TeZAG6nWtwTwFEv0V7C69a83+b8Pi42vtb2q42KMDE8uIt+3Tj3OorUn
e8dmD5O6MrJvcwcIaaFgOJhn66sfcWaMJ2yk8m84XIpS6m2hO9KVl4wE+GZueGsM0IVruvTNi60i
OZi/7GeYmCHtoCIYJaGouqb5XVOM5FatyP2qlJUlgCvMEXVIV+iIzHCQnSrE43PhX3WvnPr/H4/Z
uDyqxxtr1RHh65uYO7/ce6TcP9tnA2S2YGnjrfVjuGDrZFYEiPgAnLqo8p7Qv6HVlPGI+/X26u2I
XjE1s6PkSZAItZZ71NRcINfCanF63uT83WSooPTN8nCp2c6fLjhs8cSf42KaG5zzDsbdWENp6xC8
nieae442Upcccs1hDDglzaTdAZYxhY9BPc4YuKVTjmg1zVGiNkvGCC7ZxpkER7KPgGk1OxrPnuUY
jaPh6L5hCUrvniInifzmQ9VaGBkb9OmhVR9gK8s9R7YfnBVs1icHuQ/S9SAsCCMXK05/fwibjfgo
0BRpPxS9LqKRScuioJbnoMgFdv7b/855UCnTjh4oYp5iPoDi37RtffiSZgaBQXgJFGrQSfGGLGBc
++u1F0OkoYstJqNqnFYtt+RQH5QxMdi1jjapYz13hmxwP8fbq0E7shT9rASnvDDddS+6KDRXWrSu
mHwm2fCaFT+74dCXy9q3dKTTxbFaOhm18kfCwTTzh8LMFqqs+Rv1QsYkxV+G/rUyWxiBMgBR2UWr
P7HhY08AzvyEh/rMJlei87XkARvG+2PeavAf/iEQ0AbQNRQKNRTO6Bqx/FYRkGIiytAUwHugxhqK
63jEKTl+zRCUFE8a5D06Kuf3UfbZ6DlyyPew+xOPoWnvKS8mWuhHYhkbRxotz6zMeZK+L6pnORdE
vsV7absDWWUH4HZTs5aqiJYE9UiefXyw2eGpaPboxG6eKyWq+K2zNuv5O8thBwo2vwaVYbFEn32L
zksg6yI0JL2VgtOh6obwGk78ClBrEjipnqYhvoMeU8nOgTd/6/1lh1u7QALnms7jgdt/qSQYyBTT
IAoeSMvoeIVfrLRRB++nlLZQvibjIz0mwREC8aAkKjvYhSHhSbHQONlI1Ymogr6tDbk5jSQtMV7B
ae1B6bQNZb2a5YwqEq7VgMzLM3b7bro/XMCDnoLQqEKbtTNJqAfCVeg3jyZjlZkbeuq5aT0X6ysT
/j2UT81/2aLwAGPWCkTGWNgxm+Q3KY5MbhNX/H7aknEvXea+wJ8q0XUXBvXq3WFWEo5cDDIBaDin
Qoqfc6r4/aw1LKlxDtJcdSa4n2AT3jAaGem/kYzBRI7w3jbshvAANJvYDFaMF2uLZGW4LeseWvvu
3bEHqAVRK+EYeA4urvcV94ZqtZDXU2IDMxixsOsf3XltjEfptvvO2EiOM7C4IyTtz41Aa8XsPVLj
fzq5/lEZThgFyJjiNIrZuI2iDiY0zfEe74RJOefNGhSg4I8KlLqneqC94C8uhN2G/lFZq6dlg6t0
WesAGffQ71/hOzKuImDCmuXUaPYKX+ip03aZQpXlMGPp4zHev6AnYWlCt8JmPGu1s1dr1v6kQHQt
p/kUYVMkm6oZj69OTssqZLpiJyNsTbmAFaNE4FJEyZ+d9s/RoueCPqAuphF6D6QrmnKubBJAMJ/X
K4seObPIZ7UyGHuTGx0EuWuqn/0hmxpCXSZQMZXu5t7QUXVHFBJsneRA7lDUStvVeZC8N2DBtEQ9
rVMMNoOyZCC7BqIkeeI46E5OoR5CGVizb3lORCSrJg1fYPUZKcmtlwf2qxenSen/KZxW8ITnFe86
RQpEd1bmdIWE15WtEmBc8sjRL6at8zgyGWD5yD8lnQVX2sMhML1breBd+x3KBpEMIdZSS10tqegd
xb6Dl7dBLn+skIK4tdIOiVrelwuimXajuhYmvzCn3p6zMDL9YTzep4apcTf9LOT+ypRNbBBnULlD
J8Lcsg2P6u+uSF/pjEZPfyE0vudU7rwTrDsy3LB+CnoAXU4PyD1tWrLoJhrwH+5YpqZHCdf0r9gx
TW8EukK8lSaLzCXeJ1oSbAHd9eZb0SVBWCo/Kk3VfEdpRzDVVC1YyAe3GMbTW9LxovaMvCe4faTg
YjMjFYnMyh7PVpwSRaM0xWcu9Y0fSEhDKdns0r7kmCfu5f33RPBuuNlihXmx0cw0T8PCCtLJaQFV
dgBUA2qUEvNg2JozTf0QIyHor72W8p2gcls935r+L+ZfdN8Ctyu1qsV0EgbxU6oRaxM3OwDQ+jqK
7xXX3RIu7E/DU0RfwCoc+S/E8SBU/KL15vZBrkAWTJYUIMGrBm116IMilPesJNNa7POX5/xHKTIl
MdlfKvB7hm8/I/N7ChiDZ61NU5Q3CuJnnCi01ZR4pdTRG6GdEjutHoNab7x+x4eZKg+2WwJQzeEv
4eZ/8muIHFh1fJmflK8K6im3UpKMiBlGXMBj/EXnMac0Wd3fGqBxxuWAD6VkqRgzkvaF2ixLpeQx
U015z58eROgEXzhGNLxADqsJsDpIXBECw+h1xPXtE+L1bm804xF32yQqEAjYawRJWP4+Nt/0rzRK
3pYJVhlSlf1SW3k3jhP/GU6lD+/ytypfHJoQv99RLktz9tvrMJSjOmfUw1QIA4aV/jWEPDxl79cL
9anpHl5xtY3hdHP3XtC4RVfV9uPgbdJhDbF/ecFTIkFNRTizxoMk/soFWgxfl1kToLI8nv9v9RH7
BM6bPc/2q3HDoGlYH1f9nOkvwiIr1udXml5iLsI6vWUQk/trbSCUM+nztfoUGF/N1ilQDC+Pspws
6Lj3iKmUc/z7zhUlyXMbHSFnWK3KdnCXI8K+OtuhwzwNVBv5YqIi+vVYZ0/nB07NbIMjwutEI2ue
4RTjWCBcesZVFzPzKfVRfxSxURSfMOqDit3ZNIWyDFJ+o4hhGvTSRJeqn12rVauBYoELPNanBy0m
R/kh6uNu160NuOFQWpAs1MmkMayDKeDzVH2Z8xZQWs2KCIviu9FCmkRjFCMMTVdWFa3dgNgq5h0f
+v6mC5He4faBV6EILGTJqlhWEcTAAzDz4+xZCfBiD2JvAXqs5Q4bU2MNobz1p4Y1CjArOVeGl+Jr
CiOy6LCiEF6xyDEczuePGiZvAdJCOXQnoEKXEpGhlHDKrqK2EZOlhePMhAW5494pwoGROc5rRNvV
EJ7utaAXRGqYCd5ZY4+Q/X9NHdsNtk1oSLRjuUat1g8Q1tUHc3KyQHMRiDDGiJami6cL8vIOn3J2
gr1QzARyH5N4t2Eyqii06iSriqx1/KqoYDSnBTdpURqSxQy0IjdzPmZ1lglIhkp//bgO5wDnt8Xd
7pXiTajuvrIAh67ca7AkVjNoP8isaTAtsz54H8mIsvKNvCXsHziOGWiHOULI9CPDSP5NCWLLtOVL
fE8VQQ3MVjmnfPCJkeWZcdQ+0/6gv8ZQZMo8ItI9k+xGJceifXUHGJqgGu6DgJlwd0+uO9nBAP5+
aaxHWd5m9jAXcITB84N/TK8O9UpNDNlWtpTgIK+lTNw6p7vS0OpvMTeCgVFYRWXftCttDt8hLzJ3
2Z8q4231WaZAm7kkF+LgNuIl4yXRRIV8eTDxbLbDlX9r6iF1dka/UDE6kJeEX/LYFQ+AN/o+/Tw7
P44bh66SaGZjBsl12b4m3nTY2Hu/d8efUI8SN5Yej5PR14jZ7XSKr2luCvPBgUgnZmhIHSpDgntj
yBrJr8cNIOoWBp8yPxs4WenwHMyXdK6rhRyhExAVdA31M1FLY+U7MW44nG6dnUx67Y7ww1LbW1m6
XqsGUR5yQivvqUVhliFQED9+/rP10PLkku0jn8oEHetReVQT5AueSvlucDIDynm/yiiEdqKgTI87
sV208HKjjZHDKwq7roLuRFqFMQZ8lZ0SnesCqhjeHKaCnmld6kagYwvDE/F1prAi8TvfoLFbr8Sp
b5gl4GDBNbLvEa3e/OYCjLQPKROdgj1HdgNsOZ3tdZETZpZ3upGM3iCLbzmkMm3OaPsocg78p06T
3tsHtcDPX5YdqJDO8IkLiejTUou8XIOQVRypjAduEQqABZQbxOAB6tDc14odI/UUgRPJpMCjB5L1
f4xiY3kPRUlg/zA11PohJQTNIHrsjh4XlZ44u1m5Q+Al0g4PzAO+AEmgeKJs3mA/1V2utnZBOq5C
MzR0xtYcfxiO1DTW1e13CoZ4Bo/BLv8FcszoFh+kE5X91dNLXqQdub89Xbpi0tBL/DePT7IgD6an
i2ZMqHBk9YlEn4us5edc4//phikxH9CCK6XFoDAQIbNh5W4ysRYfADQRWJrcTCirKUoXJ058lgMp
n197+FalHQaezSU1hYYDKDNqN1n9BmPQKZJD9VJ5dI8APUYXYvrFjVMDnn3VYh5cqwOxWIWu5J20
BlS9G056cggB8QZx+OjPDj1Sy+jvv73HWTPiGiIhlAaRZuI7stZPk8RPqzZwV9hdakvqIaaUss1K
0KQtpo8Tj3wTTSkZ5rQvRDoYTraBPI5/h2trNu0/R57FIdhn4gUq/Ev5gXqyC4nL8Px0GeA1ZFfY
qmPKx0rY8hnvDMb2jfzbl+YcmBkC9wDGDewpdvfxFfRZaJgbNqeIRR0Om9+P+ESda/qOtjQ0eAEp
EDCAht/L7R7YAZhKSHh42tRsKmlYiw5025fSdHH4+frWJHhipLT0uX1KeIIBvru6274jpdXoT8c3
TmqF5/WiwdJTjtsxMFZnS8cw3gLB6jlXvddzcK3SFfAQzuiftbyerryrkyPGSN7P0wYT0EzEe7Nh
95dgjUISw1yyOJAzNzFH50ToTy2QCe74DhmR67Sm2QwbipeMyzWUvEYXrtR9na9hy9PmgwGkCRhP
nFOCZ/IvvFGhn987xLS8qs8tKhEOTjRdUGBlaNJg/MDlL7j8HTpO+n8ZHWfvjRU/BlcHydVGpUK9
yYUdAG/fZ+71s/vPVyTvJ6Jq8PfdBEAq+9iEFSFOZUMozfO3G+IUWVbwByg8/FLWgSh1f7I+NBFU
8YbuTHFWC+u2blstaGe2b7k+d/GPkcmyGFFozWgVeAKEhlNGkDjZ94b7PvRZGC5MrUNk0FEp1NXb
vB4LumVXVxo9xQKdsXYRQfPCIJFXPjcr+2ZeyzIt9uqqjV9c69W5u42McM6FHGzGJO+KsprjGs3i
Uk0WRz/uqftDahg6LJo77lgWX/xDZ16DZMFQsYYgz4623bQY3EJome0uoDm4I/6dZYatZIIzty5A
4mF9TdGFhYJnCXG+GetoztgSe10Kr3+0o3W7vaI/+nZTVrKWRCaKwo6HQ7i+ip4aSJnMpQmXNmya
oJNrsaetKB+enmjvWsrrr4tTi8ZizrxcLMtkNAmxxL2I8SETtTphrgB5MDL7UCHZwLix6XtpIAnq
T0BCWbcwn081J784nJsahoFIVHHMzRg56mNlzp2XYuFKYepGKdbtux/A9f495Fb7cUqjDMoei2He
8RWYNr7G6i1To42F0YnD+q6Dvlxx0a88FvmjKGBV0aLicUY2fm3+aclQnCOWamHH/5Js7Z77wU6E
8mhRFTcINLvOEsQAc6McP1qM59BJxnTZLmSIoDZn+IjhxhnSumSioPHuPW4gAtRX0rxuIA/35XbK
s37wgmbxyxPuG0ds/xfMp2wehAD49y0FyFgQx49Agdu3lAsEThyd3N3FMfhmbMIBNHRfE6mGer+G
eCId9Y0jV/LtZDmqlDKCc+Flui0Jt1geRcE+oBKTF2jXZFMXnhl4brr95Dhy0Ai1KTICPe9kdrA1
XJriqC2/LweAb0GvfIqX+tNk3mwW0LFvraKqLT/aSpRzEZ4W+A9P7YUvDtMAwbntiAjpg9hXe30x
MOiDZgUlEugAmW5cE47Ts5UsOA71WIWszH/hyTorOGTqNeZXaL4BLWCyZYLMDi9v8Iz9uu5i7k1Z
S5RLTVG6U4/KS387mArqU6OaPXXomBfOZxSbNDv7hlZS7GpXgKEW/cxjPwB54nalGJW6YjwAi8Cd
LXWlBGbXsMfGJzuNoIUJBuJBU8SgwAkwJxcxBfx+MBKVbNMgoSumRiP2DdLfDK9swEmQFVU/pkqd
vSoSfLQuTLmd65tzINRI7DHrxPjsSKcj4V6h0eofPZB0IRK4OHXdsY/CWCX2iQAfh46yRaseGHgB
BTV93JWz6vtohR0bTx0IiilS+FwGjt6h1a27WmBJnWar54YC2gNneE4jD/F3Vz0L3Cvd4sDGMGSk
BvdMO0+uqqJf5G5TmBBjp3B8HBK13+d3FJe4NS5EcwGzJ6vo1CwF7PaBD/BvfOg4/8M5Ux17nBia
Lz5EZTgvhf1dMHdBtSc3cXU+kFGT/iI+JRr5zCobFeTNyRO+RlYNyeHwpL18YolpRRxG7xoDAZXX
mHZtYsbnufmp3qxlmApVXPF0otSqFC8nJFEVxX5q/ZPh3XC8v2bkK6rWOmKXFh3/IAdHM8ZpgJE9
JJ8URao5FFjRUxrH0OhU6TfghH1ga9Agr8Q0+Cayg26GQc49YkFqBRIZqzDRhY8hMJsyan6fY+5m
CKA+m3HXGfmkR27x2u4IhXqxFIYrQI6L+uoMOMSHiNQ8VdUIV0OTnmm75vHMZwqd37RZSQv4+86O
Q3jq31NO4Ex2Zr9Xynvn19KXG4u6kaawLnSEh1z8YqYjQT3MeWKP+brZPBGBI/xxN1/gVvuG5U7W
bOVyiCtB67lTWhZ7O2MthEybTuN41vsEVvyl4VJu1uaB+zrnZQZNDJegZQL3kGaRrG/aU3JGKgp0
Ck2l0CXNVw0Cde6SH0awKPjfjrcYbrbVivpXx9pswVOaUe5scuf1w8s64Qh5PvfZ1sBtDV1MiWLM
CbcW1wiIsoP5Ti3zpzFw2aCuRFNNPLCeJ6jqeSanJPj4gFDsZ/Pk/5l2cfBje/bppnUI/6KRdO3k
vQXmt3/9HixKXxu+2pXZZmCXqsO2SgtuODRHgOuBIkI5RPZ6kZJbdpEXHRPZWqtTAwYRZ9QDsKvs
mWIn0KsxqxQP68egIQlVWoRIoUEa1M94sTt7n0tMl70RX0h8XYXcvWRWNVFv3PLJ8qz1n/5vURCY
MFfz3xFyrZ0MWacjamUcyeOXTnhqzGA+jDLZnMrmrEyCiqsLCYfZP1eFuAcYgn07ttCDrS8T3cuk
cZHIfdod4IUf1ZlE8Spi8fGgwlp1ekOeHGyJ5jiXI55Zj+EF3FYjO3BPu2Rk4+LHyFc5pky9ugiv
8xpylWmXtZkL783S712XbtaDwfYgHu79AlGoaARRndfhEEzb/G8alg+C/pLBKkK4FjfZw2tJoghI
378nqh/ITFJ7X7in66J3gDNytMSidw8cL2CKtJtB9YTgYlA7WxyJ/XpVoyFIubeYpcAqiJObzrSY
dgBUYz/cffOvNhFNPKGVja9w+M1GC3OHbQUnRwgsHjUPgXuEH6kXZvZ32xwwfqXiu9E7rPZBARM3
aseLmzw4prUqq9W9VtvGVspKw75hQH0HTBT/9W1b0AAD2c2OOm8tG5pjP9cTlQdRtqfrwuenv4hS
qE5A4E03fJ9I9GNGHnIATVmsGaj+jBQSZfXGzayBii3kFJMTP/39bUP/Tpe4ogiirX1Txs70U04b
XixUZJ52YBUbYVq+Js+aULIdv6mNT7QUEgqJK9yuHbE3zYFTZIkG2WYQbKyuUTZexLIr2g2wui6G
xxt+6NowPadvR6HBW3kqPUSiOy5nE8OLefX/V+X1BguV88bz4vVlaSbW2yCEDNvmluKjM6aZzB5l
7l4sn5vOMwf/z4jcr0NgNsNv3SpPnW7kmIMMUe0JHjqSPOdqMo1UsrEPsPcZuaalpatZJciyA2UZ
3LVZ0+vG+Dgkkp4k6583wwwqpphwQgCfqTRLJv8HsAzOhw53tglxhXFm152rI9Bw6yXXNu23ezYI
dKhFkDV+wIOdQnQfRzIesewbGKelj8yBxzUuXHvRskgIFTMdQ6W3EEfe5D41FAZXDXc3dBXnou1l
5YWt1dgYHHgRI/WJrpUSDEEaECWR3HcQB+3v1dWXaEkx5dqiu6B/ndojUP8H1FY5zd6t9eH6cf/k
3IAf/4EXJIcVLhIqA4KfcG1mkgI4lGsJfQ+6m8iKHzaNQ5qU7R+ZvrgQIfmwx6qaHfE1j5qFwMJO
7gB4nobViommytgZVJJTq6G0yHJ2kLbWKeIxEQcsFkV8aDmAFAPOVyvT8C+T8TK1DhB/Viu+KwLO
kNkedRQ9ZlkS7jh93pzY2BFiQNZVgRYyoeb91ytFY9VwBr4ryz8Bjo7bo/cRRmRPQbGfr1XJnZZy
QAhX1r6QPiMxi3jw2cLI6bOiyge686v0n61gudf8Ry2saWChBGPOoWqmgT6vheF6OWDIC7FSV+of
SYroLwHAtJRDzk9MSySnJiwX5l4v/0hltmDgkx9F4US2THVgh9B3CCdLKSt7PSCBgHhqH9iKs5Kh
V0g0ff7F54p8Wkgjg5e+D0EH0SedNrNYU/R76QWFgAQRQctf9EYBA+nXzv2gYn83XPRCsQqNKvKb
RwdL9o26uTokblyEumAuOGs9Q4Wm8L12+6p96wDXyqxZ4rsnlPg3bx2yl6tP7q1+eN9Ow6iJSjWP
gKpACUaGPi1VA6LlbNtBxpyGNTeKmwLWpeJ9kviEe8Ww8R/xGGkBAWTGOVKwOVdcxO57sHsVKHYL
uXPqZjEW+GebDxK+fCjvw4gfPHBsU6wtE16z8+QcEDl3v4baTsfBP0ybiqY+tgYSMp3e9VlBntwn
SmRyz04OHb9YhD/rrutPltT+7PV6nT30hpfg8qhyYR/NNGV5ZHr2IAOBmWFASZVS2UfhZZrcVr7o
qmiUlmJgxe6DCOgl4vTs2Xi8J2PLhGIYCcsRd/VmdM5MW0nVsqVlIh+3tYn3eYT48IL5wcPZcGIX
Ci+478GVpfZqqGvLqElosCxYB6gd0xNGE2kZGCYefjK4owKWzQ4EY1IjXODYOCDIdx43jhDpgHCG
5J+fkvObowQrJ1KJVHfcj8GRB5kQ76F3vDHRJsXe/2sSq4SSmFULgDlnQ05w7EurL9Usy9fHZIuz
bkODrrwH3EJIshLDD0/ncd/aFB7ccG3tzt+vq6Lp7gZzU65jN2xTGUELsXv6dmXNkNh7JnxZPrL5
DvcPnrtMwKc96JCPQSBnIdflBoBKP0BsG28bLCLdte8oOML2vkSPLFma0Y9zN9mLhlDCYTciHmFA
aMxaEhSVwb7R7aIr2tq/Qr21k9Wgdh4bysJ5txXBzpS+e05JG58nyk/s5+gCDcirRsDNM4AQxx+L
eVcCiERuAyypWIDY4RruMQVD38uvho43rxNDZL/pO9qZucLraq1lhN2DD6HUHcMmxMpmwTcuiuLM
dCVZ4nzZd6w6AED/ezM49ZFP9NMLo+vOY25YsO518GPUWAmmsFLk9/fDuCDdXfH+Y6no9tqWTwvx
5bNlXaJYzPNXAsVUvwfOSxJrAsIo2Fc3RwGQfLX5iM2bliMSmcEtg2FV/aDSraSdFBgTFvCJTlvw
LVx2B8tq96KhtYA91jjaMs7rwcaOeHkUYL2qg6Gt9m/bEzyd5QB+BHg9RMOq76pcL4ypiD4NZcPK
jtGndO8ogjxInUmt3/aIyE33LudkxOjuTJWxzCTxvbhlYasi2w/uPecmRjJjEJrOo+3psnzH0sCX
7yRDqhcVybqrdsUL/VMwmgVY0pxbChpRsMQiMlE6ir+NdYvJIiK3waI0Znq/oMF0Y7mfuV67yieO
ZKjA1zybWB1ZfRz0QkDtYnqQvZ/iz80OmuKUJGt+vfr/xyMhuzS6+h3eEabxVF7MxmIGncXTv0Sb
1PrdJctVYP0EmvGyeILMvEPHnBQXP9ua2krgXJWQkRQ78PEaq3i/7zEXfeA8/MqCMucOjMYg8bir
lqGIRxkugmqhmnwznlXwh8tLdkhPnXkAdvwRoJijeWUv/uCQMGCtXHWjTPo4NWkmXlqk43RnbD1M
13DtzxI73rOxC442b2uH26vGx6vzGdEao99ALWmCXfMKqZ2ZE1+XzH4p03WiTOuo9RzfU1KA3RA/
9uUDLOf2eEAvjDDb7Y5WkXJQbIyuD8QrSlfItopH4T7j5AzWik3BWxm0YxJ+VQteM0NUPC1jkv3i
0vsbR4Q3CvItHXXPBaTDdQ7zwkIDcYR6Y605vtmCyQVU+Wut0SBEnu3zjEFS91AS4KlDuiYP8gvY
RHW6Uv2mGBrkNtLZsfQUy3Cd7gCdgyc733ki3BUCbRx7OBuANsC9WwL52YkjraDsfLckzLMJxQ7y
K4MIyqY80JLWObrnnYHUwpTLBNFXrRPjDoVcEfzFg2da1HLjwgBZguBjTHoAQ0Ycgpd7DvAoGg+/
PBSDyp57JRD0zkrD/Ebh8zXZkQ0Qk8LK6nUTa4ETJYQJXkId8+eQIUamJ3B3nCGfwEyuLGie39DE
iYvjjsjkKzlxt8IF/57BvuuXRJrmcFyIVsoGSQLhguEm+UU5Fq/ViZVFfjUTHrgrdt8a8mARuSD3
BaodYOEVNuCRPaaWWFMJaXJ3z1F8NK3xKGI0pAma8odT/n0VvO3tJmNl4bKqYEKaOwxWRymzxsJ1
u8hJ8eDzKckLGdj6Q4Xwpdc8vAPJ86UUzRoybuafqnl9yKrm1RPnkuO7gYI4GcTeGNZrgg5rYR7U
CEsFeX1GHxuEboqwI2m2RRMyRCaeTG88woGK0JcfyQ4QX4xfBqREmtvzD1ivfirYQCm7LBUexaMN
9Q2rHHjo/nwtAACz7Ugt+wPR9m3UQ7ldhha2eCATqabDkblleYfZMMjahn1Xb2aBrnkObwEBnsZO
p4s4VtLGcmgaPOYPPn0bpX5pmeU92VUjHPU4qU6iI6BrEBJLONOIBOtnD4cjLtxhAHGGOKs2nPtk
m91cIPPOTfJF07UHaLh7wgKTPUDm0RAWkW9lj4d+9ATgSGtH2p8SAOnr80VXeOaKVLBteldrlmiB
2YmW+oS2FNTi+D26EaCw5ecoUtzdG5z7lgm4yFrFlSLZEUFEt+FNjRclRHwqF32lqaSijUW2U0RF
/yrnQNMvfGsWpKQSgwNc+AH/oDdshbbqgJ9Ehab7N8Uq9166FRv0tMf2kNFyh2QmuVX/l5PF/mSO
7lHcqRXnNxIlx1BLZsKPReo3sQSOi5u4ThRKHKdQZiCLcpYzmDXjPZ/xyQGKe7b0Zg+Vgwlo4RW4
yfqMVzWOnXA7u5mmzNU6kej5NphThcb9OMFMZKcqPRK5izHocaAhcp4uidJoaH/oTkN3iFbyL2Ox
miOYQbjxYOb1veMeKz3G3iX+Cfut6F9pBOtAdhD6av+Vzl++l6tSNQqbfan6tLxgWesApr5Wru7t
cwwy5/QsfsOqCXlOsT5Dq6lNTVB3ClB/7cE5uBgDhhPdZTRhDid2suitN5uYPoRgjYvOaOIKBPqG
9J1RT2WtC/qUFGpcEZ996aGZjNWAA+opp1cLRBIt0N5c4gTEGQxGWQGYeZy3x9px5zovryLhL8WU
s22wIFtlbiygjfMVGa0BhQwfkmqUzC/to2c4y2ZMLeGdDGl+VnoB4kHC3/PN+XDXo3riKorOWfVn
UI+TUdGB8U4CPxkyB0wKHhgThn5kVAzQpZkaIWGSB0zZG90vNTif7xXfGvHKfXWK3DGWgEP1Q4Zm
NwHEZbm6/vEkK9unNLDcSMBPqHk0nTUI5MtyuiwF4SN32IUdpNX09r0zJTwIXA8FLGxQJeRq4fT3
ukzs71KiaOPb1slVn3W3SD88Va0Sz5PyNxqBEqi7Hju9eqgdEcqbwIYtf25o9bESxKRfqvLqlg0Z
8rgy1T7CU+FAKM+TIZMzrh6l1fK4IrcMNmzXvtOycN1hmJwOvbB/rgLycaS3OkOf4FDAadygVEpA
aUjHjOrtcmdutAZgM2oRRVHTRRTmEkbdKlYBeKL+50/Z4s8cZfba23YCPJ0jr2LGjNGhEZuHgxQm
GIs84soe1lEYHLq+f9Yed7sjUM7MtguXhJWjXkGBcdjDCdXgmxl6kC/Duwvk/05Am65IvES5rgu2
t6929fj/RpD7tEA5JpdFfDzaYydbrvk8UEWwtDMsbsUik31l6+Ax0nu4yR0AJQ9zhx2yds0kTcB6
+o8ruOB4Zd+Bkpa7s8is/p2EK5XfoD7nu1XfodXSvWqStDLClqXWFP45DUsoaD3FyyzYaXcY+U55
h9vD9YThYLhYAqKXxiuWu0EpdIMfNcWbdadCSn0LPskK8e3NbPnrEpg+DVPD6/el7/681zOGAqby
sn9v0vaXXxjHVkfbXJYjXDKubfLO4Eql8ZIvbSLvc+tX8qBVUf21LFRSjjaaDVGsiv+jzStCtGI9
0Yo4vY5FMncGFwg8i9pG3s/hADx6waLDi/dEDOEWYq0nqwY7VXkVTWq79hEul23Y2ir70clL/bLF
I5vLyFRzsDxU9KYu7okAyQhpOa28YJPh0AFvCs2kDCppVSWvIekku9EAcq/llaCB6nHQ3t6TNZ0O
58v8r/gJx+iZd1SqzwH0SbdIUmwxlja9HP3zwkQXRmFk/icIvkP1uyNcQgkmW9L1w5NTPlwF2Xnx
NSer+E14pFoPvctuk6HfOTwkkt6luO35kcsuxLZasc+wZ6i4p5h4vokZ1Kc0871+5Q2B7C75nrwL
2C7gtd4AZAZGLvZ+3g/OUIe53mptLmXblIgXI/D59FdToKSsCPKN+IKncCX/C1x/JIhLxunLQt3w
9rnKzE4S4TlVas5FwCAE58ffamkBG6wFf3OwP5M6bihHRItAl3HSnSmYu//IKYh8IGQKvlWyH2c4
aIOGy5aFqLct7Et0hUPI1jomyTcVdg1wWBXKU5dl4Qao8t+CeJzMUcNgntybCkBiOR/Ckc3XpyeI
9Iz8edTdUjDAlzmvEFZXtveFnIUoBGwwQBhVyHxnNILBZlOpDsS6LKsflEL7b/CX1goqAMXvuvaJ
pmf8PoZm1T8hBhVptAooDRV2LX6DgxUaG3byGpumR9xF2nMvAA7b/BL+qCvW1o5K4wXT4Pn2nUcP
XjKdrgbsQYTx7XxJu8ZPV9MRj0eIeaI4TVCaX/NSyU0iiL9VbeUuGSwn+1KqS9kyKjS9WSHAzke8
9TMljvVbul1CvFo68rB8ppDAsjOTs3zwrKA26MAHX5O8vbyPNRxTRxlqZMRgfMN1mOcLVtOCBhr5
m49tUQl53ovDrveDE76nRMHpqbKWJh+WLv4Pi9SUTOWg1XcD1JrrMTfiWSRa4TxZp2o6mdrVDQ3O
FnqTJAHETLFq6a0CAryHp3IRMBrbSoMb5g5X3TPdra4o5IGcKy3U/5P4NQWqFS8bCZpufanFWLYO
oy1F6yx8+4h7hXsXQGM8meu3v18978ooTpmuBYd3rhgS5MygC1udNV36MNmSD7j66qrfGkxJk8IV
KZGb4rjiY0+aXAhjdmA4ablon/yeyypN3hITDD3hWkdMsM4dHR2D2m064V3kTYKpftF1QQ0yCtWf
2bnDMnyQxdn7d4jmhu52s6hdSOsCPqCOOQzWhKa2CVCRHTtKp89jCs0hioXCuCGO+wrIaMXAQzy3
YZhS2lz3zf/dKSAHGqr/GB5kAhiki3K2EauG93UuApTU3GdoEFL0CfjQoov4jh6DqNGAgqDx6kMN
Zws6Mdjz+eNff5WGXI91n84nLPAdqfwg+SnUR2b4c1RFJLfh+HYGwOtU447OBz0oRkWTbK2ZYT8w
wDBXmn5LjLqRD6I5ctGZlvU+bjUjZsguKvXqVDJR9HPabq7e8LaO932xzqZs4/49HEvw/j205R66
ji3Nyb5VH/wZMaVKDRBmDdSBtzoSW2sHbeMmx7XzcfdVB8OevEJKD7cpuMgcz3NTQdZMfHZ6VaZH
2wBXROva+9Y/BFsYeBLKF6pONajXdR9dwJy3nFrP2FOM95McEOVGR6+Er2tHsxKhz2RO58XXy+p6
13814r6Zq7SjdEoD11yuHvIegk8/FeyyIEzaYj0U3AmEyIzOdlP/Ika340Y4tzFEps3Ifj3TmGUN
79qkaoQ0S7XYyceLwIhea2Uns4xn7EWRMnuWMNGbfN9yhOj0uyJEd3WPZbyqM/EugIsUETmyK7Jy
wCG9sg0vvjjntXF8kMnLTHTCF6bUS40XD41F3OOuPucFA2JYcv9eSnKN+9slpcDn8Fbt97EYRlrE
sh3h7mTS681rSKul4Q86FTsOfWnEzI+antzWGm63Kkaz2vsoCSKLzKk2+JejZDFM6km/x6PUh7Fp
0tJjVzgwNbtnI/55R4STKvLnOKeRNv1/+ycFwF7EUCqglU0m+e803vZAOqxOaknfZOECK8Z7ywP6
yCbEeH/vfpxCN3CKfRwnv4Cbu62EqiOgfMhM7G7WJNgVVWTCNPLh8DlMeaFoW+d8yA1df3T1Vzm/
6VOl5WqhOn8cYG+rY74amYLVt1scuzItbXevAWYtH32djr/zMyMn5JbvaNJeP11eke/YXSOCd593
TTgK5v/9abuaGE7Cd37lE2KqHMzWq5q065EkGTZDwBWx95o1GJR5w3KEkaKXbESJ8IN0a6hpEQBi
yhP7ua16rEiGcBGCQyozljtOagpOS58ZgUU+H7Sht/E8Fra9GokfZtE7mq4pnLO2SZVUPj6sBV6+
cNbR5HA1FPdrlrFIETtXV73EuVV5CAcJAp2SZOnr4jvypTfDi+L16ba48IkQEoUY5xVqSrEcwDmM
vVGj1+j5mSG2GyTihp1GlhAcJWKB5ih7GjWLJ31s6fXeGYISU37NafaTz5LSUiDWig0FcT2pJZhk
cDnpGSWT/VqR/ECn7BDzXhNsrxaG4Z3axpUlo4FtOilXXsmuLdSBV3LO4OEit/mhFbDnce/m7H0s
m+A6hLGdH7G/iF2zyzoawGBElED3JAQzT+L4ahLLhU1Rss3Si4KGC/mXr+nadbK58sQ5wytGQSK1
uF4jmp3zoqHd96BWsLs8Ii5qPX1E5X9mvkTaKodTswZgkFiQBiZx03d0I4lX8EFsQdHWS+NvOa4K
jEDSdDDdmI2SWLxtDJz5kjtxNUc2etdIkJJDnQgNTfKpxMDo1BvHs/zFrjMMqppYQPRvapl8eHjq
vkrSJG5q3AKTH5LpQ9LOEkVs7vjzRU13zRSvGFPo++h4+gck40BBT+hxT507gvlXFK9IYeJkaY0Y
IPqft3iQjT3hNPZUEsax5kLjqZlejtWrsbnWJR35wYLrS4k/V4GdRStq2Yge1ijlbjgoWx17iGhe
CRU5uZ3DXiJY9emH9d6ay/MXO0XKBSmWXFMQ468MctF225uL/Vu7YLDOhIteyTeVSCA+X891onjW
yGMPWpmJKFtJzWcMWEjPYQvu2W3xF27mviSakcmEnGQFg5yPGC+Tki2sJqcdXHsAP+q4ltEPxvkI
NZ1iGA1buthmS0Y4Ss9k/18Bn1D5Hu/5O2OfT9y8Iq6Esd+WLyJGOKO+FbUh7EHSxgLo8nsKeuk4
+EHxVTNJYchlSdCXBCM7eDSn79EmS6DRyF6vlVHVQAJjVkUR2f7Lcbi20E8+OH7sP+OCAUdcNJ7F
RnEnaViqAR8MVl5TDKFMxKp9yTNnbgpsolTC7VkXdMThOnlCSHwLFIQNklw/SL/NaqoS1GefvbvY
Ufek32paHOCW+O+p5KtHqscXsJcSGVlyd3JFIZm1ot2tMUJqgBXsgEERObThrfoNnjBpxtl+xCk9
O1b1TNqnhQ3bMgZAnq+DsF5wShNEydx8cCI58xCWweQORBAwhor6RS6W1WPOHPhoTceQ1I5JbCBB
oY2CbvJo6K9mFdA8t4QeYjibcsglzv2s+JBaBvguSO+j0h6sAw0BNeYPFrHxzWEIyo0bh7bBhiw/
1eZAG+808WXMdGD1wse0tnkuos5bgnsFF83Sbbryd3RX9OeT3cXt7By+ztZSHInwvn7N96Odb2dm
99Q+/aNbZ6MpaWo70GbjtFPqY3iiCuj2+Wp0SEZUUJvxkWWtndtOs6LxYspiyj77EoIWgDi/cdoV
5JDuteGRxowUced+hJTFZgGWRJ69yvJOETm8VtGJEx5CKxcGeEdnyBvH3wJvzwBYAMCquKmn1Lig
B7IaAHfXLi8zRyxBPsRJ/3FJsBTcyyHTQ6zoz1qZ1GKOaHGSillTe9B076Ij4uJSmRVJ+O+0lHWP
8D7JRQpHHJycuV9ZO7aRCNAZ+YgEIW4IMTgbg4WZq0qAnR0sWeHGLzQmq5XlUf479cF5Nih/1EhD
g6LPaOgmv+o3D/6MIb4fqcauLmawwsj84hoefhgRR4y/fB5JEKWTmOsBT2cf4+qxJtuMCWQtr1bI
1bZjhlk3uUqUIWh+M/5LdDEF0m6XKJZCmwd4f9pZtxKjYuGQ4Aj0rWjIgovKBQXrxl0mbAPPIqOw
k/IxkKV1/Qp/o9F0/tl0OKT4W8iEUAcb/yEFZ4AgHSMJq6dCaxNfqRrNh+z+C+6tg6/56p4VaT5Z
2T1XRTPLZZoOLxpX66bYYGs7hS0kbMMYDN0g5lwKotZKxjVvbsYnBktg7kfRoFfIOnqHiWxHvgeX
QzBOqNVi2Ctym48hQcIrzRSGQJ9cRopNBYzafwpeDtXwZeGYkzrXlpDerNGl0VVm4eHcPdbPk3n9
IQzt07OuApAfnV+6OxNqXpj+OOj1sPuANk5E9YV6OPzoaui249FQAtS8A6/1vDvdlo+YgtZawKbm
H4Lt4DTuFwaYpLjlaDJE29dJdwWZs5HixnWeqrRznEjrP1G3Sw47aNdlVamQo7cqT/ZkoqZ46WoY
/l9E0JKCeaVX1sZxmA4PZAcatWTg9k0nCQD39tWY26tE+4ABmwMfJTSUrkkJN7CV2dx3VA5055MX
3fDq5irV3wKEvIKWGBVUBvOQnsZGvB4WsQKeXOmL+cT4mSPoyAMppAUgo2G1bjUSrt1IDWSNaw6r
O4qIux67MS8WfYhrj7jTfI5rUfy29oturLP9N3UEk15+4SJ+pu5mjxSlt3th7mrS5WleCJ1VuLbm
1DiGNTBtjZ79NL5r6k3Jbssdr3Z9ajBq6WT1KGnS9+5J2oUxBNh/2xU4evkX0p5VXNjM8wBxwxtL
R5KuCKFW+xaCS72uHrS7tWFLzeAk4DYIC0PICQVTFdhXw8InturOACS+I5DwAJ31Xl3ZYyQ6JCg8
sQlXoZNicqHUgdFvrV+zCD/ZgGaTafFlHleqffFrMSln4yYGdjD3n8pH3Ubks81MW4eGapm0cfvf
h8sBLA/RMkTNXZFbilo/j8+sUDb6hn+tyyPk76Sg+lVB0dOzDxWDdF6hkCBWCljHcLKE6ucfp/Ri
w22PZw/LKsZd0dL1+D4HarcOM8CpaoZjC45TGwPBKLcqYJB62mBA66z1O3xOrpaiLY40NlVdvG37
mL4kh6LU3cQOTA8qEPMOBh2xoqeVQ6Eph/DNUwGdUPU2oxZfLnoQpoF1rJYG3r1oSxhFZkXUVlgl
b3CU+Hg4preascsA8gHAPxW8WYQP5VTTA/lxI5auAK6K7UG8rU5YpDJqCS3upEzJfhXx6dMl9ZmW
mTCUfsXNSCvXfyahpv5BEFeRVlf8aLNNtnF2V1qchO4Dysj7Q5Vkrt4zjhnRIh9BE3LMrH1Ym7eT
h8QTfvRbIoyuIeCBOWMhjz2apUG2mWnmREXCoUCknxpanl9yDl8JjxkDtUsAycUMufG0DlQnpb8P
f3RwhHDXfyLPBvxc2JNPc+E5YA1e+suo03kZICuaoRpZfthxoA1eepUXDVQIY4Iyqmjt13N/E1Vo
gLU3Q7Tn2ePkVoluYafs7iuzv2mxEmN50xFshGZWA5gUHHIYRnPr8IFTTZYHIAaWkoX4RZyXUxPh
x7lqEZLAIMmqHTy19d27CV4/GNpCu9GdbMrt9Ao8quSsMiSapILxU3IbiATeZYnUO/W65Ytf9Tzx
zGmKlzgF0KH/P54dicFwnyVDZsA8OnrPHwLrhb1+K15hAfLdOIdwUgNiXcVK6dCEzrNPgNEp9Ws6
wGjC24fgVi5l/rZqoDL1eLssyAKaHO4f8+5eIniB7x3N7m5EPS24hd8rfDweILMImoCf2fGi5mMB
tBQ9VtBRKHKoXRA3MPlBglpUsbuW1EMYW6mfcpbRkJqf8qHcQgM15NT9JNNZ59eZMf6DzxEGkgh8
w67qAVO30860fY4CWOOq4ahhr+Yu08B9ke/UdOrIHlybgoq/Tc87JSExTeOeuCvo5Sx2ydAFHMWm
l6i1GDW2qDBpMzLGq1ji62aXXdU1f4J+rfVwrZpcG3TsI58bW53LxkQ/E2J7oMLiLW8M+Ry4jHu5
9NRdY6EGSIHuq6lyRP9QEQVOmj3qNNeMqs3dZgprLgxxr82IvhLqcX1e1W4g8MK+4breW2JfCqJy
IUzGB1UMz1EKqgABWuTBs/XQ5k73la15CXw/qbz8HKxFo4TEiu5JruEmzAlzUuYG0GHDFdBDBOiM
Kr37DSrB0OplVT2bHbEYTGT2QcNhjbMzBx7Wic+g1fgxWhmyGg7utIVycyWmp26e6PmQeFbI8jY7
LImlVZsw8FcFh8wUT3Tf9KaG9N2q3YYyQ32B3amcvz+hv4gz5aPXCXRqEpiRe+Vg5afL55Rmmzis
3EYHXWU4JZ0hICZf/JQr+tcMY1Q0v9Whk2mO+dSeuvRRvLzx/qvjhErznZC24WHbl2s1O3gC+hYc
wpGCNh/Ivm0Jhk/RIa9NnNh9wXJfm1+FlB37ftOZchVY2qvwyqYQ7M3C2iU1AVRz61ajtHFc2KaS
uR6sDNSOHKTms05BtQ67XHp0i0XL77Np35ytvNPSpipXN4KQebjTIka5l2s5RyqrayNY+iXQ19VF
CEIOA7UTBNvHpEQrvC6GD12E18zpeae/iVYr67aplIO7S2XyhYufqP/pMLhrQXZGfyP85IQHNZXo
ISpzzz71dLLWLox8NbHmJ+HGoN08smX18mlyiSkfZKy1Q0oR9UNRVOe4ZKc9N+vRs+B1O5uY2F6R
0W/CGDmGaqrVYSoSdiXw0bG4k7eN4XLa5gMBzpRhP6Vfkpw9cHJ/1HgE8sdk86QNbZ/Po+xNwY4N
1FCzRr6aoBowLKy6OXM7gPSsaB2W6Zsp/VR8pRVpQ5z35B4CDAtmcMvOOicV2pe3305rlL6FLEdZ
zDXpOLTjIIS7smYj8txwUK7Jiqg3fMgydfbtGVy8/ZuppCXTtNDTgjDzggAQ1k6kouzqGeZgGzoT
hV751UPW6Qo0Im2l0y1JFtU14oalxQW437s4sxoDVTd9KpA8lUkGypPe9IRY0h7EK/8bFU0G9KRV
yvolYHbyWz/n4KxrzW6uIMMYovZkeyk6rHOV/vLgjZ8gZ4+j22CFHsOQGTxggBwXiXQeQ+uBJ0YD
aZ3kfNOzdAzm6F55dEtxkISFWDTlOgKwUZVS00I6vouJhVYhjITb0NF6SMLU/xX2uZCB2RBI16hd
viarLo45enyCDpWnQ2g9Q1FTDMYZnWhmqbanq6VI6lIkRdxr4hvshhgWO4yw6N6ll9jA8Htggszh
z8Wm91k7J3Cay2R8QqJ9youhWTqM0LyBe4YS9TN45H1FJeFkrkWx7e62V3VoZVm9Riwzdfzmy2o4
qc0BAYFioIN1F3fHzOJDZKfp30c6E8YFtHYaCw723ge7of8Mi/u9esjG310SOwwAPHAtQzxiHcih
PI4xeu3AR1FzriBAIoBOIetLvgj+mOlshr2cfTZ0tcPKffHsMUhT622InB8C/2znSCqvVYPxFXtD
GuHLI1S5PbzcpYJVM7V/U9n9ptgAhKvhh1CIz0U+bTn6u9mI6i4SDm9vUOLs/zRa0QvDKUt4M1f3
LgWzCkIRlA8a6HkY3oUu/XCxDhayBH5Dfve3tRyxEd8C21sZOKwFJwqjJ89GJLVb1s3unKN+XQSx
lyjxN8SlDOGna+CpGmaujS6TS9Z/qYHzGoSjXcN0pO2IueNv+Ju3n4RRdjsApsfHmTYA/viCSkJX
r8m3DMJUB89axm17HsBdRTkBDlnQr48SiLSego2V/vJ3uJZ0OHhckrA4kFm/4Do6QVZOViePXjm5
o9RrlUMQFbxsGcjsMfggAXgz0eZ6yy8IJAFz0SOj2HBDHTPudlWMHTAJkPSk3dVJyHgP340b9ohQ
LZUDt4iEXoVhMRdsbnuyaQBbXGf6ovCqjjAtPdLGB8WDic7JTKAaRt+Ps5iWw4TLCDEv8h4f6qRE
yxETUUW28LRU4FUUhpNT6XoRGvgf+nw7ClptWVY03ZQkDofYqDDyNX/iTa7KJUBCgyNaXEr+TtG7
HfSRKC/HqvMYGyaqTdeMJ03T+FX5sZIEpAX1zQpV3rjQw6RmjmXBNFpsYOlqQbbiL+JxLFloiYaW
wIT/IeJVtuXofLTzgjml9eE8gtTind6womdibJaafinsowop5E9vspXJsdXu8Vv9A0rvapCdMxyP
lurAmLtjMSbE/t2yd/Nt+kjycbdF90dKN48ce5dnIPx8yLF2nzO0NnB4mrdJfJSTTe7tyy3ZRVpu
6DPayNknFofVJV8vQzt30+SPqZyG3hX6jQ77ZGa/eQOR5r72rfUmfX0yK5uuYq6ZSEISDl01NRcw
qdPuopOorOOeTzAj8cc4IGxv1VNKjGye85Ri23cGDW7tDoqWA/QdHWXiQdgiGaoHrPnpNPqAsRX7
fAAI+k8BCySpfbgVoqQl/8ig78pxG55kasepbEiOvGVBUKcPeqLeqgfkZHLx/lUa8FHinNPImZxw
ISgJoKUdHIY+bu6/4inTtOGX5Muqx5g3lzR94vJPLvVW/dBXPGkJ83NZZTDdIXURnf3Phb02TmlY
W5wuV1gi5Or4wDLA4Kqi5SbHQUXh7ApkH3BoOvROkHYfXwd97JykUNjDgfpRC4WkGlLA81beCVgW
pXZRdGVjgpYljE0hu7UuQ+apZNxW50iGkrHNqF84AA/xEGICJsb6LlpVxwsSqct4dCE0wkTC7J3i
c/n/8GpvVxfiHs+0frLP5R4D9GLivOMwtRbKPKpqOjGVR7BLEcBtjIRrbILpaC5NfMFxwJT2yZ8p
3EhLZWPbAd15hGpT+GtPbOMj13+FC4YNxWKaffItlj9sRmr/BrqahJQQ7lNP8tmpnDisZDdN2M57
P8MyHiP8p38J13QNcC2w0yy/Nvy8QQHaJf5JqXyFPhonohZllcl0sj7Ld+oZGoz9P/WhAR8DuuW5
WUukD/2O9PEziblboyxnJ2Et7tCS/qKIh6nVX6GHo6GSIpL4VbnxBRDwzPywAlC01LhMZu3WDmsb
zKura/8BUW6XF9frpIWtObV0BQgx5rVNBE0Hhvl3Ewgh7c8Z7BtpJ+VJFxh+BD0m5ytzgrZ1wluE
AZcHAZwL2FNM2qhk+//JPdTx5ahWDZ7Xh/F7k/lFG2vRZyZs9YYPGppqGIQ5poKYPxF51g/2Qc/j
Gq4eU4fDFCu/9J1qydT3tY90ioqtgpUKufuOJmpngdnUO3TdwU2Pv5tZyT9qGAILOQ38MagcKZgI
HVxDcj+UZpu8aP7mg1j9KTmsvrMw1YHcIhERaeGGOOPWKVTLJ3/yX//Ya9k0EPW9GKA04D3yb0xw
hjffy2kjoA6qWaQXkNPP77IK2MMy5N8/tCD7ePIHEEph7FeWO2enl6+byatOKg3Mkkmb2CPuL6VF
jGdnULsLnq8otXZ1H3IPQWPlSIHQEiM3GFQ7AeshCBn90RHuC4pYQn3d6D66sj0Vgo2wW6fwfkuq
XNcxWVAh2p+ZKeb0GRAX/cgP668DQl3FyWKb15LYmISwFY12j9lz4CHCoAWQlhpqzCQp6tQ22gg0
+BsuynHtQxjBoz512ucDz4EjeOd5pFORzMkPuaiTNq3NrH80QcClcVijW297yY8LJfROktBXDsYq
/I+gXHiSrnxk+wNkfgSbL1JiPptqFbKp2l9QscNRvyEMZ7upd+RA8MBt8Qc+zIbKgdNj6GmBdSL0
sm1vJwiZMaY0ZHxY7gkOEFIgDLd/Z5SQjnhHC8P9WStlpzf2AP7nXYYEICXF/ZTcMy3wgfkQ7VpU
oKRF4n6IY3Gm7IjKpQqfPbxOPaPMHM4PbF/ZLTSoZI7mrfb7p7ZChU/d0wML31mWDufHjbtwFjsQ
zcZ5D7emHMxPha5vv5WHqU3tKuTSnbfq6cmUNzHPUpFz4xH+dunDfBgTY5Z6EYVxKdN+uLaCqN6A
c/w+19/K2H0Coa8bLZ/zczzocAzMNLRDovvs6NdX5pt5et4K1bN/U4gHBxcVec6O9bbY57ZilYsP
wZf+XptKRk570RxbVrYDnhxSKRSfs0r5dMLOH0EzQdhGWb3qwJZaAuw4IOGwBE4USK2/oq9YIoYI
gL0b/EpZogAiwddXMb5omR8Qen/npWR227WgKzEI0ZUPq/7u63i2GF64dqREQItloqloRqhpoXR7
9Dt/myE4X0E79hWawbAG6d6VEt/cA3/zQGZl/n1MVO4IXTVex3juiQAbHlkSanXqUHOAljRFv1do
TD0HA6bglPPqtmjrkuI7mKU7/MgnXQeN7aoknMMK0GavxO8NbCyWHulO0tp2GD6n/0L9yPqif3k7
hkCrP1P50Cy1NcfjhJeHcPajwFkFnvWonKlYW1Xqr1V5WagtKzOcpQx/Dj6O8fXCIJ+nZ6nmhTVD
+ZuAIy6qKIq9PdzN4mNZ21HKzlR6wldyLtuW4VRPiCLzrhncWZuVqnacS4GwYZs5Rt6ANa4dKsHM
bbWKj7rw6LTUg/LN0/EUtHg7S+H+HMyVvyuFlBobYv7sNvSjHYlJoZelex/iSKO6pkFPKNVXw4t5
FfkJOBHSIipl0eHmbd1G9WYDBmPO6Uo/2YiR3VMNJAKwrjZcO37MXc8mZxUuyFLrMXz11ZPyU2+Y
m5RSWlN5lbisgggYUtYfjcA6C9J5GIgi69stNIMmTsNl9gB85XyLxcb4XYWw+Y/s7llh3H1iBGGV
87kl3g89lDbdSe+ihCc3UXdf4qNBK0j3uIDEKrD+J6ul7qQdR2ABOlOY78Vd+zsGIH9UND5vJLgE
8+xIV8yuxZV0jM710CG0WtEAuzH3INQkxKSirdH7FCwktfZK2GteYJDIUbiNsWLH+sEOWXkbHEwz
y49OqlvN6jYam3Z1dMLUcJdaPGZPB0eDnIFuu+2Qvre82C6uFk+3ffOssbYvURiUwkzko5t7TeXj
rQATXNvGFWfLGpf9j6CngP7LMm6681PB5y19csYLEqMJDf83gt3RX8wF3eNZgPpD0nLLzMab6n0h
Oly0g/y7n8II5FMkXuhzFjFR6EnRI+oyEob41DFr4aJGpa0UxA6ku6DTfEtmyI6B0yAB4mnHYNMc
EhXemukJ/eLSiqFnYhmkR5qsk4jZUGJrOIBvggQBnhSXmE1uem/PIRlBDWpTlL2o+q/cAzelSKAA
dX5qpZPmJfU/pKgn7wgDiHIBS0srDDZ/Mmm9ohuSiI+k6OrJ/LvLz9uJZlDXknNIMiP7M49wSlX7
KKxhGo5pBaRzkCeFUoa3lnj6w6dZgZgjsmcic0regZFQ7JFRVYH6AIKtKsmNQatzAIEWD9eDdH38
qkh06EF372+JL1/TsvvPFcp47oKr40F4Mdts0Z69LK0Lr3zsHnL5/0/oSjthM5O/+Q2PIOTlHD3o
X+XoUGqV3VCDjtYiCkzdcq2OsL5NouObm/XnKKQcy83bbt0VAkCF6Op+XYqj0q+ld0TpzNOiZ3tT
3BD7YFWDAsTwk1p3cQc0dar4PuVDEXX39yqybNVyT6tzkDXQjCWoew/L+nCpy4NLkAkkQtWHg3tf
PN8HLujT+m1+wuf6ntAOBCGzP7UOsR5fTEDPm/99jd3rc4xFqAmA93aJgbpbYzJARnwuOF4WkWoM
uVi/8iMVdxAfIUOvaH4VuuVUp0ZmsWPiSpFZA3ALubLRbWbARVlhP0sxmrU0ZA/iwJFVQv4q5vRj
A3umekburweyZ2vREGvbv1hpvK4KEJ+EGfLGRVJyDr0cGXV7lULOiLqqeet89AO5F0Afff25mwT0
c/clUcuhdSrU+/ln3Uah/lPbN0FIYWUAKCRUZjjoDOIQmDRNhGEOCSdtZmUOswH/R1GQBjzzLUNA
Hsb757bcz6kHYGdoBZ9Aq2IBslYxIf3WVvPMYgr2ImRM7N3rTTBJIvM0YJCfZk2N8Ea5verKaT3p
TGPoXEWbiAgH2KckHJ9aZzv60St0SWdTXuI4EWcihXXgpX29KvMJgg82X8Xf7zccYt6ePMuQIZ7h
jSpiXl7ZvpM0x8FCNEN1Pg2A6+w6EH4WZc61ZQ3KrcHzPTPF9mjEmx8/7NKv7xqQi4dAbiEyU5K3
MUqhCLfrvYVCn5B8ysLF9id8uCwxOBRDvOfA1iD6ISywPdX9LE4Mnq6/4yQyYUiuL3ScIYuKqMRs
ZuCXtoXpPRl1ipDIvkHJZ9iwtNd4BObOu9SUvk6zSIrtgrzL6RHUnOv339T7SdxWjrV0BFCQdghu
AHfuIuJ00f62xsIi9tuWewt9uCqijmVj7Q6UfAwrtkeW+YRww2eWDbJEPxuobhPt4NSfsYNqEMRj
crKQlmfssh0wlgQ12J/z+APALDoeOyMvJaiP+I4AIyQIyW/Ddxtq57g3ZoKHj8BINilj5KiKyyau
xr/thtUPEQqICGq08jFV1Dl0pe8sctjwoADnNuITL528OD37xZqRA4SaPniIfYbUEjjjMXWPGNif
HuKHV7vr7D21AKRis9I9RDfXyarpDlehUDuc/pQmCH+oc05kqes/4e4c4vta3INekjaeU6cUW/US
X51TXp/usSy+QOWxM5AY+QLJzGOgweyZfaMVn5BR1FcwojtspJMZrrhwdBvEDkSiFoxeVsmG0AfY
BwqsFlStRULlWdR9snV60CU0QMmySngMWGNHbWv++A/IoHDgSXWQSy93kX76t3HULNgSzJ5M0ouR
E3SzuNT5i1sgqrU/4owDVzLc43WyNsOFbeo5dOEg1E4kMOp2HIcl/MtK0REq4uAhQymMfHC1QToJ
9EhosXlMZTmEXlkoc96yRo+SWK3Ju2YGLo/7XiOtZaTDDqDhL2zpNMG/qEQHIWJsHWyoVpxpbS51
wYNyoFFvJlxTqN1nrT3150TWDoHI0hl7jO/+kNIr8+3F6DiWR4TqTGa1H85zhmLR4e54aED6PVLb
nyg6b8if0kDspJs+Rh4cYksqUOOzqA7MBx3HllztTCLBBGRz/sOoh07oBCJbpQs8uqHz/i93mQC7
Eq0SzuVO5YaxdMkoRn04NgpEP7/mDQ2jYnvEWquznjUkwVuFtuLftYRb2hudkXskRTtAhoVd68XG
TYA6J/TetSokv2yFwnr2RD98LRTXAVUN5Yx+CyRnCmj3mIderkpnRArd6yQhe9NehH8HWiKtB1gb
+66miSAVnJZ5dIyfLdDIzIHF+c2H1pAK7HETlLDmLjHb6of9MpK/+c+FyH+Norc51vCNFbdFskq0
1HdTrrCSlnhP7h1w7qlKB/zEcBOiOOlmOh2JRFeD6WvRTjGLoyaqFxzRdeEWblpJtFJwANFUbsrY
GnizZ6wUpKilsMsSwA3qAswReQJPaQ+++syez26zYi/tdOpVFdL0L8zZdxgeMPxIZ0xcKAuFsSwG
1IpvZu+3KjuDmUBAOiw9NYAN5oPdC/yP6LRpvPNqHVPttEY2Iz5unzPGYsYiaHRCsFEJ1Rr4O5D5
0Q6Onez67AJBVG8Fs9J8AH533upLLeejecpxOiS48//lD64E/KGqEedV+jVKA8euVqHCjQZGtRQf
W9X5GCk1JGzorBvUoxO/S5cjtiDSYcB8z64/RUoFT+Kv91nXNurzWZhU8CvrHMjSH/JrTqQWx78g
R41fhpwLyMmMVNrHHyXlpznJwgOmVwBDLhsUbP06atFtFGIFt7YMUnj8A6Zx/HFY9e32o+819xWi
i7INhAwtfRcxsVWiXwZ63DhHUFpZPqg9QQRHpe1l6dPrgbI2s8kTvfzi4fToyWjJ3Ej4oJgAt2c3
+pmK8NmkJd8eKvwrHH67fCbZm0FDpPl3wIcJvZJA/2E0uPOYFsGWV8HWiUZ+gJ8oZXRiia1UMP19
qxH4xoTXZRtCkRv+usN+ybvOcwJD3aZpFWNqnFgAXKBU+JXzVLL2TpdE8yiNEf2DVshDdB9nNdPN
/hF28o2tf2IrtBiVfShsIsOXPPQG4C6XR01vDQLF6VImqp4y44Rg6tkgtBm2UrCgsElB9Pz+kuIY
YuMKvb3/+1S/mdYKoA1N1sUueLAN9MVlLL2BXST+G81XaJ/DHzN2ugHhTRFd2YrcI3+seD1dMVdf
sL4/aCs9ScA/z3zTwEc6B/KAhiPAEsdpoBcUuBmAd0KW8qkPf4JJ12KNKD7Zjni8zOcV5msFIaRx
T8NeVXx9YKXsyfVidV3Ui5rB2zY9Rshxx9wERadzBBixnOHpShX/cXbejx4QCV1RmMn+HESBneLe
OFz6zSscB9ykOaFpcmitB2cpluNfOri6iN008n3GAcqBZnk25JKDZmzRoZORNijJlmDAmr31hlmB
xK0BdZjzlOd1TOOdyW64n9hpqrY9SQ/PKWraXnGwrr/UDErY6AjpsfNSaTubr+ozT/etHUKFrIDZ
kviCfuco8h+WwQkfV7pejsFJbfg+cK0JvA1J6NbspRhbOwnrkzvDe2ah0ceh7/8C8b5Vh3t2+QwZ
UAFNpLt15n4VRkQKJlHLWs7EvjWGmvT0GqKRzI7UjDiLT/26vm4jfubUI1ASozg9PDU9r56+CCZ2
Qqqt/I1LXutKj8KYdz+oTfZKoFsTc+RNECNBnx/jqkILHXY1QMb8Zr8hgiSmmjQtLZzAU8+OwRi0
Zm1GYmnEvz8jVcv+lQKkfU1viVN5A9bn/JcUiTKoRufzfG25GgGDLt7zuwmUhyDi5zsC7ieHaZsn
kOoYsyj5gXrmRYIeSwKMlhUuqLzcLMTq+1NVUPqrzSh6lKae4ukWnLeCTPoh4phFOEnAbo6krBnu
k8G7nyHMQPYvFpdIsLApemgXDDNgGOf7PsFiP4iKek677KuCAaewXZydY94AhtNed0XT5EgTOlTz
55DtcZDdZ2YV95s+Y56ODXF8dHACgVFMiNkAacztZli/2ZWPXrKoQWGVR6zqCho8bB6XuMrcHcIv
9BQwGh+AvjM3vjerSDWXwFPF3Noyu7Cgq9TUdC4cvaTQuhZ0cfeUfbK2jI+BuGRsxYEQ6WBImn52
Vy7KVq9FUl92Ojhb+18mxyhxfDipMQh6q1mws4wLj5JmDBAFUNpHbZF0QuOw6++rMV3fhP/kf5IT
QRER/n5BSnXjkhV8fBSUxBLD0Qe1KEox1w+3yoM5wbNqyq0kE0m9rzOuXjXuTWdJRxul3xCeYpWs
FqoJTUnoF8ydENt66QhIcMFOgRzb6yOX83IvEr+rseqtmslvyIeAy2dSYhtEAIbpuJ+Dbchdnigm
izeb/lFnKBKGehKIw5Lpl43qq3mwJxxO1+c+jT1+lU4grY8c2NwLTWq6RWywo3B57BsJt610tAFi
zTTCax21gcCR2dgjzq2BQD+sOc/0we+lgYC0R+PY9gABTb6GJSRu3PbxX9ZcYiC3vtknYp34P3bi
gZJ8+fCDxO3YhNBX4wk7O7D2qtaMqbaeVgu/XZtd+OyFINGxwrxf0a/wjxYXnqoUaBRJkTuJvyDE
Uh++2h4dlY6izk3JmRL3nzM5HKf5F24h1RhTA5TfV+hQmD9FaZQjp+zAIjIWoICW/D46rBaSOfRe
hQqc3L+6+gOvwmb3Wpi3Vk/NFpJu1bA1XD+sps7TZwMkwTzbO5jU9gI6YEJLedeLvR+U6eX3dDXy
3HPkW64Z4Jc34vJ+VttiMR09qzNVGQd/g/Btxn+rEHDpOAuIeyRstXhGEB2iYQRU7P0ChVask6Zd
InGGJT4tEnZxZfB5I7MKjX/gXyBtjHDs+rNyoGpFH+VpcVBjzBm5bPGS/JtlRvTgjz3qtDAQJeix
9iBjh1AhyZWBa5Mw8L1RRs26UEqDR5kPi71sPnNiGcLBLW6sKrqj8I2wTbkWCD9m0GWlAGDubKMz
A5oVED0FFzlOqWSMGovUQ6DxdtPcBwGvf62umrf/14SzK72Z6KwK15O/CqLQIM2LCKp3pwzGEmbO
H4p3qDx5PQwwyXZdUQ54KjKqSaQ8WNGZLGu7RSJEoSTGDPgiHDUszCmEJUnfDd43WO7d2zB8xzHT
OiGJt/5nvyHloHj9hcpsk8ShkbqGR1jSG3f+QSnqU2m2dQv2p3iBb1eJPTqH87Hn7BXFtXPrGRsT
Z2S2jru/+mdBgzChpbdQSpaZerrNR0NFnWnRgJL3FNdrUA5LvXSGwgHDNtFvqc1jxSSIwYkwy66z
EAEQEL3ikYg+7Rlrf/1uLpvBTF9uowhbSf5GpyE9P6l+kgXhkiop9KlEF/vu3GO2jyRiWAugEbac
3/yi18BTH77aHRDN/50/NoBQNViM77qSqbMkN7vniMLYGrPYbj4LdibS5qhKSjJgn0hjcvls8GRH
adLXGpAri6uMKcWGMuVf4UAIfWJZ62/p9Kivmq598o53G+0dxie1AVecwA9yQepaQgq4gN4jAm2u
UnAMSZ7XZ/mJeY+tvrIalPUkSJlM/NnDbdg86+xPIFi9DP15ESb0ammwNAjsvtcO2RY0yCkQ56An
Tl6FTwLCipBhUVsnmUL8NmMLn+KmxQl6Etp8DHNqIY7u3V3JBttv6jHHGwxoSATNOPztVrH97TNE
XHy2dekySaehas7vgDiR2+V61OGjh1p3QRneIFv6Tmh5+cyq4Vh3mHRmX9h3tMCW+mwscgtlBlCs
H5k3ZW46ft0c0sOJwPIgO8lYI7UMa6lPDv3fw+jT6PGR2Tc2U5ii0Xq6cxa4MbjmTBCyrbxxGCvS
XoncLwivwDm1h01fhWDPRBEqf0C4spBkjXThHDOjbCEl4D5eG2YGSyQZYpcc2QYgwv7uxHH7QO9E
Ukd4yQS31euHg2hxLGf6V5zmr/lkSoQMJgI5nSaITjNOrKtnfJToDT7tzYbQuiiJ1j9XBh7DOHds
t9/wU9PAhoeQK48sTa1BCzb2qveTt8dRIGP3RVOd4YrfWaPGC9/9/v/xT1UskL8AyxIczjDiDPWf
S+LK4NbVXcRz8MnGnnzlO1WYVeYAvF7TEbB6VvwJaxfNkpN+KMh/mbN3JHDeCUsO78zBIKOHKW7i
IMezNLGdXCjXHfkxIVXqS2GymABbzVLT4CgieZP6OKIw2GOMnKtBKwlzCds1BkZseUPRyXhKQ6cx
tQgATRu18MdQvem5LOGr/I7h0UhhF3ab3kvAai6PR2ZRRXqWZIuUfRSa9Wu/C9WCm5/4tJhGtzAx
2HNWH6oXHtrf+WoQDEQDgSzSeZkWHOmK6GncWfD4Y+YSlFaKFhJEswi1JijxxqzIg205Ad7X67ct
TFeyqqsX6/hoVC7wC7inak8O9Vxp237FNnXmm6PPTgJvydJxmVecGektuEW7VCmJT+NuyMcdVlKs
+I+DQy9UImMrp5ruem18QmCK9XkX/LEH+Lf9DTd2tKNAng5YiIE2X0ENmsepGu9kRkf7NFoGYZto
0GBg/bN6Qp70rQfP2tqFdUIUZPelP7qfrpKhQnZzm9riN56n7eE9TDUDTXQ3agFgJOGmYMLT7L3S
xF3Ib5FFpLwHYaSy38EwFUaqWQw36bo/pHCdhNdh7bnf3WxaF/9obXGhZFVRKGgIiB+nR2rYQuyq
0tbNyReiPCakIIBwW96IT0T3atNSTE3TcboQzBFP5f+mKzDxGflGBB2p5ooMm8yGOzotOmttyS1x
wny46EdFkzeNZFFtMsnUFtale0MUi/wG8RzUeju+cPghnYjzv0RRgNFm46coKIIJnxo4zhGycF/Q
Pr6S0LTT7vJ87qr80wCgRiWM5Ns8Q2SCjFKryLo9/dSsnNMaPw5dZ0c62CPzCDMaN6gFl5fyf74d
d1FMMq8yCnyvVUof36ziYl+1hEWGUWprfypqJe5sMckLsOSa6vhbFRdXH+CKaYtQarrTK4KHfX4R
7rbkQzjUZ/XUVTFB6iZEMIZDky9rYYO3GQHF0KgTs5LhI1Ho07vN68F9YABQTgqNvxdeosg1225m
TEK1pGWR6HzBop7TrAjW3tVX66DzSHv17xz/ziNzAMgJlY4mnE82EKOFirpwJTiMnb2d9uF5GK1e
NU95SuXpf02rvu3BcKs4D5nd3+G7X1TcQZ9nhDdcdaP4xvX5Z71Xg8IPFGgVjpdSJO8jrrctroWd
3RctXm+o1J9z0Dfj2KQCdjPMt6efeA6Bv4Q1/nYbyjt6wmzRQpWtBwoIe0q8/WiTCbDudvp0M9nj
qiO45mQAXs4a81TJZAT3VH9yRLj0JLUDFas6mz718DiHWhMXrGotgyNByi4CxjdW+bWkmSHPZbIs
k7vOfO5YSF40LnmJSVY/g9iBv3H9lZnQaSMJfhIFdncfoKhfNy2jZJSHcmXWY1GNK7L6n/2zPW/w
EXfSSK+9GI1BVNBvtu4pDqT3k4P2dlF/3bAuOZghAPZtAzlSxzX1p/+B3dC6yXe4sLZL8HOO69Z4
UgqpkRwCZFnRA8ISnmkH0Zp5MABREgji0L9Od9diBs/Le74MnIbOpffiy3tHio2dShAUNBqHNjzC
ObJ9Lg0QcppeDZeqTGEnpb+cT8agxVjWv9BC4FpHPW0jCvQBWaNGmbM5h1Hh1peXjVTX4IAni4Pp
bh7RRkGLic63yH3IIHK9pATK3wlVICr/sYE14amgNoBAXa1W1mlc2EXZgmIxGEIeySBeZIR3LyOo
ZQN7XQCwY8WOGJnPCMIH+K8Q3pvSoutxYRsL6YsWFOIAn9AilvC76PH5A6KSQa/1l/qTH6ulvt6Z
oLRS1RP1maNVih+CP0ypUckD6bfLsF2FR6XLwOkuhMxOXmK2460mVkyOf8Cq/eYvExgw3FAgaZnO
1YXoqxfmhaHX82CYVE85CM+Fs5Ep6rquxNIE23fVpv5DRDiTzgKOqM6kOj3i6VTlaGVB25hKd0L7
RChQMcmFxg+Irv+moNtHcrvcjHodUlWc9fbPFk5vbYAqQ7EW/9EjR/whpvHDdthVMYNXJO9LW0YK
fxusFsM8ZVRFwaMVQmfVug0TG8UjGhCtJJdOODzIPw/m/NZ24qYXsMx44zMFzmY/kUfTNwTPVT6k
dVfVUh9PTLqiIxtx2KKm+GSp8SUPCyuygpejP7mS8sl01kZNq9DJi7zKa9hBo0sH42kz6qEUwyMO
0XGOaDHhyLfXHbBhC9EJdK3uIv7tzzh+BB94mSMWZWHIHu0Xmn5qwgrYQGlxNFRfpPkCp7IX43sg
eAtTFccIxXcl2sCqahtm2opihPQ2felQd3AiPTRY5eG05B9TfL0+uL7RCXVMNoiCszZItmNQizxv
2o97paAZieFkzik0xDkJZFag+qTkNw9NZmMYKgW6LBS8+PEBwJ9xql9K83vDuCMZXekPtOF4A3bL
Mdm4m0QS30OjinqUU3xKiZT+cqMfy8TJyu9PsDcLWfw9oU/1eqPTYD0+ETENAHpgfBX8LBUV+PHv
0M8uv11VLsY+9wjLUJtaIoEKOLkRz5LksYEPUzfGRgFDVN0K/8oHK3AK7UWIEXfA2ScCa9P3QLFk
baanui5TI4AE7/eV4++6nPJWA1Cyt8J7B13qhhKlUSNkdTXFF+qLouLgOx1yljfqGpYT6NlX6yTk
cR0uB31ln8r6v0i7cViHzmD76cbYTOLkPS92I9n5Mt12ACpMJbm6LuqVp2lil2lHYmnMZLp4GhFv
yGA+6CyNOBwTsuPDJNG8idZpqzvko0/3sKCtQ7E/SnUqjoti6HlUHH0f5RwIoK38l+T3mPcfzQhf
Q1/TGysN72Gw1MqN9ArYX+E+Yga0SvG37CqzGyNvwI3srbq3KjeC+bmaGDopY2BnwVroo4aJFF2O
UfLL+NExRHxyJMPJRr+qTYaUGPfGJa5KNyhnaf0ydg2CTMcGQVBfE320gFRK+dL66Ue76qGc/62w
xUR7FIkdl9V4CdpriIOY0fhQz6J2f3rhbVfPUTnxSfdTHS+U89cGfYNUjdj367nbx9pJU0F3dEf9
1P65BJX8HgipwY+nxz+AI9Ac9rIIzDaIWuKNjfS65JPOGK5eAcxS5UigEp27MYAaq+qiPaUqnmks
0OmTG1/Ysx7TRWAZHhipeS47ipKBJwc8HvAOuDgONuaktF9B/BcjTlOJo+R2py1Mdp6OqHMGS5JF
yUcU2sW1QVOf2A08zZhS+lSoTZDzXT0FHLkRDf1TEj5MNJFcz6fp/fT/btyehzpDPfHfSA2+G9r7
xeHtHj6phYvVpO6J9hYYYHb3ItFALqtioiTfiwrMAO+i4Is4/7XmuuuZpTaZ3uhc9I/o4dKN7dur
bHGLQMoim/f1spKyTKLSPko9IS0zboRS2Y1fWlK7XWHZLa6ia0BHu3jd0QhzBvkcd0VEKRkX+A1O
9KFR+WahsnnMr4YIsTrNmmEMvBUfM/N/f716USHy2ciPNsMb68ki8NZYd0eK2NltJsEbeptyl/5S
nMXiVee3GaMhQemvz/vFSreYGOXo7f4L+6L0RF1ftke9+5y/6ygvZ6kFa5b+fDmrI62J/kHlO8om
6eAyZlFLGFoFNziNy7/ONHeBcYvCZXeN8uWJKAT1mkotIOzMkWxQn5g/bI0+nXlzC0FRtzM2kr86
vx61SwqOpS5kHQ+VwH4tb46v1Ieq+wVpQMvrhqEXTrPIZMljMysMjJIQGShWioGNdPBoPFJ9o+Rv
r6FZSjkWfw8Uy962j8tttGNHTDq4cFMo1/9dMifJEZnXu1yfwKv2GnhStCPhIl00T8Y3tVYi7Qa0
5yr5YaqFj7BPMirLflQKnkUTjGXyok9cbmuIzjqx46TU10nJh8IWqzCCBX1DKQ5nLeIEwr4ajIB1
NO74sHAerZb8UKjusE86hXLtiKfJOhYeMP+iXH4EQIlq25u6uSeglijWGMUxSanPMN8MTPIgK6d4
HfLmi+jJuBIBVSjiTQMCHYIhOH9LbLqC/h+rE8YXhCtW45FUy4JKs0OLM2XYoqW7vYPwe67RrSIh
d/j5iBchNdpT63TCDWHjLYqFm3Ddi3mCGtgJ3vGYMPQ9OPgY8wfmd0pj32IR63u3oAAxkONJoWeH
ZyzNgKS7cgVUDPDcVhEp0jUlyqi5v1Mi0aiF9636ZqDFjWVH0eTzOa3ruUGeLlq5dK3Ep1cgS4g/
2dtkWUSh/x8Q5lvN6AgopIjPDaMz4zOVAQ53wcQae4sejBC8W1i1VZyH0BoYqGj+nRqOHyYxdpBK
Qh2WL5yRBg/2LcjZAknGDNx1cG6OE121/syzqDXw/ZDGHGBCOSAV3I60e7c8D5cAliTHUzC6n7Ne
SOSQ9MMboc0+ofHJi04yqp2YToO7OxoWCCaSGgpoq72avDc2OsTe8NDyFuQxP44B0YZ/vkKyBhbJ
g0ey/uLqTTv+eefk2ht3gcqraVuB/YTX/Sa9G6QOEDxr3f3tdLHzAoILAyF9C5JOLHS/i/jwoMVv
8sSDQW5iioyjSlVB9/AYcFkuW9IFaq8ea+1RgjZ8yFL2auxz7r5L50yHYhJ2mPofGXIVOkSfQTAM
/68mQDTAHdXnnCCTyIDvCV04RGJakzbbk8BYT27GmD2a1MvSX6Hi6dfKUhdnZAf68cyhItJAja6Q
kVpJgM+oi0Ywn04OA26kF9tvNOIY+QvTZsvEewyCRX1b82LmWC22AuHzSKg+HGXT3dm8xj8CY0KP
0ECPIn01MRsscSUDc5sF4hojwVYKqEmFKtGRdPh9vfm2zxdI7pdYm1bJ1flC0GReO9BpUT98fhR4
ruNo9cOSviGmo2xrpm10IEhPPjO05n4yZX25KnD6kTxqIUaYduS0pk6TmolfP2XwfXDXM5Wyb9TN
/97UiMNBRdgKYzN2/bFMXPlXLSFOUgDRIpvRlFf13wSO5NIUyb23ViQKofhHLFDPHb0mNVw0qTKM
FeyJUfES9Z+EHgdzTu/k9nDTPi8Wt4EY/qLRjtx94p/HkNAnyVGdhj4Mvn46NnZXpgHSpTmnM46+
/nKdl8A1ncP1/siQPTf1KMkOTvfTNW9gh9SojMfslYmbREFVhTkRotW/FxxUWOJT4xhdc3fe4qjw
3H0nMxXhCzHs76Pv7F7cqlijFrL0KpF//dXJtEtxI5wHb0l60eGcVanyGja6TONznPpJE11NwvVV
xkxTVhlBjVeBnxZz7Ur+/S0Z+admEz5EOoOD1KLaOFe8BU+PSJ5oDGm70nwsq8TaKP/n5QKYhxWc
GdlacRDtNFs0aZ4I5G0Qe325DIrB9oyVIFeoeNmO6d3GvmLMvcb7MFAIdNAhg3gF3d2NfQcnM54b
wQBDyF6CvWGX6YaDIS4xi7azVyqp4++andlR+oPoaO6ekSKlGr2VXw26tzpmRG6j0BRkdLH9jysu
/nQ/0YxFxShvxkjU9M0fz4QBw/zTysDeEIwz5YXTYdAzbMfumJdJ+YVDzrhSREZocmJ/fRwes6j+
9UpzUw+65apvNx5i1C8VBjwiM1A+O2tiKau70UCKY65AAe34eO0rRcNR+sQz1LXj1SDZjkw4IVEe
XWWgp5DovWU6o5qfhaCMAfwb6sOhlkRcJNUZTTMRjfqa/qSe844t7DdmJTuJB5L1B1cGFhjNPjpM
3eVPcLeX5Fqwy4g+wA+dCqiZ79oothvbf5LOJeI1bdUym6BrJGpfGFpVNqbTUi6Q1k66bCr7jeWo
BZ8Tr39SkdhVx3TBxj6pLguiwNydsDfaKOffD3IWW//eagZYqs0/cQquj29DZZMPpeqOeLqm3B6x
NadpsN2kNS7jrl5+4vSfjLmcdzQRk/7jfDLIIhjcBYky/Jfj5ktGxtYSWkuX1mZVzWn4lRJwaqzW
0vOmFbK4I+8Z9gm7ovnLwTs1HTgNwmbCd9ChidzJ0CbLXeVBqoxuYWsLqlsnLlVsiIkwV67uyi7N
YjQATmIFx5gPek64StzdBxCQzhnjOYJJGbTIYUcwPBotjwrqUr1Jrzil3dWptCmgHBix3kR1ltUr
0yX1sEsO4NC1TwWI5cfbfuRF2nnqGxbd2QRbdMrmwkFEXJKEO/Nl9WYawKGk/X6x5ddkPSlkSKyk
fY1/9T0An7kjmQKFQdxffQbOS0ulcNxpTLHS6AjAkUaBvSDTWGatEofVtrPVXDBjnbRHHNQNMKR3
rMUoHbXkmvRNXqTNKsyowLVCkblGSnKmMW7aeAdwuKfVvKhCWfXH0BykjhtDw5cmG3WmiJmmG3fg
6F0XBqgT3uyiAAnuibbAYYqpFmdXmGc6C1tJL539fTmThqdt7z/I0OQDq/xoVUywddr5A1drskFj
cmEOgoHLDXaAl1/Z+xLKqnB3WuZVsRo2KqDUePdzqqKuc9DfuIZ8chqOlX38dBiuz1LG/hKv1LWC
YSbMXoetHFjYdLjvbYuMKP56sC3B7mDIKE84aObHVv3BGcCpPobWKT1FZo9gHLjcqe1+n8j2MQq4
ekCNb4t4sAulr5hpvfzmuK2GdF4iburpTub0/V5AxTGojmdDPNVFY+K5o/c2+D2G12LoqH8lZpB0
Vei5668jvZ6M77fShEusJAI8KjYqhmhN6Tc/2ye7iw/MCRkTCkbt/nKMn30cvIN0RaseG0Iq1kLr
2amArOv36Qddns3/LTQaSLpu2iaTBbmr/pXIbmL6E6fYUmn6xNNDM8gpNq05yf2MtJUK732PPeak
bBDJ9R023PLpPBERig3cbBxxOgLU3WFHPzlexNeopQ5EwR6Fca8NXpAqRl5MSRY6hzdhgQ3OQciO
h+NgWyOk4mAdokb3FoxtTzx9KFsAP6iU+ieT44cJqk2r3UjxJB88fQagrmrAm9Bj9NSRjT/UWX/r
/r7xXHGsbyQ79tRmlySI1XXqTRNX90XjYd9WvH4K5Ff3PLJKhIw95/3T1eWMI/APYq95N5tLI0xu
WWLVISad6cF/RrLQ9vBdihLJ0GTzyJAvyr7SiGAWgopmJ+SrR3uA7jSMaRo395fJGCLyqPpXtqG/
4EpdBmwNZUHHmLrBdFmv7QJNx81Mw1Pg3Ct1W1whRnV0U1xQrLDUyxNQf9W4p2uXZlGYVC3SHAxS
qZlrv9pZfq6dyDyLZX2ocO0SXI96e8DlnsTK1Fo28xiepM33XWI55POXeB3pDI2ijSjUVidKU+0s
oNGptP3FLuSRx8rZyAi9kaP5mGvWMIHr65uY6B7/IJgcdhZ1ou+gHJHdujSzS3vc1oyAD6uImZus
LMSrR97Vh/q+bc/hs09p3MR6BK5aNLB5MoO49zwg0BaMPngD4N85aClnbJYi6D8rcGWhQX4oSPKO
enKc3y1cLF4Kj4Q7kMn2jXBh6+Hun4EaJewcnbMgw3tJpImtzIh3hTEcRnKvnYF3D6rOmd/cbb3s
5Hihuuwwg+OrFJUb1ivAdIXZPLTijQKk3QeKlHlqvPZlAO3Jka2Qe7IDcn+LJqDYTos4JbEPQKli
kFKUj0sE9gmwYWNEtX3CB4sMp4LsKbwTSDyu5v4VJG68IWMHdNuq6S9u7g6WtdCXq5w5z0GLCPgI
1cfCzE4OWkbLdigS4SAHWO2Dqyq1/aj3L5KfoMxu1DI4K5g5UKBOMYu68n3bG8cC7uR4AHY0IeZg
lH9KFa+0he8B67VcOIA2AQtXPGWPbU6jYAaVZr+NBfgulqdGLiT1hz+qxx5WlI86wUn9mRYSkV/6
TqJ3h/UtQgUhxiPr8kqD7BpkyCBTKpXk5P+ErlVYlz5+UTZZ/JEmrFlfcCUeBh2aS79lVxigghpo
Wyg8aHml7aWWcCSpQq3pzXEoR/dSVpEOJRQPSYk98kLlqqC1Qs5qgnzgj2jqKOlgbZ94boo/5OhY
9+FCJLF35gAq69KvmPb91xYQ4ddAjRpRG6whtJeJepdpLS08aVTlAr6ga9YnDk/m/SdclkOdmiJ2
Q/yqKEjJsfQeYgYx+N0RWeTWf5QsgV4g+NrW8IRbxEy0f8CoJCAMk7kcn1dEn0kHnqBNKqCR3dWv
J/d9VvwgdlLjW+SGQyJuBScakfXwVaM4f9M9LVb1tf1WCIji80nA01GcoHt6bBUdy+iWTE8eJQeH
XlxDZY9HVABaFRvjiMBKfO9vXZ4qXXv+BoKXzw2SpLSikuRXUTQgsxCxG1CNpomVNI9dO1K29bzq
REHzT16luZszMX5Oyo104w6uYUA8pD1tvunAwAgawGaCx6xyq5Bns0If4b4Mkejf/uawza7ZVar6
F4a9cP6aaFJBbuyc1KZDeGpSK70CQsHrtsYJWhv0FYMHR5gqGmNjgJKLLQOsuNrP5LSFkhrhf+Mn
9N8uSQb/pg46RLmwqFDeWk1VpOzwXjqhh4pBcfkyvOPTFdcbcULp1fCjPDcxle7EDHBINSC33I3A
AgC+YixtKauPre4aKhxH+q2XBT43fFqNq9oM/DFbYDJmqDeD9DDVsLTd1oZNFBHP9+/WbfqWwkQ8
BvnNwdLv5yB/i0nXyvfq4i5wS6eejZrReeyA1ZXQU+Wx2xHGSYrxKM5xAQt/N6yg+cmTkYqdmazb
jK3PcfMHQ/N7E9wKHpa48tC+ueq+9/xw/Kdn3XQnenuh2QuGLKCabLTNQ9tgor6Jl2KY6Ie+JTTy
EiBb4uTsksGAzDNAiLVCx4fhjcuBSz/i6QMAyS3U9ttetUr3NmhOmpYBWhBJVQxzNm4lU56eDdfs
hijojLr1ODOs8ivcvMwSy+CXLkTZnM9yBiKshXNgtJZotZuw33ysEFPAOcSeZJ28eagnljT5CLvF
zYnHHnkae5zywo8c/Lc/WZoumrW6dERP2lTXhdQa9N8ngmWz3Z3pKxRbeUDQy1oYjjpu0eET2j2C
ETOwb/OWlxI/GE1MzX6jrWT27qdA6KyxFhMvKqJbkaGvGz1WPfHO1a4ixS4IXJ7ahkU4azUrRi47
esvNBqRZGburZ51bVd1YtytrlSc55zEnnpmTLbpBBDiYoaaIJkKsOZBeY/VjKsM2nW1CFPIlL6g8
JEcBQH51Xp4PISL4pXcl262nnM7LfBSww8ZNJXxPxc8Z/8vHOSeJwkf31Ug+7AaXjxRA2nyCeQko
AoY2ofxwI0K5v+r/dlfhHdBoHB8tWX00w+2dnh+J11B+LomEp3SUtyPLWYmfnlXd5ddy6jOWYW36
DYRfR8wrVl1sZRcBw7CeaWSryw8ugCBf3cO5Z9J/KxXKqUQLk7FOeph3eKn4fcimcH2+4fhTWAjl
dRaVI+HujjKWjqqdWKaXOLJ0AWdbgPC6CUG3HLj1iK3SXpeXFWQ5G3GFFBblxzlzfnMh58DD0YPc
9O2MO3ttHIqgiYertl5l60yT3UV8+xXLbaZN13YmDyoyBjKa/kBMcvjm8rweA/hynhmhnkBh8h2N
Vko8XLbKCUqgXS5hRhcebO5v6vb8nf0KXF71O206Zy22Bfrjx4V3VSP3/O3CYmuXVDq+sg/e4S2x
SHJLk4x4VDtxED2dCUKGsu3MXLLQWiKB/MvKdSklmnWKC0otRjfXkIbIPBLM/VKEbpWLlvLIarkk
cls4wRBru+PhCm3gzmnlheCi1ZU9296vTWKfavHqZtFUxmgWuC42lJnDdl66WwC9uylziANbjHDq
9b08vMHUaMSzE1kquqJ4AlLifcXwjR9/f5VNtMijQmzPZ6HttZPlSYLShDcEAfhsspK5vrN776JA
Y9kZTS3ZsgLJbqMxMSotvDgkTRLeI1pMwBQ7YhPJL/8A6QF3cFcxgBCueuf+CD1iqkio3pYFyEMm
5dKYttnhDrDVGUM6NYr8/MECynuvH0uW9dF2HyEIdds2JIa0WBBh4rRWTiVlgZOCM3/wGWrhk17V
sVv7XGnDEixu2OOXnMHtVkJoaoT6I/kpj9r3cTajwtWiIvw6cS9z9heZlUdRgp5P2bIGnzsTGtiF
HWtfFOWYseUmrb3G1Gu0Nul7sNk7gFOPYcN5j/om8tPKe1VDovGTW9hvg/AModYLMLEfVJVuBhkO
htXCCI7T9MfulRBCLm+wtxdQv5bp2lFsxYFa/Nms81IuLT2BvrZ9o8lfC175R5dFrw0ReI43CL9X
aY5unTNmuh2I9TWCSYdQ8r27A8qaKsUpePB+++Oyhu09Sfd/akVoIiZFVMNfxRGC2vy6kGSYFzKu
qSoJc9ScMDUPjOy+gPOYl2GnoNtrUAB91Lh9UZaCQZIsw9ol5WyOEtJV2hb/LyjWdlqhQPnBmJS0
DMlZmkixd3jwtL8DHZgP07i5Ze58pahA+JuAxLgekGjjcI9b8ltafo3Us+037a8GZGyMdxqQWpqw
6LVT8v8HhLAD53HUIM6qLGVW77m9EB7aKZSAEfFo7hS0PpMHAKPk2ETvbCYpqGFoWOeLmiaUJQCo
FtNEJZTrvIW6ZVWci6CoMsZdW1GPBtnUoFNKR3RgR2CjhA8LLNiwqAsE/nCe5m/B5Bc9Ozx4Z8vL
qEXiCDZFyn00eoy5flDGGn2KlCguKg4f8UKPjbmpfiOswA4HERWFJTt0Z+8FCTGgcXVpp5NtBNOs
yOIgAy98CcD2rNiji4650fSCfEIirjZn7gpywUEt7ZKizJBdNzh7wtkNuHh3mGlvM6ISAnZqqmE2
4xzl3ppxR35xIzeo+dUOvfEguWBloMU+Yw9jjboTdNjPeNJgGcUVZ88Rzwc0meqmbbsgl9gx4B+X
nhml1iAmueDRfKkU3VR+0kv66aPCV1bQupPWLtjuDDJvPZeswkhU/qiAgBwBLi5b6ubtpa7S7dJS
ago1GbAaxrHgcVSxXNonqSZaTwDJEEmkHmzX4++gP2fy+DF9K2/1j4wuaYcJEeX+rakRzYkCoI6S
coHsNX8q4CJ9LpEAtBawgMeJ5e19/IWTcLGY+tUJze4Mb+AJKQAZx8aF23mFY6UQT48GXwQVe2xb
cNsRfCIGhDH2C0o8gjcY9MQh7KPkUpMHmPGoN7qOceJPxmOciI5OCsyEZhqAIVcZH5GBPXLLoL4H
XQLUWK027Q8NOT7qmq99dOcblH6rv2lYmQ5eZRboMI09q14XOJI1Wd+MDIE3m/bKXkpPtQqZCdOR
/5npQHGar7mq240zNrsWb1Dq8/J2jlrwbuzFCFEs42LnMrXP2EC+LnKPCg6lZqeES/nTqSWEG74D
rbJNlG4CgK4D/4rLrrq4fqkgxzWFW5Nus+MDLUt1j5FV93dE6jSczuGzbCaCwvmQp5H2sxEqb+1l
N9PcTWdyhXz5FPT10U40QH61vgcx1xAIaTbYCH4JtYaQ6yAWdyNh7PQlHc81YD9jknINxBn0WW7a
mm6SaDmmDOZVcBpa6ak2bKkiML+8fSIDb6FPLfNQO7fEOGQQzoximQWbaT33bQnJessepC47IIZf
IeQs7KHlyLHPUesDhHnXDDdS3Ay/lbxdhgWu90FMLuBFQsHI0f6umclY4mBfm+huK29SxTONO1ws
IL8FoDG6YKN/eHTZHSactLKLrwwdBt38J5ddXDqvuaIfz8Dm8fAcbHp7pjvDds0ky6YXczMxTyLN
vajHMpr5ogf82rTxgMnnEvYAQEzJyXyW8SuasNsyveOEHYoiGupw1Zzf7dnEYK8M1zgY9tlXotlN
Ge/pf8oxOnPqswWES72U7Pp1kSWgFADArLrWhYSql0Z6G7sMKLo/1w24AM7XaNDipnOq0UYrVO97
i3BNnG2aOE+n/UNgnJ+alA8skG5eIuMLlGb4f2Yi47E06TnnJa1I2i1zn961SA2RoUMEliz2ufGY
q5ORhyz1VAtYe54ctIOVc1yGp0OZX0M8ts81M1IrFMVHsKQlxQlIEfi4K+SwqaRKoAzJWyqSw0ov
Is8ER0jCxXEys+1GJY623xM8zRqdMPXdau/tobPzpkWWjFhniYmywMqH2i+CizDtA9HC5Y3ObYFt
1Igao0ysl9j+A3ESVwDhhC1LziM3Xp6ETosLSxyLrpDizIMQaRuUhOvIfMMe4+ajugjHOBskWsd4
lsTJohfaTK7JGofEq/GtiERLTKv9m9m4mdWg24UEuVI6xhG6ODiTYMi5V/4SIL7cMZLtPAXU6x0G
mgtgJT9zaImGHbSC/wMz68yz210ERuXeegsNMZc+R1Zf+S7EuSoFGGOpsfmpwi88oYXiV2MPtFzI
+SW9TdSYcZauLmETg+IgX+K+ZeC13XXe09BxQ8Bwk2pkt9gJkMsfvsSUJ7uFwXW2zOWkkBNqmDkD
HaPFE0/fSCLpIfjANx2RPH8qWfwgktwo6Nw4vm7s6CE7d7Jw2m7g9JBwm2DA5gqWA9pwA6ofzLMt
Kx4VS03O9cKfI+x1xRXWu+qpJVZLPw1s3joMeBv92VaESpykBt9M/5saCPWq3wcZ3KO3+BQ+aQif
nxp8YGGz7VzzstZroEBRV6wlFHdbbY24RLnOw66rLeqTUvJZUpRbO7+KEMVLGA12e5/iTf7+n09B
9+3Tpe0G8g+/zwVwFl1gHZpALDAV4wa2iiXeInR82rY/xE6+SKSVJrkNrZxRHKOBt5F6w3azOL34
FCfc+2SraJIoBH1ullmU9crIF+46qcQhTkrbrjymEe5cMp5dRX4rnDMJsuIpd4mEIkE5w/gvqJfn
ugQQFXTQDSMJwipVvDhY6o4VwLEIDv+hMZTAecmn86agZO+Ly3oW8yYa57ZWPiGw3hIvdUAhG91o
yXbVPRhNfDTa19ae4TmCubA2PJepc5O56Wzn8IyP9xzq8YV5JXB2CgxwPMGBi6h69vG8hWOipDzu
sOCM45RO0+q1aO3LG4z7CtTcxue6jiQE9hUH2M3r28gJl12H4NqYVkZ8S2CLC5STV04NL19tRzvN
VPg36DByrFhj/TsBGf3Rn9ZRYBKcsA2i/wNylM4DH3JZc94qJJ5/AvIUTn+xWuGWu14jy2t7rXOy
FE69RDwcVuhhNfHC1oQMg1D9+QY/pFqU+tFHxC/bCd1tku1ZX+VGfGB2LLy3wzpUfvhvTkYXdGA6
tYPYlhH89ec4VLzFZIbM6vQCCF9Xc2aNsd9ZZR4q0ngskWwPsnMFyaENl0WNENqCLaNLGWCR9wg/
ElljaBSKsEK7SOjYM0Uu248/dOCDkB0oUmESBmkMiD/UHoAL8UD0oq1l9N3rKoSK+PEzOeQRJk/r
8S6c/gcfWV2XhtYVuVfgIeU3/XrxY7kECaiZtxo3X4ytpUfWFb8Z1siQZPxGiFFPeUCai3CgLBfl
zwoayxR13hXM9IufKMOlnwdaq0p7WfEZk+1MRywBKbTbmNDDWlJQZaSKYsBcVnlZnOQ0YSyv2cKS
dsntX2zTUnk4nuSEQ1B0jpK6uGCo2fpiGZ2TiMbwjqs+4QtcigHNuMTK/2ccTY4asROE4GPPoY8W
rFU9BvNinMOhdqlyY86K0HQHD22NG43xqCZJCYc+b9Ix/tIeCyxoEkIKoOw4zLXD+QdqCNbnJivo
DFczWa5f/Re02Op48M+4w1ojV2qz7UnJie0Ubc9Q86wtwWYAhQRk23bzlnCQNgK7kpeGtStL3Nfq
SOlV43dvEDw4+YLP0qVXYSInS2UP+GqpnkX7TqZgip44KBc6b4vWex3U9JoMcKpMKyUnuz5ECtNB
V3kObCcoZjgDfvBW7w90v/UJBbWQ3+ddbSNS/bMVdpZQi0DeBrMccLYX4iTzQXuDmT8yx8iiHT3X
h0HfVcrkXgbnDM28bD9DmmoA2qtGqRFD7sJ9VzcGa82QQhpuYk2HJykODXlHCVxOnXvaXglWoJSz
wZwdu+SoJL5alUrRYe6ggC7/lTglVrUXTmWLd+1nCJqmD2uAdKkTzfSmsj5Aap4RD3RWe7fUrqix
EWnHgfPvtaMszJx+SQn5LstVVffRm/5dJZXh5C/zDPQGLdzvVc+veybzrUh6qxe8PIhv912yHqjc
M9OaSESgQZyAw49ZEcOvzxM5WRj5ir6xGSKBt1cSCzAV3BiKZaHpTMdo9lXoiUmffo5EDd2WDJQJ
nbKyIiIoPfgSuonU+s/nmrL75PbR0NE5MfHe7duE/6V6zeHO2VDQs7ZrwvGVI9AKGBJAk/bksvBl
sqafTVKdV3GUy2bRLM4fHvATHsVKfQmA1Elf2nR/1m0beS2WjHXW8gHlFKekYK3twzohr+S3b+2e
ZJPh12yxkOJ7cWl2q0QIUDJgzqkmCslcpDxRCQFO6zBHrDGOyTx0Q7fz0HgdQHEWfAUoM0LyoHFj
SNyCeJ+ZA5RXrOq8U2LMgP+iiAxoPyBbtdrhHZhhfn1VfQQTVacT3yOx8pUGFAc2x7dsEJHrTf22
XjjN/IsSTymkhPeY0Lr5Qhv+FR1MfDv3bEiQyRdmvlrD6ZM6sAmZ4QP3Z8HkOo2Jw+iuhJntX2xA
wsGQQdB2FRt+82uSTaW9Lfrm5pqx+VItBE6eDYXyKgUiBBdYZTMDxQ0FTflyKmFE4+kcDiPkhwju
inGFcuvk04Pl4FAv9VYkY8QfWpFDB9Tcy6PKrnopyBKLlOsUMzovf+VEHw6cBfVFNtFYSLWf4xSM
E1a78uDZMbSaV7jWAAftc9vsevr0+I4VuGNR9fm99GMuSYyVFDm/86vAzQWYBtXRTv39hBuJCnFM
afzLmLb7s7ygpD5S4ur4bHr6D9pVlC+ZekxXWUcBLAjlVPXDK5ZrRTYgdltXJZ5c04vCg8ooPotE
qBVkSGYRL/AIUh9wdcRmjJFnSeFv/aMgBGkdn+nrbNKEdjy9ugNhG7FzB7RtOMsvbiMgNd5GvXAc
BR1zdelUTNAlui6jrT2qwejriSty7D1IeIYuamwJoam/jNBoloNYD+rV9jHo2FiUPjC0ZulOelin
nTkp+G7lr+OGhmoHK7FH6eUF+GVLbQS2Z1FfAhdmG8a1X+oOYAXGcpsIdT5Y/SEnXkK9ejkGLUq8
wo90vj1qnhKkWqiLakW/Td7G7lRtsGrypK+1elcBx6KqAdaETa3umeM+WFJkR8l7++YNbreLJy1X
0wBxRUPYCyCNzKee30uCd082Ztvx/IRTVScCPK6rdexqzB0O2bP+J7b/Xhupl3jA7Onz1z4DsbWq
hF81ASuAD3MtHI4ilxh7NWUf4rs7pfahc2+phHpHAYC8DJmTAnkoJQRl/+sxU+WVvoBi3vOY9t6Y
pOsBknYXmYx6GQSxODiUw4xZgA/h8bMLxPNfvyaxjnUwse+oOga3YTFN1b8980VUsS34pTlWSSHc
wL/isNtYdb2whVJ6HnPZwWFOLrtsH8EolvUSTOap851UXtpDxDF4MNywrIH9tj7Q1WZFmIL9W/v2
uw+9GG0uFsrn4Tb/vPxJ9Z+tVess/+u0NikVuaAQq+1WvfakG26kR1wrefoSRxo6jAwJ3vWGSi5N
XZawQ/pCGdB9lZ176EEZBcBxgvvPhR01+VCmfTRaw9020fyLY/g6+09jNiIjR7vSiFRFNMPeiUlj
cMPJFOQe7/myn4RV/wGqd9gWV+9P7XybrlqoxeHWvWq+5w0rKDX0vy5l8LFRhLCiNLSItAzeqNoE
+MWM8pCnM4CpGvWQU+u/gyQsVOeX83QgR/zFI9GBz5ynI45aA3wJO6kjyuZdXWn5f+YhzLVg0a9/
Y+KiQjyj0M6cmqBnBSoJwBVpOe/JtWN9ENGwc+kZbVDO+kC3ANnJ62Zt8NsQZ/a4eEMMc8lXl+5/
q0T9rYf8XQdXYxvWgy/CxD49GwlnN2LYcYRDeb20OICrrEe1aSS5zsK88DWOYTncsl4yt78Ws23w
nUfOkIR06ZJ7UT/5jxUviKva6PmK8ZvbH/XqzWPhz8/QNQqbwPFlX/2ZnvrVu9R04FzC6lacOsWS
di6d3y2UhwibyFdoYILspYRlh4vINs0hb4GzNHclfap3OB1MF/M9B7957nGZupG6mUVXZl/o7zKu
T9pjFk9zMwLSD8lDeBQsOhTc9nXyhFpTMFDZFg+oAE5dGQh+uij5UXRVijuM8mix70BtRUhVaLTs
grghZHbzV94sAvib39aFHP4xcRVvHss444q4BgM4XUcrNzMIJ19jufltBBLx0++ACZcOJ4bNBDr2
MHKH3QhOuL7172uc4F3Diys2RdTY12JCrAsPJ/9Zgz5d6RPlxPlgGdxUXxO4YmPysuPKDuwlrpjQ
KH/YMOzle1Y+Mc3IZp59a/jIB36TVMIwIVCVd0vSaKtVgAkjitEeuB9PeRzit8KoDC5S0ws0cxTM
uD8ufVkc5zIZ+YipdGTPDiAfB6HdUcFaK+YFvw2zjY83b508egQh85ShWxZk2vBBSp50hjB0RDU9
8cp66dusaoVqdnGNqxMRdD6agsPpalnN5sBDUTZBye9pVC63f8hWDIS+F4vD2fbLtZ4vpHHT7Dfu
iARqZD4wRSvR33ToJsOtIcEQtXpoxakneVznIyEY/ZbFgIpmPupCB5vGBTJFp2vVIYJyfK40SBp7
ZVtnUncgLmHeDhz/CHsVaXHcpb2VSiCgCkXRdigUysLH3ZNcT7t+qtci6vHWDFfZUwnr3GHPv+MK
rz4odBu9Z8cU7x/huPd40k0/ydKmpF5aS2R284ySHoynQRs1n4VJQGuxd2gUr64EozV3UGzFn4sz
bgLprnAYILOX6CPBV1PZ5Wss/zW8+cyersqKfgU6mluh5L/B9vfylw6cworzeajROqvbzabCRqu8
+KO94PqL/IF5i2L3e7ltsjIDrLULr7jsp/qu96FcemADp5ZWRQh2OtuCZixKcVujdNn6pb/KXFp6
buFdQ4E+PF1VmjSZizJnftszGIgHs5kZVy8oYsNdntv0ocFRlOECdkIfzx9H3ANSIbLZiiHe2y/Z
GkUmMHrXfMjKn5NRpPc6O+pAm9qrxsCsBWRWOgCLCkah6GiS
`protect end_protected
