`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YNZOfwFmq+EKwX1iXTqpnCzO6NCkg8iVZ15wmEqF2fK31FdwL7p+998IAHTcmvJXXulOlBvS6vH1
+iYCkUubZg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSuLWicvAgz15dAyaBM1McguU+c1OlTxM3rwIjZed+XVwT0aj3kC8vBXZpS89nkrz4cH1M3IFZBK
zd+c70XrF2f50b7PhHzi1/zvy7zfnrDsI3RQtNlcdzxESKaNa2OVRlTl1FiVvvM0flfMEoGOVBEg
CInpOdHF1+GNpH3Jzc4=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c0YpjGsmE6XFKBplkrecWMiGPy4/BXTRGoswHI3n2HH7rRfRrIKKFBskl5r4MXDh+36ObQ/r4PAk
tfwFXdRBQQdjX794wIxcy6RXY7xcRmOpxCWwo0hF7M+Du5JZuTdvu5waK1k3RHlAIf9fMqtpFqa4
/KglkgOK46YLWOg98V4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cUsDUT+TuVyMSf/EEh3e3oVg55uMy42ju7dn2qfNxoV/6aNQsmopR/owNzHJ8w2iRIbnD/sWUeVD
YfC5Nh9wQkO+W++ModGSDC7LnmRkQos1o2QXsyGO7CwRp+BAnJvattDBYemVwv4BYerghJyYxugG
VuaHyMph06OOJqTM01KRiHL1l6599aYPL6x1/zhvgxuLp5p+bcz4yWnxtE0ZoamT2LCdP7gM6f6C
edWtC0tvUpoBL6a3+CkNW424HNzG7euC5cgFf3whD5KjxK0sgU3DOgHfGxtZT3pY69/36mu756TX
JZSijhFRV50xlcUra7R9ar0hdrBRjEOSw7W3vg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
msL2o+GmDoFk+NL6vgip8zUMztiw6jKP1JrnEkE+4rDO8UAEw73Bp+XaWDJ56xzku7n2eZey3ZXo
5t0kzk9ueKFNecgIlJ+KU5U2yQqYWSItsRIQuSu4rKPl8Rqn+dE0pcawYSBPhVOsFFtaXlpfXI5E
/6dCGckETNQ7yeYg58KrKQfp5W9zaaEw+sE6ym7QBzCBb3dmWjdUqH7paIeYhjytGjAkhoofSzNg
g8k2NBO+eeLdDWD+xxiRjuDbJXen+TTEMwG3QFWPP6FJTr097RR19HGV0ON+WT7z7zJCaS6N+Ajv
3OxS7NRyD6qW0oN/CBWf8OZtJ5pG6dKBLcxCJQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kXQIZv8mrCnXdeUXTei22vQEDigOjr4M+bzu4+tut8y+H4BU8tqpgWzAawYjBx0Q9HqqEYYKSACf
UeawwsHxb2466iL/YrIN9+RqC9NKqlbJC0Gk251C/dmXlDQUuvsewDbLU4g9y+zb3nua3y4dKwNC
QE25LX/Sa3SyQazOgoFWwhfEsmEbi2LDvoNJWIuq7sSOK2Awu1VlnbJcXjjblq6y0akDL9wLxa0z
9pb1oK/XSraNLnR9asMy7i1xZ7fwmuxwLowdIK1CU6T/qtrhXctBLMsJlQ3gnD7FJ2klrTuK3ilX
2lNAz+VBfdEokkhLi1QPBxGu0q6x58LkOoJ5Fw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
BR1Q16Lyg5zz6kUNIT1/rUVWp1M1MAxsi8GRvHObVeRDDhUtG4HwVLWBhwN7oZq1PeZ8fiBCeUnY
GLuxSH6VPc7Ep4Q2rDBs7DAz8dfWQb1LnMEB4lXwtXR4DJwittOqTklXJ0bv8Wt7aEyWWhCNKKio
v3x8RzWi4xSeOJTcl7VvmVRF4ZCSbzSi3gwZ5D7NkqnN78x7qvs9IaZ7+sUk9tqvRGcTKJb8mFeh
383QXS2Odp82BtHJontYNTFemShoOdmQUtt3TCT3z8DS6apGPx2XCsSyUzLnhCPQB3RG5LJgLaKP
OSpTiGNIs2Y3voZU7+8ATsTkko+1szYoG32QramG3zNz5HnHxcasFU56LZvQ8G40S1vZWwZaqbpq
8FBRHEi/CRkCJq+z1w4DxVQv/FvnFyfVVglAS7WHs7TgafDag4ZAgpiyOlP1hBy8c95JR4kv3SAX
8ASRqInPYY8HLN6A4mImkIX3YQge6uPjx3Gu6yzUIpcL3Dr+qgq+kNiKu7UQnXZ86IMYeiZz9Uw3
gEpnq00YIaccHMXqAvjBrljJuBAy+QEKZ0tmpaJhzBUNRwpW8pRZXpzPb8SssWvQHQF6UpTw1Ncn
cGF+TveIZkx6u8CbTof5tY+pGoxAwbKXVHpQGy8JI/YApoM4gFB3kO0yGeMVsEZ6pMWHyLr+uWJY
hJ8LQYicN6CtmGkdKgHYp0WH0W9QuE2bz2A7lCwsTey9NpPVppgw13WRweaZoOO2bmrhmQWM9Ste
Pz14BsSz5StRO6emnbc6g/bg8wdkdEUhAdg3Q9gAtUTtKtAgdOTaq6S1h5z7163v1gYg8jJnuO5t
i+v8FpXHhjWKetJLwjJu3wgfhG2zeWQ1zr6+2nEoZFSBlEpocREGBPBbqTENGBxOmiXeuVQj+j4F
hbS+n41nPbaFEmm4MxwCOWF8igwSUN/QjN9RA6wqjcY1G88cFeF7SLMqFlNsxA/c0WnJlC2jCcIg
ZkkIvUPBeBe0thAxkSB1NNfFBTgW15BCD2inpCFzX4HWWiohnhEyKmMlXI2DhNvCr/da0JkOPpXV
ZK4qG1nHxY9afOsdsr80zjOklpilxqv1yA3GqC1jjsoN2G+7DFX3MqT3WLtZgO0c+TAfh2/YjkHM
z4dIoFMrYz6JqFxWCDU80e37UuuU/V56w4SSzUlFxsxVc8sj7JnVC0D/2lhu5i/csncT/1QkLvsA
gQailKvcsWcH4cZJTvwNlohWvjVVX69oAcJTWtA1Qsn10vQ6FaOXar7rHmSYrLDJwVikZQHM2JsH
o8zcngFSO71GAzB9lRx4jbVjOVYo/t1aAuHH9XQwiuba6il3yIkWmxvPy7VPc7WuDA4fIl2eG1gi
pSPrK/2o+scJ9NR627nnUkBLSc0GcZBgHSbbtf6kLV29YdIe79rruwgANFjTRsaQJxmTbh6aDwTQ
ZgiOSUj7Yh27d1GhU1TEhmP/HLBjnCXWkmjt3lIULjR6ktBzulf5nK4uONilkUrrM84BUGhj8Ctg
JpYEu0pQ9fhtHvZdagKs/4f59HU4FwCDsgBf7yOBSMG08gfNK38kT4uWzO0sSGjO6z0cgtf4UzgD
gJdAncHFQU0XDg4+Uh58ldqUQNs+xj+Gb2OoaRKW5ThG2u1VPGGuFOud/11QuHb3xnhkzxImMims
JGdrAQ8/zlZghI+mQGI7fugi5U6o2hgiR52YSPou491jSs69Hr4o9+31Uk/O2+qLgB0iQmroafVA
HvURSCmLQ5OVjH3GMi1VJ8/dY0i4kNxTnGpYwr36q1VjxeCN1JJuCtw+jH14xC9dd7jY9NsIBATU
dwyw2D8vSx+m55g1+FMlj2WirC2fToU/EXBnCCy3xvbCX2T9mIAwti69ziGNJanstLKrNns3dfwE
IVjvXIkrI1fmrovyFJQUV8zFtnHZjK7OLB/dL984VmPVLS14K+yPbVUR7HF8452myt8FGuqVhOma
D1tGpzWIc2qwTVa4CFgAQWbmMoVAt2bULpy88F9NQ1B+6OAUd0g/4SQZmrhfL58W8ddIOZSMd/nA
zaHh+zUH/+N7+lwGQ4lF7cHnp1Jc+tEbssDNxGqVPsYrCXb6M9Vyxqh0GOZtoJr4l00CLF5fn2Ho
6G86be4szTVe4TZheAT55nK431wWiuDCR8SjHJxkPpPxKtEki14IsUrRhnnQdk+ubjbnS4Vnjo2x
JwlMSHr/W6IFPk88iQDjUYXQKDhZpyfvQqKIVhGDTzOuB43or6wt/Yay2Ux+VfGU6907WqjZu/ft
+LH63N7k2ySUbOlK5OLz8k4mcRRTDDXaCDs1lc2h/Bv5LQ3Rmr9iF1TXBeEGwcV80HtDxjP4vD4w
JIwiZc3ypYouya8NtbvXbbfEdVh/Vzrx4CVGHybD5YXCvQHABHcgRdP2wxRSTlc1favJyU58gsxf
lZDwsfuuV/mc+SZuYxo+kZQNcd7J9AxSRO21OVPVdlNnVk2b3e7NsVF9yMhVALs6co2FWrca9rYr
QawDNpQD3RhrhzSDsuOglPMxsX4IF4GLNfENamVh3pHmXbD+3aR0Rz6ziB8GOP2A/EWbuBfBX9jh
AS5KigAYwf4UIvSm6+U3s6wCeSpP6O4dci0rL3jo4bKllVNcPuO4/tweZKafgFdyn48e8XM9f6zq
abEfoNT7izTjBdJfzh5oiahi2U0Yy5LWL+tvdkEjSMgE9iQ7A30yHXo8MfSb3haME8n4wfZP3WH4
w1BcU7EWYn4hozbJ7omyOudp1GyROpgMVVZtu4HfXuKxGblAIg1irSg7Vk8x2xm16H08bRDJZp9Z
v7UDskSoLjQ+0I+VjEHdumlOpUA07/Yw1x7NBJ43pA6M1w5hJjpawm2AJJYPGemTfWW6DhNy0Yh5
CO5E+SwQymR9rDhe+MjDXrfNxESS7eQXm4rUkLOP6BzHTmgQ3ULwlx7ChIblxiTtu/j5JndaJoho
YS3ugUPcZSA/XygT/BP6faJkR4UkGzweUH3OO2tSWp53KMC8sqKhYfMiArPqMK3eDozMEyoeJ2so
C4DiAjJG4mZzRBAPzl2RtgWDEE9gmZNHKa3NltxA73dHrad9qdKB0OMtOmLX2HfYIpu24JqX7FGa
h0+NWZlBRPuTGV5WdZUg6M724pJHnG/9PDhseTqjG/LfXITjD0pE1Pv4G6PyDJ1D5YrDrsgdrtBE
RACjmYj8jHAbj9QiMFM4U1a77UkcLLacxkIxiv32FLOoYQI5LYfkrZprtuLbekpq5HUVRua0D65r
SBRRnxHR0s4Evm32yhGnoGGhGMqHzl/OmBs90jbLwXQa+yR6Jku47XStOziHBtfOteQ2EWlswhdo
Tft1JOCce9uxEwjAOJTOlaQg7sayhSE8KkF2qllY3lPwez+bCMkWvC9KFX4UXq4ToWvh/gIwVuSP
LkywPwXZoLN3hZjmhrSUQmsrNp/JBoGW44jCtuuvyczAnkqguIFjVdEhfRkty8QFHlTFz7GqkeEE
1HrV6ffDOJOYdRndqdHVNdp9SOqGWmJ+dfT5BURCdTxdgjqw4iRIhBdl9c+O5eA8+H2goPsL9LUK
6tx4uOx+g6Pr4/01+Bp5aCrsiiqqDpTGi4/Y9mR1YZn7n+njtA9gm+BAbDO6EzSmPe/fa9Cn+cZF
ndzAjkZ0GOWi6Nv4QXM3FffCCAWUYKejbzS769+rXZZc91akEUpG92iPuEykeg4KAy3pZZh6Afmo
z/ja7wBXeuLFxNZ7LHfkNAqq/PL9DfVYuotgjxQ/UCXTluPo9u4hVyfN85EmjeiVIchysrlh4V3u
d8FDTTeRaODMPl/Us0F899qnepstx8W4ZdpONVMxlOf9hP1+anC1iN2h5gauKgqQ8YAh/L+xLJ/K
3MUh8jRw9EHg88NeL2wIex80Mx76AwGb2S62cSO3f0yYUkvAJsC3NydRwpf4qgGvMtgfxVKmwYl4
RkLPmCWhAnoLuhqveWvvEirP5txkHZd/tYJ3VRCS+1hl+Lb/IRXNEOEdH55W9jtAdN5JqITmjk6O
cxpT3R0ez6GY+q32Q+kPul9ER1gBzPPMWWdPBxZ7CJsDJMJLRCK3f9bJPCHe/y3cI/gWF0fY4iM3
QGgheDrSUeVKrTSCjHiGE5qJ6vcA/ddJMQnDeuF/24AOK6iNHHIkxrCuVy5hkKvG6Y4sryVOLEUV
alshUJM4J296SJjxNSVpd4q9u2jTvwQY1mXbp3umx2105H7FO7ThU/Lf/rNpdGOy0yWFUvQ13lIM
C9bCmhkkpFvo2h9F1YvJmvHRDK3NZkq5xgYxb8WH+1vryrbA+Aliop5YaAAIXTxQwJt2lfJJXcfZ
dg66dTBJ95Kq+2Tp1z7vhggalibPOttGx5XYAwCpYXZXmdMnNLUSTCOXDWQQWvubRgfD+MuspBqV
2eu2FAgn/cYid4mIoubRztD2SXVIVfeZYAgIJIVcHbb+AZeBRsM/DfmhFUdYm8uro/43s2ez1Sgo
+Tn77TR4umfbvll/IwKyfUoME0HDLt1S+zmis+8rkOGun8nBqMSgybe9vSm4nXad2M1oZWyUoaOx
7KPbT5Tt0RXXtivmmKbchL8FmSr8niyjjMG6CSyEQL46lY3Y5KfUI6TwGLAL47EyiL1CbNxfnKa+
B7XbCdYnLY8PuZjNP3ntyEhDr9mJr91uK7HzfKrEFrI/Do6H4rDHlWUDKC95gLcw3bqAV56/0bZP
UT2NY8IRAZGwi11YmDzanMy56oAh0WIcJAkNGhzwR4ozuIIdxVoJUXMiL38hK15jsEo8nf4jeCnq
WkltNuQmtGJP0xbWtSiBCKRBu0ezci/ky3LKU0EjH+TbfHfEObfYiLjz5ElVb24XOEHLbCk8BrRj
8CqPuFOIcWe9ex3VhVrOWKYPCuqVwxwhiwZKhvUNMUs2pwa5XQB+OK5Yxwly/OMX/G3zJ4qgz024
gTmOrJ+Y9ft6HTFBhrc5DCEstIxR7IbJlVGgzwaaW2LWZ0YLhFOQ1gMQFqKS86tu+gISs1LgdPP4
QAIWY26C9rDbWuZeBNI6KdhbmL8c+yAnQ1ir2qPeiz0JP3KZZlKfTECbgM24FsfdEIr1pt7Rx9Qt
3rTY8qmkAwcNEUxK4BDAEWw23aNimVxXO4yPkXJ8Dc+q0ietgW9mXaFJTmJvHSl24sOVmwIzcjUQ
MwbyjdFIObPlwr4G6oAsbwDjN8rvhq/UOU2rPvyGkuk0otim4do5ul2aXX80gok+vLMiA3XZyob0
izSnDBk5ooYfqlaPDPFRqdFfNU0eGzb/t4HvCl89qT4FKsRynkgxAjbja0JPUlJJP6Eqm2sH8aU2
0BOYSTbCABhunP6NNdJ17SEbCwVVN709q53ZplfzU6yllCARZRm3jBLbUD/llpf4a30wAUmYI3xu
XV3OfrRJZSMSUIGn0mDnILPtm1vCGKhH4RHXskwhrU0EgB11kkjXJ37ecmoUQGrMQcNV0pflIxtp
w4STGBZXkv70WzmKYYExXcTPk3gGl9DQytj9KCAzEF0N5gxYp2ir5xX6d2UZFIxtZSZcITsSYC3X
2lOeEiNDos6nP7/+yJXBgI2zsHZ3jSX6VIgSCxkW7QtUFpZ/VMm6kZJYzerC4Hnbn6T4RKaoQDVz
OfQMsqW+asrudukxZyEC6/gaG4uFNNnXkV7VseuNqdOiwA0iluvBsFFgR/01tkTvYaAnxCHYG8vW
sSMQKzPQNrvqasDXpoM0abfGqR9GvvVFMsXuLw1PhArVu2x9oWXun4bmI1XrE8lbbK4CbWce8HsS
/j4XE1OhmU53iPAx1e/8pXTvjv58aJ72SNEEfoWH88qQFvij56nlmlHiip9aHa2S7bqss2d+2qrg
4DcxLoR9LKCoMD1hO8OOrh5kUnAkEj9p0K+FLGTRJR5dq1Xw6s4eCBrWgEi0KI1ZMm++K6sJ8c09
Hj1byKlobPmK1sAcsfq8503siyNJpuDWKVvuAr9whRVZHmYIH0EQSO8N0bp717j9/g/8I3OnDl5j
vsJwl8u47w04HivS56Veunvx/zcR68IjyKcVGYXcwG3pObmVfe3KphK+YmG0k4Ddjbp7xnu23wH6
b/bLqE1+5+DfzDXTsMIAg87Yt2dDx0+y+5/pi9cZHLlNsxIbcaorzv1PpsLGZyd1qY2gGM/d79rd
LIwsvbVZaiWeaIa9evyy7jALJvJvbe7UU645i/lquN3Ilk7dE/RDGcJerMdIl3J58p2g6X7MxCXW
4W91NZNcn2BcWkOMAGIJkigeaLdWQxy1v9phJiORHqbdIoeLQn1avPCJRCnWTnWDVC6hE9dT/Ury
JGJMLDADdMQBeJIc8eKG2SM2K92fzdf3AuF78MDM3M1J7SDtVU9J/7qN5Rzdg4rS64rhT+EnGByn
uHAUKs/RrJJx+TtTvLiSNid0zMNMKH05qriw0EdMEw83hm6wkeNEooEi5ltcziCMsLTXgVmAj2pc
Bid76IQYvZZg+GfVyuZCfpVrcmislWROpw3fKv4FIlyq49ZY3zdyUvtnCMZkNcNekmvy0R7I2quR
Kh45SfO7PcOGrubW4H9Vnt95GtCLiVvelbNsh0Bumk6op8caUIHyedpcFM8VVE2HxYpx3NIhqBdh
czVivuiMfKTaSzODkrOyY90DAA5EqKF165SThok/x6K7yPVOuZnu0LxEIlx9arnzNN7cSLwx460e
DiRbDg1y65vPJ2WJ+N0OG+o097XNEfFcJUIUQhOqaPFMQhU7ynav9TYRbjlSu/EuGnCIqvBZn4oM
4VwFtb0xlVSXLIrcSqKOgGWlhGum/OID3NsCWVSRIgn92x9Kl60ar+2j7Uqt/kMMK/Pyufmkz+6P
UQ2le0WoYXUrF9ORuuJaPklkt6iA7w0niMGUDw7S3EYjE6uOrcanqez+KlbxFxb75o97uFesk+Pb
b/0V4O7S5WAuJ4qVQd3300ZYN0EULUMc7uzvcDTkk+Gw2EaWoYSJHanMWhHklnDeQ4t5SrIQUwwb
O3Qmx1XoOTwGghv2ytqJdiZI5z113urzEe/srCkZ3fsatvrnFYtpvQFFxkIPp5oP16C3sNn3ADbC
ur3kqqVEzwwuS5KM1qQKNKsOh+wiF5efUSGb6wKxhhkihGdV3pzZniEWucq/o2dAF6rL7UeB4e82
TTjMWOtRM2oGA2+KGV/mpAAcZt290vstpOy2RBHsVJDp59Bf2tnHIuy5Ls6xjAi7urOVolMW11Ee
Uel2oDZzh6DQBC81Lsl43LFFHLdDjPcs695d8qRgWbonBfNpvVBDUdPdGBrGm3lSRw6FsIH4A1DQ
Ejpms6oNu1PFQtmnpzBtEGdsrIfFbNfBYEeysNl5/q/Xu44H7+hxLFwwVKr8EpVFRdtnF23lvn2Q
rHwnY17jlXivPgIN/p+woSEHgre+iTgC3h0ndrn2j20kgSGdD37jJJJ0H6c8OqaJEWvFKhAN8enT
cyvM7c+DqjY8GtaECTPEr1NJ7gqvKVc8u+vXGgHZ1oAsP0UdTFu3aDeD03oqVxC+wFqdvG3yqCZK
bvoUNNYE5c86giQjQUK+JKXR+8EbziMeQPE0VdCxuW1KNtECcSR0rEzGFIFT01lvBjy4VX305CDf
ediwWyRxsCmix8XY/dlBw/+h9Al03W9j0bHCgYZHSVt2SRrTLufj1s7LOJ66pt5u0v+fk1N3vZK2
Qotq4LBIQ0ku5Htl3QMnDz3XUs2jijaAQ1M6L465ssh4gTdeJKbQDw/c5ByMgi+70xDwLoGY/X00
uDGsPygdyUUNz88waf5cPGEepMsJLEDcpj6YHe2DsYdlFWycZG89UWkbo05tXz6qVmZZS10MN66e
FejGWBBmymaZOAtCKnMUKNCTT/z56pDIG3vsRQMQLn0KbyO2EOyvy08GWu9gvRyT8SyCNrVozvjR
xPJe5FhgrJyq0utal5efWvLR3QKxTY08V6ht56rLgANt7lipYph1UG9rmj/DRghRCTXeYpP/V1EN
o3fOEUUQ7UbhDjwJ44RVWYPaAUjhm4EoiginyoIBmejWCTPOIaRQHb/wBx5rwkEKHtCTaojAn0JZ
TiXOmZL80zhhPzroti+QMveCnqoH04b9TpmMsJOYgN9+5b0OQb/G5FROgOjhTxD0LK4lh2I2LUGy
eTQWGCvkN010fYgI6IbPybY7K5NL3fNBXQ45WxJ26tkQBxRQHj+1CeOvk53vKYbhT66mCKsszJO6
RW2RE56pGRNyIjZjXqf+IMw6G77eRalpb2hUdCQR7t4HYbbER4dgSZfzKpY+SFNaqpaG0L2ha5t+
Q5blpq887kdWGy3dRetuvQCvcFnlZ7pkrxWt8+Q/GbBaBxX3t4O62bFc/eqyWu480q2ImQrDiLy1
Opt7t1hJQd91KHTE7ffxwB6DF75xAp37OZKz7ixS0lAGtOCcvV+EkthiaohMUhEClI2XaUt8Hzh9
pxoy5FyNajYfN6n6iMaQs74Y5rqpmBHAU4jovBoci9jlNGSiZUm3gPEQmAGCvAfbGXB651m46TS1
iiGCDrqwouZmI4S1jDva8Ie592zfDxWf+ArGULOeEM2DJN+r/3nkgIqfBNXLwUl9QfQMyN5dsli1
NoQ4cZ6butVnpxZzfRybrUE1mSaMZyEekOK3fGbsMq05mjfRMEZC3A10eaBdqhGQ26WywsWgRSwQ
Xb0yuCveCNh0stJZwyZnFXTL4qGfFdjCcrwE2XDUD0tMORbLKwyX1WycEDw4AUbLKAL32pqX9gSJ
pZvGKhwjcHTjpN95xYpEC+TVW44V3P1XbNc2ofI77ewBhtb8hmEIHbxF0pHp2c3cCvgog79SYUPx
3KqZ+GmpM/x3jRvQvyW3E+0jIyNYOFTA5S3Tf6tVM/fCMMYU5AeyuB3fi4HOl85XVPp4+tZc+BnW
vEyV0GuhLBOgySvGNOa1Cz0gKw47ISsJYysuPzW5ruDYidh0zeToG6+iQXXN/HrBMbqzmIuAAV42
BgaPudbEg5SXPHpAPaGxfSULJMlSu+6mklELSTEh2mbetT6IE6nL3v2ipVMZ7OoflRLY2CX7IRpI
u4ucOEppIDYNbGjbPit9BJlh0mSN0ONclQvNZ8pGFP35m4Q/95B5yMFSKjrZrhy6U92RajzXAFCo
aSTGbehpMVwRxQFs6I8RplcpwPOQGfUccd8vqa+9MS46DfWD9pQIWfoyIcIZPCFsWpUgoe5iumyJ
EsdBFGaKmhyF4+S8umgUae+SWZa1NOrALEyg6eo+pVjo2q0/T6wPNCWNu/yQ93vXvKuUYtXyAlNt
tQbXbPcCQVFUi+/aFFpPKXfaso9lcJrpJcsmb+OwL68Jx/x5am61Gu5f6jneS8ZkKVU2XSpg4svK
MWSMzmFr1Cf80ByP/yRB+68Kh76zInmqgEuroh4PUhbUG2rUqFu4/XcjODWfKe0a8vXaK8RMP/1b
cABZeqpjaQxEv3lZ3vW/lwjW7HBcLMZ+kbTKRyD1DHQ4K4mRfZiyrY9vQg5k7A1LTHELWij8rcl3
ti0ly7F2lVxJ5Gz57Ab8WjXT+jKw4ARichRj3uiIGZhVdY88TTfQHJ3MdLfOOBcyaA5jtXkxUrTO
6eED548WTN06oK2ijnkJeVy9A1vjrETB2DFdVY3svHV1S7e3z1yX1Y1woOvM8Ki/fqQMfhTBFV9M
A6l72IMYBEvn638kzyU7PxG5dqFypWtuO0hLTXMQcBJBZBTZzi+LjUtsOSE0dcqWAM4m3OxMFNek
tpNdczeLp66j8GnPxQ+TTYXGiaLgbSKiXoXzrj+Omg2CylIYeNoMBJrC8vVELBjf56l+SIfATDIu
lfOZYktfRRRHt7vPWrGjoROzh2+BOurZW0eoXyeryqT+0ZvXsI6uEyqVYElm5URg+2zfPh5Fq19T
efd/xfIl6nKLEtCgDlzZe3/dQajmCCrr4moMTIvxsiNf5EYpPEclw5XWwPxxlZEWlWdmkWgQ99Tk
1ho4KFPoYNRvbTTibS5avBmy17dx287+MGFzCzRv3DQZ7rTsvIWDchECwikCQzJoOQyMuJ3R0zAR
9GGspEw9LIEoWj/JgodLPbFosEQTWVi1F/x9P+DgFFVrBKtA3CNxhdv4JQstFtZXvl8q/TrVoSh9
XGl7wO9jlKLlnlfpU+9wi5WhdVH4vm4/2dPgt4pNStp6E2VX2CaYl0H2fN6oemDnd8pJ8reRcGQ2
pOfpY66VANypT9SwD2Noqt8M00XJEdnC6fsFQr2THr90SovPaN3USHB58a5o8tFrrDBc/vukCVQi
Q9BaBEc3qtJ/165NG8DcTMo1dFS+QL4LWgQnR5hgZngI1DB1OUqFvIOD7oTJZN2MalwR3pfD5cZS
WHVX0fn8m/zWt+3ZxrPpeHySd+NUlSoins1W9npHgfOPN47JUGjoguf1t0CYmZsWg0xLbFgF38a2
dEJVWP6HJKaoP+7cQa1bXlrPCvqrORZUl7gNhaakOEnbaQft9dviaKbCXsUTuUFJ94+Hj5sCz/2f
tAoF5O6F2YWUC/MCZEPqJeXfN/GGrpBwjAhiuN8a+uIsJ2bdyd0+BezcPB1VAZu0ydkM4SVxt9K8
hteRBmwGiZuYfba+lZ6jXv2GftfJB3NnC0oRw2/yUjRLozuPeTl8Kq+PguNorq2dttQqK4o6BANB
u6gCzHptqiex5iIINKjG/emYNszSeK6y2PbQ+uS4wDBRy5JIABsIiZXG2l5jy/CZA3jKUHnI+EB2
go2sF46w2B7820BLpmaNUSt4e4SfO0W5lZjICuy1HjZOWeUvg3IWESvV4E0erd7gXsM65jbpIDfb
Di66ZzaXKaULR45IwARDLF41WT8C4FK+zVhClH/jam32idL5dxFDeqMMLrJj5Ue8ol+UYeRerH8C
y3hOzyJsaxXb+Ojtk62SN3fqT6XTpM4O7WUMkhWbg2YJ+wHaF/i5Y6kgFe9VteBSDwhqFY40QKzZ
ojHRssGWIcKCbErhHV2b+mBEesS6b0ZlPq6+Ufw4AzdJuSqaFq0jZ9uZKqW9neBsrNl+dkeuDSLY
QBRzQW/wH2+pzqrR7yaxAzPhZifCJ1RGxYzptPc1MjuMYwvWyYZwPoWBFCyj4ib53eVNpVwMqEV9
hF46W7XVJ9S0yseIR6MWy/nqMh7lKh2DzJjubOksTZwUzqoI5MIdy7xgnFfZnNKFkTlO8I+LeGLq
/jsgorocKI/eaov/kH+p4ntxzZ2eM41lz+N1QYJKm//9E/1yDNS1HYLQA0z/qfuAjQVirAuz9iFY
iDeQivkBtvCIIL/7ldw7oe9lkOLnR5c6/3Ggl+QOxUQhqSqmyoizhlgbR01UJ4/rd8lhAIdNaYX6
2j5HjYgOpipKXpNXNpi6W9G5cfmiFZxDCnfeYCeUXaVOHrIwHmleu3W2s2Jspjdp/Q8235xlaDLS
337LfEB45lHJJUJ7K4j1IgI0gm+WC8rAZpyW3Rahx7nFtdvFKvlvq6/FdMmIGDUvNwTz5R0YId4s
wjuznAOX12wmI8WCXw3garUvcqrw0R+/9JF9qboMeSCq8uLLuHnbkJ8luo9lbrt1q4VebTpjVQLG
uswwTq8H99BlrUOMHMCp9UIoIIutSzKCeleC4xGT/ETiik0cU9CcdiTzzOr+XRsRI3Y7u30ex+VI
13DMpNY5pjqgYejMTGu7I+Fuw5PwnE25c0YCeAG8aoBhZn4e3Va0omVuXU6m4ZApuTTvQor7tov3
gaO+afdxAStccTq/tE4BQr8dc7NS/rQlxnSImjoi1DZP/u3Zs8lj/4MlcqqMVKsrHhMACKCulB46
ZBSm97bVlvrjKNksWETEWJCWFn+8sNZru6JnwGHleZ8hEJyEAv3tD/YJ+7bwozZczuNu3NELNw3s
LAAI/AE3xroPjH4LQN5P3rNmzw5lpiXe8l8wvKkKR0V8KvuRFNF5XkAMhH0Bb7qQG5a3yAZWsgw1
i0wpcaKzB414famGkPjln7BW1kY76iVZw353waeulfHtb4WztHYOOLg7760vtlQovtCMjwjRAkNC
ZOuMG+wywM79FUuj4ReVVKt7+m5pGMoi+WI9y8bzhwxVWbgc/loPe/Yvjt+oronMcI00tXJTyDU2
R7Ov4VakyfpYRV3PY11paB+SAS/NDLZTQYes0/YTq3ZZOEn/dqp0blwhLxFp7fHSFzSNMxdfUPEM
IIDeo9W+JyBH1rdrAwVbKjv+Odx9TdlYSj7sAuWsM4xi+eZ2M8jbfb2nYrSTxdCDz7FEq6GhgJXn
KCnAweiBPct+i8HLZiOUiYrm5zg6AF5Dtt+xRKJu4dywIxT2bLZCryxJ73Onp9ps0jmrdb7ashpM
h0XROh6oj+Xh2tDZjQ7UI4RGqq5+vqEoke2ldswDEQN3cT2neGB+wnBkBXWQz0TFQoIhqTGgfuiZ
CZcpaMkGEhmhrqThGsGuV3rHtVdHrF+lPfe0uPUCCag6vlrFP4doB3cuykeqX5OrcwrwImcF20Wh
zLMIO9WsfIUDCI3DUXnF74fGl8ZH2jOBAl1cuPlpFqjd41dhQ8cP4ocpXK0Q44xu6uIPaMvk20yC
L5C4x0D8YXF8ccFVEeD2Hk40HD8yBljjdj56lX4MV/5Dmpp6E39OhOBiBiDHwR2f/orM2pOp3mTw
ny97EnuNlEDlraUJnSzGZb9l3ny3b+7Ip0aYLrz0wp5aNqVmLxythHDztQVKs4hQY9tncW8Ngp3Y
pdz+I8m1zt4YANLqt9ssiovGfOmzGYR18a/VBTzAfjrD3V+mQyRRYNzs52cIqVzY7twTYr5A97Fq
5TyD/4SiJ7V/TQoztW6D4lNxjp3pbKM/UZyLZXWOu9UAVHi2F7yRTFl7zBmxfJkUeIJ/kVfDxAR5
Mnx8kWqVGv+Fa5md8zEOdAmjYJioNq0wjFqRmbgZxXbuLKwEtqRZThkZqblglD8LjAeRH5HW1ISN
FY/WPenQIfK0ABpH+Pjtp2MsWKyQMrD9uYpjB7s3TBU1s0bOR7eBaP1Wh3R7Ks3NBQayXMoYRcZG
/LN11EMPKhIoKw+4xVHp49S/TsKGe6ENnbOIodklKMW72XqsJe3H8lihpnKFj3WOKkKWklRXAide
I5NHqwNbw5SFg50mhmHf4HdmJ12lLycmEVUneAw0zB39kXODgDUyhrqAsCtUUKUAWIZVlnnHze40
h1tDWQwYIYiEvhDi+Dl/MXqqK+4OVZTojBBW/Nlbp7lWU2ERiH1812YY+XC4wrUlpEbBQEHLb4ir
HiqWsSBOx4OlsQPJ/arBaR6LkNHsp3LjNbkPyAjFEjuGjIvDBzHTJsSQZON4sZf6qwH4Yo97O+3w
5PLLOhbKmyTmwmwofUmnYYQfShUofVkqZ3p/HaLDcB6zlPZ8+dq0jBdTQeOHOfoA+L5+4cltfdYn
lzh8qmLhaK9NChE7JC7oT0o/uCkM0+0baDl5YaN3hrh4e9puX3A7OJsOID0JILtIjBzqVStwjIzB
+rs2qRVPRYrx/74OGfBRAH4hODkDzXrFk1bjd2RizcQEGkjc2+Ahww9R0tI0BxBMaeMnCbSkWJqO
jwG8Rj4kGkeWnBbMlQUPsh+DNaYAK8bHgM/cU03ebESCMbI3pExG69Rum7kw8BgVXO4eCYeZvmoE
CQPoxfWynx/s/v+kZ+Z81UzlKRYFRgouM6Prus+IY52y1eUlDYcVZ76TEGWPVFvPZ65ggiuMv235
kBtv7b2ULT5ipo+jGdj7zeLMN5In3drVfejlLyiz1jE753uWpfrGWf2aGpcfxgOIYhuwrd9aBz7I
AJlpthPKUFh4adlPRPvfrS0UZauQlWE2/9zH4TfbaO4MaAPPM0qDRwbnlK648Fd8COVmjjEsFvqv
2odIbgkqQgJUybr9vXa8SmWQbE+VPAjDdqrpzN+C/ajN85Cynxo4FxJVsOmG2qteFuG8KU0plB74
0sHJFpCBMm6h3XttFDCU+z1Ehm5cfiWEI+lZQduafxcOiYvidh1lcmoZEd08FoRsQ6/z8G7rKkYS
sU5dvHiyo26iS7oPjbtmLJQ9RkLuutvCSl2cW3U0Dja9nRBFnCxB6VjmnLs1vwxOp88I+IgXqcM6
Lg1RmpYf8YQe5WkT2Yz5CZAr7We0eIu7dP8RbJIpNjF1LRlHcxwAA17Rr8309XjWbHI8bjJavEro
TrqVAJNBk/mqJQhp76ZDJsruF0LhenCB/ryuNV7jd2lscNldk8f8cscYfT6muEnFn/dn1/fWru01
sKm2YIshX97C9Sucan1iDlAWbYx/7VFI3MeBZFKs8geSxCh2I0uBxaR6lkQk87GBzOF7CBcHChRm
4p8r4iuZfdpYNLzb49wTcx8g8D8P4ejI0+qPe1byIN8yTLnfNHe+n5fhNUUFo4YbNQPV7epZi0eg
mdo4n3xonZhNLyg4XFHnRRMxUa/CPu+wqw4TLXkkNqu63MoZu4AjyqGlpvvFNSL3BuD241TnedT5
XCxBhkuy2yHQgBno2JGQXliDhUZB4mkJbYf8qyRl9Y65IqgOnWUrvKWiQSEBaBztwrC4D4T5uDB9
1tSdbdiCP3ghr3REsmohLXbf8aTwPxcqAltP4+09zSBv49qmccwxeLNrgnyO0IfYTr3Yc0VVsp93
2agbHLDW+h5HIv58tHEUzRBVWXLYDyCfUzY+8WDpMBnWO0ddOMhWBuw8OcxfgtvR2rfpuqIALcIL
IGc+IOxczLbpVYo/NYlxyZB+uCHSXKdLI1djJh4R7HrLC44z7UtDZsVlabok0bUzIm9lfNPW78mE
22nOkhotTmlugk/4BN0nLNjv2JqSeagKPJUKeJd3G59D40OQw43k0x+HRYOCGD+eSr0Lp2mhcup2
e93to1buNpWkZskuLZNnOX1tOe2L69k4snN77yZAFdd55PNggrkpp+A/ltHDc6oDiCmc46DbaNjj
nnYRmu4WzerhLgvpFpByYP6uXiEVIauntwb3hhMcaJKf2t1VzQLOf2ThGXhzZuspJ89Ytb4gHsGk
zhGhKAd7dnyNz1cWlCD0M9PwXWJAsGs1ryLDJsP4GvGY1BOvBMRGwTADTEXo5Nw924xG7QieYiyl
87qUUiPAizlK/kqLFA8/CyHIllXLlgjybNI5aIaDKw4+OilEA0kfT6rvJNNthDE2ooTTJdFkKXPV
xozbJFBSaS41v0eRIqs8HfaX/hz+2NE0iN1aR2PKmuIOXsRPDmhEorMs0QZNFVYxw2sKqJVVeya2
S8+YWZ5/4m7B9OPlJUZZ9+w9GvpfQMmBlnslL6rhGqadgxl5GOzIH8xfqhmOUc8vbMTTAnrbko9N
NcIvIzmwv8GXHXv8Yk4sNou0qLBM/S0DJN2LtNueZgjtzDGx3PSkPkORIy/fdtHySF1WIaFEbxWM
GeaQl08L6OCggFEFaAB8O9Hz+ESJxq5IG6LKM729dH3ycwG/SsW2m8euBghWHyTDtc94eaubFxc4
B5pT6Q/puOmvKfnmB+CRXoVOgfQonp/zSaw4aoNvbK/Pnd2GdgBzjl3gK5NBzS0dTiPVLB0aXQvH
ppTlTBTKipY0AB2s2Vy/Hkm1gne6yNKVzy0HcB4Hsj7hCQHI7pXeFQtqE4bJ9TK9KldnJ3/6Ezer
MGlfiKLyhvoqbYUJjqipyZUj25WLXo9uS2Hb7DUgK3Tec7z1tyvaiOZJVZ3ckFey+xxxKYLLXVD3
osimiQafaIdpxTcnMG7Q8pAnM7WcRCgS7Ha9O4sOyPAA5XLDrO9mxZAfjLrRMt+WpmzxlVYkSUtb
bKHUZgiGNuNEpBsbVVVQ3GWmK5hVkvzKpcfY79ZHKdAj57VKyEAyocIFoSBOGu3DXRkjKs1k96EA
S6MlfzZq2kstnUKN5J8tMXtsEXmldmk6y/79ir2M+TiZRPV+cCapva6DQhp1lx/F5ZDkq5j0rpYW
LxPwCvDZ2lbX5mwVxWr4J0p6E6waq2DQOury5z8nTR1oR4g33TNuGsaGDXdw3LmBkwpEKHmtULP/
Il4557HRkFG+1vlgfF3NDJkhVNmpKnAoPqziWahQ/NwTQu8GeOTmFE0ZU3MBe77KcK9AUey6cmDX
5iR+5uwi+cIkhXY9gG8gVu5f/c8AqTRuYJem7623NsIrj0Biu+rQuMPxES8kw3+xxf2oK0+5Sg7e
lh2Q2oHbSBySsyKl9vmPTPnp1L4QDRO/PnZwoeB6aj4Y2Fas9SQyP50vIYJXGqdsG1jvIjUzE8PK
Wyupp1KBka20QhUAWtFklTHVYYzZzBrfWQnOIUzqyj9ZwJlO85xuc6X4ecULUcsA+oq2kPSKpVMv
S6vtRE7xAzcG0bWXPSomBVkPyUpQRXHaAtUw5p/s2fd+PTyurGn+lduIe20Fu2Z+ygsoXHmyeEla
NvjNFCnjGSegbQZfcbGXIa3JiVzw4eaElRW4gOweydy2z4bWRVTGGqh2uVZnE0LaSHgWS4dOxVDG
FCsFqmTYdtL1cZnJqxOpprcD5gNEohq/DEcf1tDvKsAwbIGBwXYzje8BgDppDgGe+CwH5Jcal7Mn
N/L1IcLt+BGzEZ7FQHA4f2b4OJFyh/ZO/8Ro9IXi8HQ99unPVV8tMcaZKJZwB0ZQhrS7JUo+UWsf
qRttZaehFc9ydHWPVm60AXjIbTyLENtkw6URiESoQfXu5Y4D0DyHZiaNnGAeJgcpV9DWV38wBqdU
z27cezYkDijbn0Z73Y20LQV+/MsbTJ6ta/iXTSxhFSXV4JCmwxqTykoN9+8rDZZoM4vYu8a4/TAu
OVq+MqQ1r2ZG5Gf7UMaKu9ptjhzq1pp5HznvJMTc5y2F099OwCGVjNx70Obc7RUPe8DcSFGX7oID
zP6h0Rr627dcA8swpckTxaS5hJmQ3DOVGlE+rOoJ8BD1XafRMdpZ+bABSvkKLSJMuXZyYHbVc2gR
IhTfR89qnIe0wuxpiuRFlkSk5mb2efvxQMnkNS/MUmfPbmujR7pBCTGFneyuJM1WJdHEF/KxV1Mz
RCqCQzUAspZqfHEsQvNqSldFnNKoF2UOyf5Ku6NP3YtPa3Xviq+/UNY+Rlw9lkhf/jIGqibsCj8e
m1ebY93RaKKTJsmBcNKnh3nkrhqypRce3d+OX7rVnnsf0ae9CTxJUA8Xcsjc5DF0ohtK9StrEqvj
LXttVmYZjJBSamcyXy7CIcnMnT5ErK1cUp7p3GyBz0rvKRw+LuPmUkswLVsSxNv14784Xs61UMzJ
eqHtD+VaMaCPGAH24JQVGs9UF3X0XdODHdZMAjeWcekRgDZfRy5mzro0t52xgXYwSvTQpBbbBmqt
wZtFwBFD9+a+VqR4HtUFd6iQVU9JnpYaUmOaHA3oMImswNZcuidBpObdTC4ZyGqRZSaxbzHJOrqx
oAh1YYi2XOEztE1VxOolr6oZm8G6CoTuyPulTVBmiEp6HIq0WpYyAwTI/SUxlaYoAehiCAelne0W
mLDHkHA3ABngf3xugiLJcP82O/ptbCj213/czV7YkfyLzSosKz1U8CTXuuIhlbpq61gabbrajSVf
xuElqyS6XmFZgdZihNcsx3mJj3i20UJLHmNh2rYXamubvnYodBAWZVro45+7z/A5krtiPswxs8qR
9T6+TJOzXvxd+4aXO8+EI8BbTbzdkHHzhnMonq4YB367ArwhaLpCT0RmsloHXV9KuBdLUxRK7hn1
TgYGudARTVNLsGtnoxcmIJqGtf1J+2n20ZB6cT5zTVrsBhdAe9+2V7EBTWfyI6AuYeM6ldLzSD4U
3RH19HueRmxth/xYoQYqsUc9iH35QBn5dyyz29lioUnB6NPQ4K27atyStIuu7WDnCRqNxH4cT9dv
pv69TnBNKwUruCciAcdFKQb+nSf1MCjfK9Hp786aBBeftQwJ+Kywf+V57Z1TmmSO1qV/EIulb74D
1qS6vcFmIwL3cs8oKk7nED4Fp9STXHlAXCnayIuZRCyvfMpHtX7bBCpXwYinxXApdl1cZXCod2IL
2U0Pdb8GPMjSfsGhr4LNzV8m/z6Oi8a02BvXRGXkuLp1pcYwBypec9oSCX9P1GWsb07gBw9/qS6y
AMLQm0D1W8k9E4u65rwE1emd6sAA7sQMITlil12acAOHjL5fVz2DaeJWLysEr2+NwrRlKTbHlUJU
c8ugXijABJx5CesNS0SJDvTx6o4qinsGxL6+ivs9EiWTyRIzOZvKRatnmP2NAGYaLMGz/cJIQoCC
8lXT43jRNGfy0TNHzhPbloPIPick10fW/fbfEQ4RROH4qpkXAT+6wfycHevxzMSptLaOYjk1UbeN
WwZZoMNxSIQvpuHjUtiWkcvVtJ5ENKQilIMWwusLtRF8jDp58sdA2GFBDKRqIVLOUXtqvb+QUXOo
53/abJzr/s65zoX9zMMxn9ldGS4AECKSYwgcSbg6PkVQvdWyUiRk/h8KLzQxsps5ZPrg9m5KUhbU
swk/U2Mxhi5Ehzq44cGKuBgsuykW6dYSmpRKL9WUcYdEXwArNXuLz0wVPGikgd5WhJcLxXSmVmZK
GPI5TnVHsC+F5NdgmG+ZAztyMfEmd1JwPCX9ZUrMuI7CCUj2S806Z4Z6Hlfgt2xEtKm0Ugl1XY9g
vpqCOYNEllzYbnbPsaCHMt8A8a15cC/HELXUd8LNygJFw8HnDjahWwhC95o7hq8GrTp1aQsLwE+w
WN0of3wn7EbHuxQDuHO3mojnJDgGINYLDqJZiHJlSHWfzzIaWyhqTT4RqpOxg8RB2Q6Bfp74ZLbN
Y5q4rYB2TxHDMsjDJmaqTHKHFI48IBDvT3aJtncNd4aXYKKb1QF+BLyM8H26gGhfS3dmwXIqxxqs
NFG38QgCVwWr6VIR3dBozX9N4xiZkrX7h+JcCIt/FUrsA6CeJX/2pJbdoMhDujgyWrCDXjUXn0Mv
UFyOadyq0DIfmrRWgewHjeWEMdR3mlWomXBOKEh0PlHk7mOlc6dddaR5e10adx5sQkpKEPmhsZcf
jjm5r47zPERRLJ7VGRIER43MXL+j9AjYO6Jz2YQuMCSsPh0zruRYgVi5CWOBKOTxPyVXyDbwbP24
Myu2VHjWWlQcJ0ohres5FVzMFMikVeWhYQTD1WRmvYDb1ckVG9c/NvvrFzf07Vt+hj+wducefDjC
V1XUvsNL5QM15dE0hjuMqoc5tlhM1752Ov8QH/HsEJvpiuW+fpG1O4e6DTiTg0XN4w9gvM9p+oVu
qScs6f53ngh/p9oLsKBLoBLcxS+0ivgvv2IoXgPJp5SgN10w1IgWVy3EniacTBiyOWsWdkPFNF84
MJ36xXNTIU7AH9DFvnhvirP+vzX8hgsIqEkE0oH3gI07WdNNdtV2jYwnZAIs/uMWJm1n2zfa1qed
HjdgHC5vaiag01/9gZ5oUy8vXDqS1kMVy1NGH8bW2uWmqUTW+rnS3H4KU0Y6Wxk54KPK8dDCo83G
9GS3ed4niBKgnHLYFeIrGEon6KmaAVYP0ZIQs8Krgms3HeFvIclNM34SwSdPjqZVc6Ecz2YQNMer
RsqwTEck+XYWjSvhSeRJnZAJ7dQ/n+EMqPyQjHhFTcnjM+2MYVpCRPSVGXt3U6HUDqAQxN3+Oi0L
y4XvQy9ssyLoLdVdleRC7BOQOzXnkBbfHDjK9z64v/E/5S6sHTCvE4pveSIO4uk6PMsj0u0ZBFjK
dtwUvKPa0SNF9uOj7lN4ogCY3gYC5SB35dywSKSYC9h6cC7kyNYGaeuZVPB55wM7D0NnAHsWDxCd
u7ayrBlLY0KAMNQPsaxqHR3ItfZPXbmOuMHKhCxD/rJ4k9HAFW9eAC5weEM0am3IXHx9WDVhFecx
dSsUGzqN2xRcwUXF97f+hNGInABUpuJ+/Rlx3ka/sYsRPMcHwsumg95pcXwiWgTFXdjTgS+fIP7f
IH22fgWIrJGPbG9ftNum8CNJCT+hAPJqtCjvy3HtrjR2z7WkcfUnislZXL56iiEZY1iB92b8603g
Jdb5kP6IId192oVNogWcxyOv92cvZdTNfOd5zoASt8JlJaypEsGJjzCFTEm7/aZqpYTTxueWL33A
voBy2fthhoxPcdXjxwShRTpuxdg8nlWR3vTi7at2jaP/OG7uW9q3JkZpGEgAhyr+2kMVGS2nntAI
LFe/0/xSGUYhA23go0ZKieIjly5L7ZpfHDnpy0duvBHHl525hhwaGaie4zvRb2k96kI3CoKLtE6q
s+mlI6BehpNQ2aii6x5befLITXinFLyY191Y7BuQg7i8llzQQO9V8nJLWYzDr8Rc4suqTmBwQ4M1
6HnmAFmfeUKTeR+USIwm1ULuGPBst94YMmoaXUY/k7s+nBPo7jogyx1pCxQ5BCiFfR3Ug/I+0y3j
rdrXAThSGQz7moZWNLiTh4QIkDPoC7uBHmeJVe5sFYnBd6hPZAcgtGjN8YPPj84fnX7JNXqq9d+B
9GOSJBP3C8DnyjHH2KUfJOEhHg0O9MGjnBk3gDjQxEyFelasUuF1WqELrA53C0R2XzI11bd+2oUQ
PGHrqWXcb547PlRLnoRfcXEBtuOqpva2I4PzSlikIFaIek8+lL7AR9d9A6PDFVrcwHK/0Y4I9s6n
tGYxd9KqeadcJFELD3oioMmEuE5Y5btnNOwYCNFjrIbb1KHTc6Rg8PSDm/X1Hu0WlRfPeVWu/+kO
Nlh1GMpGQryzu7KupxLqqIaxNa8m3UuNvoexwPLYwjWd1ihN/H1U+77rkO9Kq17qWDYGSAb+AesR
gw9JU+bax+lId4zWbLVKBaF6/V3CWNmjvIpfHWw1L07lmg3OLqD2ZbZvR0xKy3sOlW5vgJGXZLJF
fpUxPaHtpXyFJ5HsghTpU9kPhYhEm99pYs9Srn6YSQw3PTRanM4q8w0yykGITF7LR0zyu5ZK+bzd
IQVpj9Cfz1hHuhIMEGaeCGRRiaD1/5CeEsVRbcx03pjHfXEVfKG5m4DfnjYPIFSDXZ6nTypPSgd4
fq9YDb3RH3OXly+wVlODDcKDyynvC2f22aifmrHPtuh+aGWTXShqMRNTum9b7QFVS1qwv5mRkjtt
dH2hpKfnjaaN85ei9YcJsBpcwc3SjWoK/Dr5GOOQgTLM2QyKc9b6Y/wbvPmkrgiv4b75t+AROZwc
HHMuQqdUUlT67P8bbbKHrTh2m2XwOgsBfDkEXz6yzMr+HBjj0hkKdo5hE2Bbu1/UOoyYcGIsCoLj
6e1Uvx8LsJ4KWa5z442mRMd6i5LKVj3rW78uB1MJy3wcAlvyeQQHCadP3rmNdDg5Kj2gJgbvSCq7
IUu5dSY5K9nf/n8cG8rgsEDE9evLMJnrK9GUNPgq8CmxuOQ0SqRsvRcDrC0H7MKhiu32zs+hh4Z5
m+oKE+yXXoytnz13IrqX6p/uWgeGV9D8PmZ1Fn7dR4lLt1E1ns3/lve3t1CxGVnNxczP9g1ApYpH
b/wNqb/o+/g5OdBLAxzHhF2HImH+dMvmZUEOO8Ad5a2+wsVNaLfoMdWDM80eqcaY9zAp/JwGarJQ
d0fefX/MO9RgZl8eCHrKgv/eOohQekvToh45eNQ6CITkmze4NsxTGpSoLsbMNx1siKxaJlVZW+bm
/wqTUxtkUpV6wD9DL/Ie8rCLeC66RMBrlIgUnFRXI/Om8quJVKEWjXtWEybWV8B0nPcIfmNuFuFt
+GaighWyJu55mud3EDDgXquXI9sgZTibmlDQ4+eSCcAvGFEPu+B4AEJB3xp388ocNOeUQUS+X262
ouTfr6PUvrrYIVg80kehoHvRzgwMErtpdMUDqi2ZdwNzg1pEzYkDid+SFCcuh1Zdvsc8BsnJ0GWs
ikitNbqGd8W33fU5wcGs/9iUSD5YieTI9C9HxtrRJSzGshwNeE4Dv8lXf2HTJgPhhXGNNs12NcDI
Q8P4HC4lGzAiNcKi4ZyQ/smqgULp1Rsh2yG2KpMfnTpz1CkwiQ9kcBBoAt8dErDHXQbkOZgxcnrU
0CqKbQ5rH8R1eIcw0sCjkgXo+jlTMOSh8K65csa9YfXfQebgLb84HN7NvG6jpGvsaVgPI2H9ynHs
AWiqxvbvDYP5HIScXIkEQFE2iTuUx3qv2V0b8TlMLmtHSu8RqyiXAnFgNWA3/UvKKVLAne7rgxID
zFCx//ERLy7aUkdzzCe/Rx5k6noSMYvl/GN8kSztOxlxo0CLxj66khk5ymzPs+uwUGbw1qryCys9
jBKs9qsls9L/F6J4Y9y/Sp4D6Mqpf3l8QdWmcnpyPyhqlLl0Ue+9kGOTWgcJ+Jg69DivdVLv10Ab
Cd4APD73053yTHGZ9TMAm5beQUGfD1/7+4SjOQjEv8TZ2AKkgZ7FSX8sWCi+AcJ5E8c3GnM2oEkT
JCvvPHGB2wE+qko7VPfLPn4NOLV6vkIC+EHsO7fBtwyPpRlSlevLm9h17R/TU7VP5vJkGKxVWnPV
kE2wHeSUqwOD2kDZ6cW0HpkSozkn1XlvLINSQ4DycXce5Xh7g8d3IS3Koe0wkRUMmcaAa3A+Nw5q
iJqgr6Ym5lsBKHnT+2gXDqh14CDf4pE+uBtcieeqo2LgeOdDDXvuBiSTwWMlDJocMwLNXvGdAVgS
l0pEWJDQDCr/HZuIkSvVjbpWe4nrYvI4PH19eZuZktcKaRmyNBPn12Ma+WAxDIKoVBlqk+PNKl/H
kH+7ydNkEn0oPPkcokHoY1PYAZExvDsmV3A4eFVuvgkruiXHLNkypKj/UOEWc105UW8V4sJaMltl
hXQze+jIDUpw9NB1U5gwkFWjyO/5wtV2Xwfo8pEfOhd+12fEJuH4utOQS6hLCOdDLzTZaJw6i7hs
lINZEUFwpnleNdX5emr63MWDxml0Gqr6EcybRBG0/0VY8Lymn4POlYBOWFS/cE0M3fCcOeJboKIO
ZHzl7JCeHcYhqwKZKcMe2CTE29w0+pXp7KkMKBJQqwTb06JHgrC7wi9Frxx1pJ/uWcN6kVqSjfsp
QY1TLuaZL4scUEn37f5zBvCJ5V/9wqPegPVWn4Ku74R+Rn54iVjNkxDPLO+UpuD19wXSUgjAzEJo
Pe8YNWHN4IkuI6ofclCv04xzOlC5dCRnUe440pbZVfJ7V+DWVs90NdnYqSpvkGHsiQjGM4VeZK+k
YijH+wzUaVu7HJfNyVQtDD7WEvYoTnI7Kkma9/puBybP2+Dtsi6/KP9RU45Hvo8MdHlhd1tY4kN9
Le2eX3MVr8HwgbUBNVxqGZR5e+MPo6NnXcEOqjDXSEdrC7fTnCgy2vkyLWHT5qZ3vpCFq5pmVEFo
cU0us7ELWeLfbluwi7tnGfl5tPgEtr6kAB9HiPaDoZRWuG04HjnYYKnGeS3xhkR3hDpum1cWq6Tq
w+TOFxWOEA4vfpbqXKde84VROmxcYpJsGCjK2FiPcUmw2FzFpPY/fksrR7m4xkW8GBRFbqGFW8ns
QvkswlkokT5boSfsiltaBRSEhlpb9k8gEKjNADiIM2ZAWcDZbzDAZ9Td9XrBo/zN9FO5l9bygJ0W
060RHjEZaIbyu6ssFjSraiO7s4XEvTrGC+YxHG4t1fCXtS3nx5B8JBnh8Q14ZeoTmV+bGBKiE9/h
bydceh6l+3ZQR0B87sBGQVm97Yxuof4voqq4RDD5kWDRtJG14d9mGEqQzkOXjEp0J6PZ7W6ul8yl
/SNCD8RVR1GJHsbnxVN6uKpWf/Eg2qi52/LIBfg4f2rTbOX83GPffJ9A6DOPTs9VHOhee6l1qz+B
SZloA/s1d4JxNgbi6iiG/NRc2NOYUhdojat89qbBOb+uB4n9ABlLXO2D98IbfbaienbPBPf3n+uZ
mrlhMlBcUlaJJFKLD0rd4ff+jKVYmbA/Ne7Xc2RIqQDHvTRQeVjY8YpUJWUVJKnDxtwO0/BZ0/Zt
KwaipXjaoAPXZveaSvMrndhLn6RThDjMwTt7zqlrsWuhCv8JRYy2riNGnEl1FmUUIe+ciydnY+/G
cqNBk6PgeOXSiLvTbrFHA2ZJF/nYbo9ZXPz1/8FFC4CrgpsZPPoHN/TlsucQeXlggrvAIJ95bkUd
8GshnN3CFqE9I3IAx1WFpT4OncoeQdYZB2T+DREmAWn8JBYRMwf45fw1L20eXMGDXW8MHaRkHvdw
nqkBci+3V1h1cq2mkuB9usDY3j6r9ZiSBeEYmXzQBDNzsEtjmmtFj4tHL8ig/6ZTHZ8k7EXhDCOj
GtALGaEuO3zAJfDE4lP/LR7EFJlepGgy61f+6wvgNZjWaS93qlPDnpKSeY1+8J+sn2VRcE9PLWew
hiFzkCFnhMAphsyhpTGvy08KhB9G2upq+bYgTlU8zzSSmKpkpnw394nGENvGosvlvTbA5jeks3y8
aMeH5D5xJ95h3zZZ7qRXw0VDpbtWA34rbKN0Hv5Zvw7/qfpH5jX5isfIQtJvYrWtiRiuqVSNEzXa
uhUtTs8g5sYxsUgeEtgilzWw1VmZtfcxhgv2DGDqfNO6rV7tCVs08uA6A3EVvhBnUlsklYd1ZMGz
rlx+2nT6eWxpCrfzfj1rln7dC3j+TlE5/ESeaQa30Db+I32a8FDrIe5/zLEFMwS0Y2DLvDzRHkaF
59s5zpJtO5wHezQNAoQFpSSNgotRWUo8ao6ElKv17Lvk+fUGDH10EJ8jjochPWQVR9fLbmc9gApZ
CdrZGXxzfiq9I2C+ADsIkB5ZxUZQiAUM5n4oGY1FqUtLwYlhFZSKL6AScoDkrG2fJRnxTdbz3sin
g8oJS4eugIdwHb0W/Oamw7pkhau962nAv8w8rkHANoOwXoriLitR3W+pKWV2SjlZ1LxxK8lvemY5
af77JkBu4pDWXODeKwljS/t8JpBGSPD1Qnu6A69FLbSN7Ml59OV9jcTOnBc7R4xRztLBzHenXVeT
x+L4+xILlDg/LGuUmPKUB2X5rTAq7ZCsFuuYqqOc37pBQtkI2/01l1O+0bsUmUWowY0MUB9gM/xo
fjoHsQnCKP8YVXMckz0i0xgquRm5nCThCA4Ke7wul3aF3c1Dq5QYKAEghz8x5zQtezZonz/6zOZ4
frznn17J+T1D6/lutSyFW3hzaMRrpaeiPrVLVyVcHDOVJl1VnKfc6l9Bsc/rKiUtpzYlDz+zvPTt
KRSFsdJ3hV/OEPyQk8Zp28Ay3to40Y/kXxuLrJs8JxUuW3oo2BIRwY9KswDOariPre82yD7SVqFl
xrz/n40W3nijAYiRk+7vbac2dwtb1HDdiw/BT9l8ikrRzf0h8gDjWxQ8XrbOwkd9J+QbmPHHl3Na
zSXxqdImqmJKxNKtGDvs3vkWij+Zj/SbaBI4wP+1ZfpuUPODuPvtWmuzGnEyP3YoO6U+f5em16CO
iCFattt+DhZ6t2bWOssuI/zjvItFVfX1/gTCOtv/2oTRrZ6aCQPCPpuiyIyz75bG1MiiBe2fOi4P
k53TlZZSr5PnU/v1Q1UT/QLaTEU+GsgLUfRIkjDrjbZm5fkXBCch9UUCv3jcXxWunNAv6DGEYxtF
Fs2g8SJ1f3iBoG7M8UTvcd7H8HQbxsnD3v6zN9oa/RaM4GE/XTHmXQvfMArpQF5tjXNPS5S7lbmO
D2zJU6OnZu/XQTpNA2lGZkV2tDXeCiw/W29sRpaDYb4iFnNYg0uVXHLszQbsxeo48MgWUWpFMkKG
BupZ0CI6peYp2xxkMIyi7+sKuR0RUVAgM3fYCCjCh0DMo9hriKbgcrIcdR7PLai2cdfq48FHUE1O
qOjl17mG30PZHVu9eoFm5BB1eXjEQWTpFEDaYC6FGoOAfaOFgjZ09F9pOvWAMKTR1LrbSD0L9ZJr
5N1HI5hLxOd6rvslxtXcJPKNUyufisKLeO2yA/ysj5FtQ+qh8B+p6KJHSxJ0WsrVtAFgPWKd9UzG
JcYCoHDZ9PDDK+bZsqil+ZtOVlhpG/Px82jFj0dxFvEHMYhMNRhFIAVkoCv/dhDbSZuSCihVZaKJ
yHz6AxK3shbXIDgI1hOlKMTBIJ3+iKcW8wRLRe9PZOgp3a5O6w5aM1ZcYjyhwMVVc6fAlFya6suf
bgO68cA+KZuAHd+YoXUSrp2KIljmsGmlJ67rAlVJusVS4P+8+iNS/hnDuwtzf2AwcgrV2NNDxOBw
j7RigMiH2lel5+/+gC9yzlt6sLauPmZtuZ9b3iblpc6JOCfowJLGZEd8Fnly1vD9MF8m+8vcHcX9
IIic98omcmrESSpcaWCIcGzmfC5QQbh9oiGYAiD5SrfE/s4luC7KRoRseC+mi7UO4gXOGt79cbnC
cHFXEOkV73XAquxm/Kh7HB1x9k5BWB9ZwstpNTj/uibo7fhfTt22qjUSPYG8jnnxW2zGv9zdXdIC
aQd2XXPsCi8BR0DSGWYHMA2xFJ9Q2xhcjhzaG08bpCchXULGJTGtclrOmtRWBHRtGrpMXFI6tvs0
5bBpUxI5GPR6FOGBoKW6JMy0HGKH8mtvFM5ZRJfpiEGchtjlJiFF+OWu7W/T3Esn+tLv6NHaAKaO
CA0Z0mevGMi3wwFbksEiqCw1FR0mjrPOQ8SRx6GIKB75Xe6ztzkmA4Dw8yJyku49M9nu+L6mTKMU
LJ2Y+WH5CxdOfNB9n4oCGxrsZtvQLcDgkyWV723DJQjeylC7J8VCEiQllzwnURhHPZLSTwwd3Axj
L74LUKDSNWVflFOkzaNg2F44TKbG/yyKow5atzLk3GRtITK/RVRLgGujzQENKO8vqCjj81oBkd6j
skKQpH0jsxynpVakJkPf9ztfwX1MlMuHtZ/hqOq2TnW7d66Nr1o6tHfIIreEUCXr/VoLaBDVIOuN
JYF8JXJM4yL3jtkHVDCDxGqdNyIrbvgenuMFc5pr2w5DlYqLMVdS+4ZkolbpleDiMlstrw00zWTY
PUZiRZNPU42Zty1ivm56AUkSkNyL9UHR6tMca1Qc+moc4ZVIt0fUvxQm0hndYS8nI6fpPpa+2G+Z
fyC3MECf89vF9PuQtFVNvy9XqnuRBLLdq8GHQg4Y5xNRrRj3jLR235vlPkcAJ0SjzLAxmCfydheP
nnZxUtqaD4X1XKmkEN++8bDwkiLxFoVOICjfKL7P1kcjYHs9U9AiAftb1K8A3kO2BNaV8r5OJ2S1
uCgHPTAVKgPBreD1qE9Y7TRv1lIM5NaA26jGynjqGHwWln4wQi9DB8iEqi6UQ3VJvb+0i2kpj1pa
Kxg6wiyLtv0RP4KbFTVoslj1w8yjJg0wEqoc45+M70IzaysmTCguo+ZX7Gg1+hzyjvw2GN4NpeDr
WfRK1nkbfHpChkc4kl6LaRHxJYfyXwD/iB7JMIikghPv72BJuzmKZjD26o+leLyKlGJZ2XLqnQ2p
6T8sgoqsmYueUEcz3jdOiVtXhlSelRSRlOpW9PxDNzGpjsK2129aB9ggtCHjTRCqhTxYgAxjVhWW
8r0eFwRKEES+34bbRiA17G7kZKNU8eF2x1j3P5Ze8AHfp1ETV/05clkHvCNkYnPYMjwkKiEcx5dC
ibYu+XrFMoAiv2Hp0isPHlhYIRFH1OdQEdMOlAOSn8deidaMOfP08m4XlPqIuN+CgosszSyh5gD5
kr1J4YqLKDf2DYggEwdZZypwdkHniiv6wfc73zSgUAUKpWa3qL6oPFBT4WqNqGCagkd80y4635z4
bH5BV2qyhSQLNGB3HSS4RIfl/ltdlzbj9v7/Hy34sn/HZyJsNhZlpSimSZCMegxYmoshZZdHlkMG
zsZVb285nhW81XRtygX7xyOZhvTSdWyuqUrygXZ+j7ea+IEJS3WHWd8rMwmX8aYNBDmGmlLl3OfR
1QVTheObOAFMEFVJUXmIbCW+Z2hR2YiEDMcyLG2mALnmiKDxcUZewoikpSfDK1NuIpga24EiRqig
nvsM6zz3anLtzQ24SGvngg90cOwuqYUzwODs1JXO/UmKgyQNnHjFP6Q9FAqPLyqRobRDBeSPuJ1f
dQgAjaaLSomgAW5u+HQ7YlDbfXZmEN3jqoyk/ZA9c4umby42eNGvlwWUMcEJHj4V4jF1ZANKcEQt
2Ah36JoriVzBIukipoBNvmQ9iTTWFJiDf5ygo2QPNxwF/ets/kXk97ww7xhZEngGk2V6HWKmpQVT
UViLjh8Ndr62YQfYkXtH5HNl8hQXsjpdUdjqdciSJoFbeZo6tyGRnf6Kgi04PICkjYcFSawgyho6
YAyZ8DePhlookH5CMXMnOHKXaZ9PDvKGfMelz5QmLfYnK0eEn+WC9lG2o0ds1SzsYU7ykquzSfN4
4FKsHIRVOqAOUWp4dSZSS7nonBeKxy0S1Efa1KG4PXcQ3o2M6a+WHKleVmf64nixYZ1bCmEA7Lb/
U22k09GR14L2O0/dgfrXvTMAQ5x5SuN790HviOS828uP5YSiLoFzrl/gRImHEzesnXLqpJkxYikb
HIiaWVqAqaV++3ealRoqw5rk4LheDxL15yJxDCX9+mnVlIlNp10RFArS/Gvvb/mLqHOjQCEjdXwc
+nIY4rJTwimFGWg/UeY0q2RybR8EL6/AAmDNptKs0BwVP5BSBIEEUfZZb9oh2ZVT/3vyzoHhb4cJ
UU2nGvK8Ze14/BO9E6DzU3MJ9V6QimXrTLbahfLpThnmtAONf3WtVxKii+H8c4NeiBmD5t098/06
/3AlStUMharR9vXb2ysVTinmPBG04o214LAQhi5chNznwMBZs2xnqNVahFn7kUI/176+cVJLMjL+
mQ+pMZqCvNJIdCFYa0Up80lmzy1Kvx3S2qVHIC+smtPckHBTtymzJtMqvgoutLblehTkr9VDxWTW
2FzJSFe6i6ud1Ks4MbDMBYp9BAw+e0rA9V+RGYvnVaDm1tbRCZRTS7LWsvA10MfpcsXPI1uPNS1S
otlDdvn6lkkwXU0PjVrpDO/fsGB+oRA3zu60I8rUNaPc8Y3/x4AKeHgGP+55KWXa0Ijps/bQtMgU
xRcD6leAr/ej7TbjIK/lIVfcncD/SJCdYKaG7zb8BnakKPWLDYCpCGGO/2cW9jv5WgcDeSybO0qa
tQLq8TUNiSzPR2QokXhE72s3bwhbijxUMDv9eMLltm8VUeeyZRs3v5W8SlsIXxMANc2R80ILp+4V
VwMl66CWGKk+iRmYMA1qC5jmwQfTnut2YI3ZcGYuqyHprazNRr4muT6Tb+HwFb2Odpu2AFe8WLem
IFfPmEXIVHRqMlmMPZaqDuchIBo9Qip134y1sPqqijHbS8QeM8bsKJDPZLl0/LObaokfAhn3bIjC
KXEOZZyLVzWDyXOTG4/S28UX/IymQkQtrchAa4MAGvkG4hVwpnkJ4Ws6uB7v1QUPuwcRbXw+HPE0
O9oZUEX0GhbdvsKCeW8Gh85U14ql5C9spwH156xgscVM0rLpNjiUCvXo8py86o628QV9hfU7dPRB
tPo2obolMpWJsKuMxYSGHH7ey2b7lhvoERtMRtGBpt0J/nzwtdKcgd1f940UsCUeQkBXk0FH6Qbt
kbtV+5kyKK15FqScqnQU5dPkPv2JPUjj+zSiwHiTZ/mTH6luIC8MwdGVEacLPxUJTjZ3lCJF79tH
w9bNbUxMSxTrKwIhSImdHcQKqsrmRNJWKINeyhgmzcqM7zFjXS8aik9pFDk8bk18lzKfOpwxHwSt
6iABG35XFbVpAcbQ4mI76mEtQaIOp6uRvjrtLDZPj5eYnHF1j58hn6xdKyXWCjymf+8eoGshU3t7
wa51CKUWqr5xMZEwhcfCfdW6PTURUBikmR/VvHR0ArJ8XK/Xucy1nj3jXrA/GqKKVliR68CC1fEA
ViTBVKqwXg009AnLhTkUFD3xzjBdmGfybm9C0vqAkxtHmms2laiLoc9E4+FLkf6OK86TFuUyI+is
+7XSVFevBRiJrGBOsayAqvOeKg3wcBaIzL88HJkA/Ls+j2tt6PthTmzeTuQTeEgHhqVwb88eRBwy
xNBZLfgARUBmMQt5Wt2xCAAkYwFNMyUFLopZtSnEWTWGVVxxT9IVINFX3S+wDJAjpc5e6nsoTgTh
sC2DW0Uvg+WSgvwJ+cStLhYuMOQa54LQQQzlAbE8wIhFzc2Aq2ehqBTaJCPUwaH/NoKC4V8cFORS
DEOpSUJzEmAQOOvp8TKFj6iZ36GWuhLetIenFZiRh/KPjkDofO4stPeIruF1vtEk7dkBPr7N3Ew4
9zsJx7JQqYOSzmSUYemQpMwFOsQwN8mTGEqYS0MVEWuJYqKgO3Ge92Aaqq3BTcHS6uX4S8SgLmlp
arHKzh3zM9l4sXwOdUqjZKMMz/jOYjt2ySTeVRdM3J90nE11KmmQGKgSLT+7tD2mkev3ivvaYlJk
Tffn+JuSzEGY3/py8MobWelNMZNYHZa8jN5yADpR2WuLHi13Rtg1tkqr5XGx7B/HW8wVrGAm5v2O
iACHKGAuSs6L+MA3e7QirsLdi9hbZzXFmQgxmiwVuHVJ1va29Tm7KOrU6u6QdogzR2wRaKkJRlU0
dmXY7YXpY7qiJ+3BBSHaKAQpXIotqZXJm9PF/cdX0BBY6Nru5PjxZ67TinIAnzENgi7IsPRuJ+cr
tMZQFE5UVKT/tGhb3/xcS4nOD42zB9lizjxeGp7YASRA7CZLldvs910MyEbo+siwQnZk5hRW+Gnq
j/iUgRgSylJE6WjpkPsYar/SSBtBAZVydm0uBAKuGijmhYN0ilz4wI/TiEIRJ1eSj8nka4Ycbkjj
ZFj7FS08fjE51DQDsS7U5Uf7J1Tz9Vx40prxxPQ1j3mnQivgXwCW4PAud1Ka24Nzar94wOz1BNq8
eiV1c8ZNoJJc9At4QeiKj3ZWr7/xpojGAaUMxYsJ3j193/SFLclEpJWwBxJQUKNWh0fDkryDvQZc
ByWZr8jG8dw6ykSgR/RbZvc9GBvfj/fqhOnw4DADOxBxImBdHjAS+Fe27kYXI854hIHf0pWKZtQf
tb5tqHn0gS2tkXq95AIBp/cQs+LYqjWgSA9Z8hB6AYh78RxhzL01RkmyFqRkbI6K42LmVoAoLRXH
i/23lnkiUir/vbO/ujR5CXanKCWD0IdSldXreGXBPE5R9p3pFeBe4FrXsQE8QqU3m4356LqGG+FC
eknB+1F2Bmsj1TDPR9UVzt6sw8eA/4RLxXM3xsZLIO0DzddC6UrrKeuU24z2tU/ArEESNhULA8EU
sA1Pq/j0ef3IJk4XzoMF/EQ/5y/JZj5Io+PADT+6zdz8vkAC9g5G8P6VjOuNb51h1wMTVb6cpXZP
3AfqsTcJTHhOL6Z9gPJp0MoudRiWprbpQwaeEutrmMZtWGdg6czpwfkBOBLwUr6717O/6gH8jyDg
/z+ibpDaGVhujYb8xv3x4ht+Pm92vjVxKK9hmGqeCBFiXa7WDBIOpax/iT8K8y5Ae3jrvB/w9zne
VjY4asxAxbpImv8+gEk1rRM+aeyQlcadZc04JCGCv6wN4q+Bkc1gIYDR5gk+ChMVj7bahZ9dEGCq
HWDRJEcg7kdE8f7sOGR1KOojmoDmf/ZKGJdK2EojdJnpQDfRoFMyW0225cXqqYao8XI5NrLMph0z
8CQx2rJyxJUAw4FKdLJzkze8lhjyh1SwSFs5q5nkxbbPsPM5BwaD3bHuvzgv2+6ua8Hld736/eD2
C3Py1ei1d3NQIsM7zad53GmQKHkl6Gdnn5YOqXBrF4G3nK8HK/Zvy/NO4xNunHhdDGi/FU0UlHH2
IUXcdEON7eUgKvPSbiL5jB0/aWFZns0Y0RNEQkRyhCbRtbTBcV/3BdStrC9FbMSm0U8y7g7BV7qi
1vL3nKZuX4QxG5iqEmKieNZ3ZTjaih1eezKMgCNdqVzjTWg0AuvT43hqvQcmvj92cfJ6SNq3JRp7
bLSA3Cq3HyYocQSX57sgaar3CdArQywnWGdxQ2ShDeDzOif3aaE+iYyLRbhKsI2YSzICZuPrQG6t
4ot5jyrkZNWFuM7JEBI1pV1UmKe9Arh8zcIfBs50wAJrDJkLoIlBkYSUSPRcTabAbhbi92rvENYS
mBj/phes1eXAMK0nhq1A+UcxbNX6fdvPhNwtO5y2ApqzO4mzjQoxqBAnY5dMVfB1Zxu9vDL4ZcnO
ApKLQQ+mL+31DP6mqZPvH/ZWPcRXbTVYqippO0jYCQBZJMrKpPxLgQZbt1ExzNVYNwcQb2TI75nQ
slGvl0TDR5gItBZhpLpvtfvR/JGtPjZrkZpSatOi+uGPYsNGC/D/3HBEhSTBIOxrINBTGbjxFt2C
LHoadyyrQxB2zyLVBxGT4NpNCXzQri3Ay+ixLvyIM64pz4wAzvWvuq5WccX9wLdJyTHr7W+f7OvL
iJ7I/n/l34Rv1I9KmyPI8Y4wRHTMxptwpUbXKOq6HndDAKk2wTlhEtwRTA8wJ+kBVfxPJ0tQXly0
WujqQhOY1gsYcfL2ijM48tf6827w190SH0pvtoXh3VsLbWenVmYLRpy9vtWZS0mFHjQzcOFZz/U1
2qSUWbL7GDOOM6D9Mbbc3d46yROBG7pF2JwdvO8U8EUYL/YvgcNdaBWpRvXXP3e2vq0CwJHSK1R8
yPO6zBowXtbRaGSKK6dgn5oRDBdYHMiMiSvOxn2PWz5swk9vcJkUtYv6jJRdxTChB/T4ExdPgu6R
WRa8jyYnVQUdekA2zn6Z9/YcabqdpsZH8A3XadO/LW8PZAReqEeU0TipxF7Zlb7UD112WmzxgTHp
0sDTkCjpmlljLnlbPEKSfpcDNl6RvR38GpixIpyTKAl0h+yINM+OdNcDl9dACLnHX/67AyDPjr3b
6NYLMPnhGmMRvtwneyndKY0ZEzzLYWHhPthCh04Rzj2n+QhuelFkNnPdm4NIg3wIV9eHUHDhGkKJ
HAComoCtci5KpFV3fd7g4JMZh+0XCIMgEyQ8c583aRu23wLwz7YVVBPdABx84Ruu/McqiUdPBVLe
9j6xltC/dMjxU4F4wuHiKBZzLZ9WiryeYU2MPlsc5V+XkhniztaicjmlkGRrLffJi9HTHJAEXSuq
hZBfEWmrQL0lP8iTzFHHUFeXYIvKE2vnsJR1t5BzHf6ZES6XH3pHYbYR7xpXSn0K3uH8sQeG9GUj
FCXktjHYa7CUzD1yZYLYktVTiaoVnIr5YZKDZhRW7MKpCRpuM7ChcB1bPYTvHd/nuwlxxmOw9PHD
7NGQg0Bn8l7CTudOdIt02jyPK6ygwpGU+M2+RH2NgWChCZLEpu9m7tMmdmhKW91Z1ePKyXeIhH6U
Ie4HZhtRhQebVqMubE86rkq1xj43gsXJYzfcDEUtdk9CjUZi4KNtP5SaOk+wX1iSsxazKO2miAKZ
9zC+EarXNyCyavwO2FZ2bqCJcyWgRUT7a4fFvLuj7oQOw9TfQj/MTMUoetJ4QEcMdaxIY7h8dciY
pSaCseVBB77HaeSu0ZpyqYlSepEKz+3horcG2mCey+7dpv2HRHaQxxc/79Stczvkf2z1EMfIOrTv
ITWkTVKP9bvyJ20cOChsxJoP/dtq41y1tzJmxK8ANjQJnR7YNuH680mxhynERwxyxbKSWm+CGyrl
KC5H/MDt6PnGyXc1OMkOoNxBuMcNrLFJRwOs566FxyxPBBwBZKz9pCRmHbYzqguPcgyDtnc1VXno
IaADgUZ5WbweeoWYRSnH4ZdWgDrqkHkp26P+8/B27x7MH7nRSzFwYQI/dBus/ZD7e4AVs2EhD+28
H/05/osi1Pfb2xns1tDfCS3C0iTJg6pmSPVo49mcNrNjxFj871GLh2qBKm+FSUT5/96BC+gUPBx+
p+TEsZ7VQ62M9LNrWEBfmWj2M02FFtWqCVkpZXiclCMKFbRf/whsnYkYZnqvHrV3Jw4V7VOJ5q4w
NTiJRRKcEyhfmZpaIcc6YIaRrp3CZshV+MoewWtCrkQfxZnJinFy9OOqQBNd/96tBiUJufXlb5O5
mHDxmdM83QRsfT806CiSovBtrv3jsiJ37jFFU/TuT8UTHzqJbA5ruUa5YRY/QghEOdw3cQ2bI2G1
Uh8hOxEyg/gusnZEcA8ExPn9D1x9IYOPMexOMZr6s1nK6sk10+gmVHV5G7arCwDc37UCyJAz1HV8
YT3jPSwSgXpm0vFfbSqt2S3Zco/sDh0sTCXtSH7/LSXLA5M/FKucmwXrjuaDEnmDN268MWX/30k0
NB7smsq0hImaqBWej8yyLeBWhLt44Ah0oOqhZF/+RhfWOnRPluXfsCjErfsHZ7P5krdaNGaxyHZg
YS2DEvkcGD5EOyxK6waOqjrlocYuHtCCzEZnseeAq1p4na2kEBr1XKZPxHdnl8GL6smI4CQHE9Ie
8QeEnmRdsMyph6XVwlOiAloWnfisw/FMzzuEdpU4nW7PZ9fdcdZ/PclPxDgf0UxgcPBCmGO8i/F0
zSUULu2claNtSeMDr8Vvv0Wev8caIfT3P4yQQaCNwZ3UFMrmGMIKHdt9SS2ZCYke81nFv10jDmyw
/nEX+/SO7UZVCnbHEKfhXLMJcDX0pkJfxgGZxYhZUXjyAMTVA5i4OFp+QuxEvskVSxHzJjio9crO
QQIAJNIWwzZ+Ayk2/5+LQAShRYDKBa5ZesMBJ6CcxW+AL2fwBVS2AZxDEdgq3YBo107OA+Dp7xMb
JkQYHVBuQOGmh7/gya84mntEfW5p4/eAgeaJ/xR1lb0/x6Z/JW1foU9yBT5iQLZe5XDbYN2ysp+G
xHsFdwgvdpM6Fou3/Xxoq7O2nEoNwrm7jE7WygRVVtR+bOWw7GYIFjnHGsnllqghKZtb8WQjUEN2
wr47saf+8FGDfm73rGtSdW1d95yj36rhHLlcMfEnFMWReCh8JbIHRJCMlmCdRpDuforB9rCfN0f3
LXElhJHZvVNu+PYs1+OLnS4JwHJVkm7sC6ZSD9S+NncPZ1T+ADbzBZ+evNIl+zPuMSfgkICX1iPZ
Jk7k9Yb9YmyqF8gCTr3u+MjEihRSA15tWH2gyDTRDPUBA076EAaE+LrPuJ4eyFTT5eKTFkQ0JQI4
xE95MLfs9P8a/cziEKxbcl0pXnABbtq1L1Ban9Y5rgdL8nTXbR/u9Se5i/aS3LVdEr+JAj5yCsXk
7VT0zOsgnBOr0+hPwx9RqY5AhFbc0SPdeQYRbA/RDgzltz+Uop8Iw/DKLNSzIxHNXe+5gArYZuy+
gAVcKIwkFebK2rBg5+FleiVlaj17ZqI0WaaMX/fbGHMHYFAY5qAywCwKZiK7phfQsbTMGt9DgXhM
CNEIn78hTvmCe90eEgedIC+3j6rABJDOhd4OMHjkIiq1wdURGvNAxJU5ovPTgWPILHGdBA2jC0Xo
2TlLxBmeqi105x8deCpC6ncdhgz2XBggcqwZXgucTp4lzXUBbyBmxfAg3zl78B6ZMeB0mtSRy8cY
9c5GrwJWmUfmzKg7PX8LKh/P6YkJVoA+ytdlmx3Tk5nBXiBTmCZOv08lBMlI9HwlduRUs92THNH3
vlFSQv7zT5iPr5FQcmi2tKNegfHtFYaZ79mwlicsHxCMAaNXE/sIUnrGBMi98kRTkFekhxr7yq1h
sW0vJt3eDHk8EIu5rmTjaXIEReYZZU7VrwDa3gQbWpt7rhdjMxe5tuhZ7qUzjJDxFakyHAN8Wq5f
/FvtEkTWJEtE6zi7mm16NGJ/Rqk62TCTAWT/4DU+MjVoroEimgRfV57KqJnffFe+dnMpih+IBRYv
PKU8AL3ZL1mUtIhnmKWliyzlt6eM7R7+tWJNro+4UH81Btayg6jMy7Lqipp1kTxCp/QzW8hQiFw+
9sX8tu7P5kDnV3mDAvL1LV/LYKAHyPUkksLEjWEtvHXQ8beKMjP4ma6/OtYZrB4GA3hDxLdEfx5j
nPUkpsp2iWcUbJ+dRyIPGIteYqPi6x8N/PRCevYNYsnx6gccV09LEWik/fU0NNr3i9n26bD9X1+s
amD2xuqoOQVw4gFcEyN955gYwEqj3cogdb2EeplwJcQqfVhHJ8pxF4a7kVx8NEaNg9tiSJbclwci
kwbPG1MnVQAfBYMkuCJG+5pm9kx4c2vkbdt6vapBh9Aj4MQ+O4aZ8G/vTNdfBzF41qwaJnpraND5
d7wmoDB7xvCJsdEreCZdKys8FqgM6pMi3iBSyLtLHOqACZjByq8x7MSW/4RvL6njS0NQKWZzWIBo
eC5Q2urhE4FnXWt05Ce46cCYHEbXoK+CdzQRqrq2zxIwhcaZmzUzEOOf2l+cZtNcJXKfUMKSpheg
hdzdH2ya1EME/xOn+LSKGag/23nFwDBATsoe8fUgGfV5/4eCuAD609SYFUEhDFCZJe25lJemAxba
7lOEDHSqzZJteVxYDBvOZbGeyOivCCKn8FLe4p5QwoaazQCTNEKUHeDTMp/32NW/qCC7i1MFsDRA
BOcCZoacQmyo1n8Elvmc7qBbzn2lTJb3mIQh2hFUs9/n+MSpcfOCrmOK70XT+LhEtSRxM+gc5Vdf
eQGBLNywAE0rKJj+uKade4tiG1PAWKyh7z5pPvTWT4BmFUWonE/M9PQQwkDKTthFeduaLgH9iiwa
InLIYHqjXa/O6rhfUqDCTMLRg9r/Duz+Qg3onT8SxM5Hr/e6SEKUzrqytPnR4ynkjcROOKOv6HzA
ZC152JknN2xrWYewIBF5JpwCaUEqhugDg8F1IoMiJ14w9Y4kQxtPJA7Xk53ITBj19+miqTyMokG+
kg+JSEOZzKB5dRKmFcGeKL+sIfsw2/86LB11Zg5grfVhvA+4Wjz49eSY/ZS7QBjSaFTJF+6nd/Wa
HdvBbKP1YUfkO/pf1RAHGlZNJcj394P4C3sjzWM+Bex1zyfiE3NL0MfTFDHSsdDlx1oQwAy5FkKB
f8FXIeiTjgdQEj4u57sjN0Xqn1sOqYMaF+4/OPreF2mG2trdOD4ftzICHCMy2w90ioGGLoAJTJuq
11hATo5Gzi0s4a6GGWXbqH4/T3BHDwJQLctK4GVk7czCDJ+OvcWlRBRuWgtuEpZwCIuYoGgI0+cM
6ABi138+vsO6CdFfANMZSaepO9rnHx6OsH4cV7Zz7o01B0GomexCIBZKpDdOuzL4DfMnAWMw6uC7
oE51RoQicBVQ5/6azypr1229KbWRO9s0duWLn0Md2Bq1CH+aJ3gRoByOUwydP7iHos7jM4G4joJh
lCfJC8pRp987mGbySdaWrzt3DsuY69Zq+1nfRys5S01D2iVBu+diAyGgO6aVTBeye9VsKwFp9BRt
0Ola34WeDggRjXPaLfYNI3t+Y/XWZdYEPwUgEHB0kB6N5okLqIUNFSE9bR24rFSyZ/7/IeEPPGBr
laqUZ/LUXyLQfmiFlfq4rkXSgoFiXtG00idVhJ6WXnhrRi0iJyTsDNB3bEhHgEIR/qnlXjib/ScP
3bgb6E4TDfPi2BWrsS7x927a8ujU9V7HxTJw4lw7bILygrFGWeW7DJr1SNOX8zDPrQFnKSe3tT5c
gJIMVMlORcUz+BdVAfgzuC/iZbQhF4lDH6NQj7RPgGbOtYW2M0mb/upSUNwBJ7+3Qmo7Yb16SNrd
rn0FV+1vPNncz6WhkKh2cTSKwALfB2HovcYRkWGH9z0lMlQPGYeHGsk82FYnrLEBL64dBRuT6U/8
dK1D5w2DYwVTVI70T1lVuCAtUgJPLgVcmKzBsRRRyx08REhYQtQFXFpU76jqzhjAF70WzyTDkegO
6xFdq5YXayP527tyhlUraFlYlv5JdJK2F3YPjFMxuQ9O7lCm7FEyAjQLhv+W6aEoxR0EBsYiTgH1
O8fgdk/8h+w+VAEvWVkgfVBdQ4GngiyPKq+WDIV4uQUF2KLlHURaq7u2vDXaZplJBIKsxlG0lV4I
BQqaCPaPQneSF86N1CRoAUrOSAshg+Mzgf6h9uvRmXwuY+n78Y/tSeE6FIzlI/jPb2OmwIcPMvl5
0MvC+gpeDatmPQQv5bUPiDEIm2fsNSdS3AwIyCcLn5ine5LDyho5L8UEhC/swEDgI+UFj6svE7gG
p4xKPJ9Qv+o83A8DdXtiW7wMWM11G+YYsB/joCsBcMy7roweP/PEXC6lOVa74aJddnEc17SuqKJ2
0NyuZEyWPUsLpArzZKKD+mvkjqt42erLXidrTtk0wR3aO/4kJfhzP9VZS0R8aKRbd+meJjQ4Y0tQ
Er95XiYDrm4mwZIPzHFeHteU6VQ/ds3uiDRnPzeXwbww+BenFRqGr7AK6JhylAdfnmuZNm0T5bkq
G1i3KNLPXPwpCA4yC/tH+ZJ2rNXwGQT4hiopJkf73kgST7vI9iywN2OWGEPYYlGp1Dv/j5RtABYR
62mlGFgcGdz9Mq3qSWjjg3ycr8JL0LJa0Xw9IXOR71d95yq1gHv/OwQBzrxE9n1g+O3BbjWYrCxe
fia5SWoGceZIZRcUWlBADsBEvCO+75hGIDzQ7n6x+Db8gMYDWjTkaCq3ITWC/gZ+YM+68X6rSkMX
AJe/B5zYwjV2LnAwlBGJuUaZoIePEp62lYHrHLHmFJHXrdoPvmEVVpljowTyRqgfILtYBCKC6Llm
qz+XGVxzk/dMH7n5NRz4GI8Xxony8jqM44UCN9YlUPlTZwvzGiikLJ0rFaue7pHE+Mm9kMP5zUa7
8CS22ibhUvNPkyPP1SC7CQm9YAbPlT80ziSF6CjezR4lVkPWUytVQ1pKQp6NblqwJCIC7yyu19lY
pCPBfYzWeh/c5ojZUt/xSVT/CTctwIICyIRlAEGp38lhZeLXA6jFJNlo0ISEovHhHHfwYQtkI2p6
wgOUn5ALNQo75/vmh0esXN57ZUh/kOhcqvOmvIayDmoDHLjhN+XFeECAM2MRBinQimRlwo+8ic0W
nsE6oy4orxDb6zKguiDOsiIGO3p5QiNP6CDdTAx3x3+FVXhlz3rZzVtcM1MWmvaVz273XgOYok2p
edKS8tyKdVOyn9AKnR3sTdUbmJ8KjnsVydvBVw4qfO9feXnEGHyBMbXJr3yYUKTqGleowOogK1bu
mIy5miaIRqTA61KeHIc5D6tb9X8UktP/pd+5jEst7nPUD0f3FLYIcNWcOSBMqnMeKDw2eBx5Oo9j
MXty5J4F14asaUMNQMChgEH7UBd2TMLw4VopxBWZSRlsINAG20F4AD3MNauYAM07e/DfHbkYrdDD
pV1gkPZXnYQ/qU0Dnb+uVOZwYFSxNUljvzwSxtjuiQ2xjrwyQRFO45jSenTC4dHEVvu+w8XSJ/TY
ZWa50wCMyQj7WNLtyp4lNWzMhfKd7Gt3zbvy+uTeFEYIrIYgvez/yfPo24YpnE6K1TRRb1aLkZZt
1VPR4MF2QL4ipC8hxAX7m9u2XHCCHccbiOIis8sm493qnUGsQ67kxL8yA9uN5TO+X43f7ewbZhiP
WTBBxk9tSDIE5uJ4zP3Ugvv67KiP+XXd5kNE8DlghaBYfB5U5f5bYcKzOWH77R4iM3sX3GvcfIEb
YVLbp5n1spvsrzKEvbjHTlOg7+d3T7MOBa//sqe5vldL80b7D++gG/rvyMeDAH3u3rH5+gKu+V6x
brbkzleCYETNEp3q88xZWecoOi2Vg2IRTpZWIQHtMH2P9tFkf9288vuFfTasjz+4ryxViXj1S1BT
bpHaHrcqm/P6ovNlBjSDnTKnQd3hmy4IqapEmJEtZLV1L0n7dFIzVEd0a0cOdbwPwyNY/EelxGi2
GAfHXGVxXRsgUX8rOizQWuulHXJVLDH3UsOCo/2cStnK0fboQL8KavRFQ3c8//v5SYUUz4Ch4LmB
pBmR5uLOxybiBLR9k9mHpMx3TnCMJsqAWqncgWqg+9oh2b/FiXXANC61LRfam8hD5RfdI6HJlvSl
i13HX7kdHdDY/bSRj/rRcgR1lu9NqG8Vy3zbmqgc2stxpCMQLyH8MHD0Sp4w2KCXJADRfh9cfcoj
0yRhkzLhffxFxmZ+MdZdtMz9fae+PTTD+9EN/nAuxBEclLpkEkMNk7o7FzoiRC38yc2qeMJe+izL
PUjJ2MNHjqsA+AiyYJojzh/bi0r7y1jSQEqul6iUXdPslNtIVAP8tuSE4K/9bK7vmKIzsLBmepCj
ZkKDPUhhbeVfOpMA1LV7xwalgXlrOIHyCMJttmhK1/IB6rpwsQyRIXqKve8npVqVYZ8v3BluDoDK
m7LzFTcpzWAWzBXoc7fEm8z4M77eIJjlG4AXGtbFrrOmVhH/q9iCJ3ejjffvOAKgh9ua4I+pxFpT
m45IpPFCdQWHKlgxfjsKzboWJTX5xP1k9vIXdqqoYRxkAtoLk5lZJUuICBBHVYKrcR+cQxkq0Ksy
hS6QaTE1CeGcN8PH6s1uC7CTkK5Qt0AKFy90SMYILB8OtpajOUSLia/PRDvtfewBxXyfz/iUH0df
4+32Ai3x8mQ/JDVVaxNbnezAFmxdUnjY/n267JhNF3tm6bx+Tf5rxzUmJUOD7lnjah6QkLv8svog
QUqMiRswqwsAeOkvWzvFjD0nOTofNdVG+s5Hm4tK7iKzn6aS56g7e6IHxpzGG/FZ7HoBywZkfDRL
H2qI8v+Z42zpNj8VHROXC51qojiZmtcAt6CIT0bJifPlM5nAi1LxdyLuZxavCWP9wP/GsBaKJPbR
BOcYxzCdA9HZLvwfYnYwINQAcDxf9BvxrKt6B7zEFlXoCP1bfgVcj2AfLTFluj0TZlJirISuhn1n
P7TlABqhPe3tJQqJPYEFhiFalwG40TX+eCaVrhK74bC7fQ3uaOWaorLsjzQ9fgFbbwwyd68d694F
vDGGqI2gem+mTvfpmGULYpry51//17O6VBX1CpTqm+diVFskaGwYqwxfSwyeoNs0NHncY0ZjMdMK
bfrAD2JnZ31tScTVYF6YVnSjy/p2gGiHR2b5nxUS2Lav4SjzoK4jvzVFICE6UMrDygIBGZIn6PBr
yBtITb9UzsT6QilR7058w6jL/U5l0UKNG+7ROE9CAiUc/P2aF1TyP39DlmyCR9k2rJRSu4vwpog9
hlpUZCa91yVqPj8qjcmzUE5VyWDl9PMB1MD6yTYvD+UULCRFxY2OT2cYeans6lr3vKMQQ1NPlXx+
x/VMojZp1+ShaSpV9fftSaX5E6hxQsxGcjcAkIF7d19kNHhVNgaFIZipLecipVaAqVitTANEO3J8
kulZlYwd0WGoxRzjXepzEXx/wlVWo1Li8k3xwZSnRZX0PvCDdALOiHyRug3N3rtXXGimynb+QgfS
ttn66jWbuI4gRwZUCNgD8CYMhTgWkNAJsoaKgHdsZa0xicMxhqm3flWqFe+9/VHETzvTSy+DhN3F
NkL7pYKfk2z7SM2D+sdN1nLDRCNui7hSuW7nlPJyUXtGADIsE6Cbo5TkE+U9/vt1poEM1o4Iej0n
rlHvXRh13lcEVwpLS62gXqGgCPJLOsxPhYcwVC+EfCUxsUvHCaEwPOV4L5zWvH4y19mVdDRoOpdQ
0e5CbkXm+933X2KogjEpEABlpEcSkgBJ7R1pj2iiis/wf/Brb/NjBpb2kt4LY/Pbcm3mxRS2CvAQ
DIX+6Jy5k5opU9JokAGMekVNgABrD7o9K1P7FYHyQjvbPNjKMnEDozQDfgmWft36g4kaHUzjH5CV
7f5VjpwiaAolf6Am6tjjf93g7R3BUr8enbPvi4rW2U+VAPjJvDwrBd1ZRtmkKo8NV4KmQLi10bKd
EVrR9WSF9aZdQEv6yL7cUdSRLYSxh93hVoIWEv2w26OGLvC7tPXxtj2Xxfd+7RoTO28Ooa7Sy7pn
kFGYrhfrwaM07r6YdeYE6q3NtL2mGFyjRb4mSKB2sZbRBBZPadKNsV3udkewtOqK112C9iUl1YMJ
wszepCzXy89zO+18t7G/HlYMVA/Awe7psc+yakFvuD/FzYOoL2SZQ9RKf4eEPKS2boivDAwIPb4g
q1miBip+TyKDN2EsHz5bLdYcwbJCS8eQ4fOjeTg4xu2uwgyeoISJ5FCIBlaXSbnNN17tF0NNNC3O
OEESFmcuSrG9LUKPjWgKWqX3hgfW8mqI2ozkf1nsBnDmmQRTVBUOr+rhcg1a4pecoORp5bs0oKn3
EtcIVYTetrM6R5lkpnDSoZz4YpAxih7JmUxsgu6ia2HnHtWpgyRShUwwRFrDws91XIURIFVpODbL
gwpVS0okehJFk36jnoWn2xPbuFUBLwFA+oECS6/wXi3xkELUnVWOjfVs92DyHIFSLKtafotUZDR3
fwna8lHrZFHPVQQ5TBF/hrUn0m2eztZ9P2AoCx6mHRg8IW6s9nBG3SzYcqsRGcTd3VfVCbCgPAhM
mm8ocndQSHO1hQ1BYsj/d6c7XLvJHCJgo9oN8U/nXXuSFpT56zTaG7JV9dmmEcdI04xCMvrqYzmN
0zTt10s8FjcXaVrBZIUznLqHGTEj22LtRRQKXQr3nRN1Fbrc1UpgyfjptsXvWH8v7PeRToxVVY6d
Us/DDJdjV81rIp4cFr4q8s/2LHTVDn//Jfb/EtMSzGDuWVxn6KU46o61nE73I/HBTT5rriHsPsse
Uuv/7RlOBEer2mqVhJ1WJFR6TlYDWIHXTXbZOk80YNBS+tAlZzsrK4z4Y5mL/IRItf0UjZ18zm3k
0yy3+NpyqC/G8I8i5V+oQxvH6KGoXmOzLdlYWQ2ogrMED2LDO9121JCKDnX+xdB35WTh8ugypfoj
QDuQZdFuvoM9oyrCUw5EDubrOMX7f2Ngz2+8ZSRWU5kpwKXUMtAmcLssUCKZXj/7zrtxa20xrWSb
+o8US6h+phl4MSSv+FEYT5DcGeEJhaM5uhlgkJ31FjGYH2WhtlpK8Q3f5AYYI0cjPEflIDgpiUzc
NQOfQ1+LyzBAiRMqkmkc3o6wSjBgm20HRrTOSLWH1Bt2lSWsFiyMfzhOpj2JF2d6DQZMGNpwwVUm
9Xo9Hf8lZR+VR5pC7n4BHDalZVi8qchdZcMhQyh3968UqpTGOZfFsDuPgDh+GgwastzII/6nCYCv
w0fngQkz9SHkSY25WMJthPoFRGEo8hwEsQcDMf55QYVndee37JTS7spISJ3lVnU0ia5qpoes1K95
ggjL9RgxfS79oFVPK27+pv4OdjqGpymDrhObiG3Jpys3CZFi31TRaSRt1+VIK7VO9LVjwEUXUrPB
q8QdyNp6NWNIjMvFOGqyzTfJdve3c44PxIr5Qod0MwJGobIyyoJIDgZrjAHFWf5dFUqIYfhZgcmF
Bidt2bVPRmWX2FFMe75eqYlk0/498dYfA5mYy1fhg3JxMvJFl2Pf6SY1+fxMMOteLQ5ohHJgpB0j
d7iPnW17pA/WfGF7/pPYeReeqa9DlIEKprymubqcz0NsCR2e9CJyACEyeJM34ljiv0nSgyI6Csyw
VOd4FdeucGG0k9sVBs5f2N+hAGRK+Wy0ZmJJ6XtU49jo/x5SUXldF5gReQ6q368dReQUC/2Vkqan
4bgC1ghQ9V0EhBkFONwP15RUqhkv1WEvfd0yJK91/OSkIDY5Kx/wz4sPRy/NJTInbf0w/5B81+xK
iPdJRR2MYRtZ2vXg6m16EahAlnIPFO0zkbYoozG1ygS7d4SqYC76LFd7CaR7YWG4CSG5y5awqPP3
x8mS/SFbWufQ/eZZJsblxBuZ1FUU0M7UN/JH4JdcLWn5EVLNpReDFYyd0RjqESvoLRyU3zxEGWUN
1muxYNFga7a43UK5t4zX5/piqz5Lcx5+ZFJKOGdgVSjDYim5afrp4pWi/iQJs9KGMKVFsYkqX99H
bRPen6L1hd4TAqqtk6eFMfyazS1fd7vuPUR6uiX+hCTd0bQzvP3hD8o8tz+C7djE7dSHhArFibnI
zcSQijGIzDsfi7wFuaRHb0cNa1bp0fTLmsNfnXG71j9AIME1yCDgwFxs6I9Q7IBhCW0fyDF6Mc7U
xcw0Gm66yRXnf9XhnTZXqjvENAgpCIySlGDjF/oHimMObS6unFcD5qk+L6nrqmAVGmX4d3U16bKu
7NcV2HBArN6/5jUdYOCMvuPUET6lhtPFqW2ua+2gmwMXhHaDwnGjj6ZJmOU30CaTE9EGt6/qN9im
jXfoVieKntnMNVqXYzyWBIN9/7DMbRVcHeCjFghfQt+8nJolb0cn6q+ltXIYNBlYScDopqvGs7LT
dZF8tQmn6IZx8V5DlD5MH3o7x1btSnr43j6If6p8rNzgGhIrRD3P2PQ/VWMJCl5Cp+F1lsla+M00
gGdAK/DsKcCLEUlnHBhus+qDUABWOBzd/IFuDE4yn+pKXlo5+NgbhZQBAsR0rhXaZqeFUtCETb7o
aWF2YC7hjYF9WxniooD1TSbPQSRKOMcJ8atOSZfvsvoJ1R6hHs0KwQxP9zdYt26E9MeHelmpU6/E
fjcfVEM3bgEdppvYXxGyoJdsRwcRT69OxYh97BvP6XC9du706hlONIwgSyCQGBV3jxwoPjgSCcsh
IklpKZ+/fvDfyS1TcuA//S5Nfngdx7lsL3uO8yIWMLs2Fvngyl03s8wz5BOQqL47l9o1SQuLJe3j
nUgZHGHuPwZ/sJsBWJNFw51uXivqo+f3hPK80Qy1I0gW+aZe2fS435jUlJbZWc6KJQYm3+3nEmYz
CBnZ+bOQ2BHLiKfd06qm71UhZeSgcahMOy2qFI9Wh0R3W7xhE5zwRizM1o6e+8piRTB51beJN9Sd
b1VLfCLbaC5mknYr3InIZSKiHMAYocNeVIz+NnDh1ErdB3UHOXms3kHFl9bEPxhEfUO+QzEUgMPZ
JdboMif0sm7O1q8erkgef8VgvpzAcUKetrTDqfUgogJfhV2iQL45ROT3vTOPuEB+AHEypKzLrd1F
Am+hhln4n+isu92ID1HK/Tzm6kSqoC47VL2vNsdieMHO8of9AZ0rfaGfg1JWmQ+cFRryt7ekmbgq
Rj3PHylb9F3Hrt5Vsa0lQD5rri3idleINXWDaWT3tzEK3dnmW/NOjBVBGfzBjZhspuOJH2EEKR4o
sH6H4Bde7rvE9eMxVS35RDeLh6GjN4dxKmBD+ZqcoWm8YM5Wc6+wa7WzRYSkcwaOUsmhKJJ9QYYE
+L+gs3JPra/2qy7xlh34nW3YEaCpJYIDOEdJhh9GcWLHCLsVnpbz8+eXlDt2Xtgz53WnadrB9nXE
K7QxwccbIUDv8hIJGSFtfo+/lAdGKScQQAq+vkDSSTd5c678vUBn6UuEZXNCn/HO0Qzpqnmp5fKl
sdL6jtgowVcnF/gLh96lV6ZR4Tj95da9zMBdzr8jEwv/Y4IJj+Z7Fzyd3rKqAfwl+LMKup3+dJmU
Hz8SNLtUNM3jYYHrIlfIRjVp++bp1s6Dlq28u6tsG0FDHR0iY3vZU+5aGEoCr/xHvmYkRLqxgL/t
7KIO5qwullQxoqmaaGy6aF/xk/OaZctDZ77uk1DioYUvNp/r52CiK0VUqp0OYz/aMlisuMWWiW/d
hgTVdSyQi21h7MY//66zamh2BF9KvuyZpst5NpXT4aQANAKMWiA1EdaUCQEAzWU5nRoRa3/s5DsL
mCt1k77uL3pAqCdwKItSNqHdqqsYRf3OtNpfCfq+iF3ZN7+kuaQjf6YMjK+jbiBWFZPK+AuMGzVP
DKdvdi/dLIV7u/38ochaN7SvmMPLr232o1BoRnacD45Z7Sk3o0SHI0XrE366HKa82xVLfZybKTiM
54lFppu592UCczLwcHoGkmb8Noy9KJmCxP7WzmDbQUNiA/HETn3dCXcYl7vjs7+3++3OSUA7Qshq
oR0l69aK8/T+uTPFLTsZMtALBkOgyQZMrhTkn8YVM+MDJAnKqk5foiDt2h61+AldC5dGyadWnsEf
uIGjhWzzj4SVPBJLKINSwwVvLPTGZpONjioE5KdTJnjJC5fmVajvtBXvFzHW11CGXJW1FNbxfsgf
s8p4ExVq8ccdSF5CQmIdiT8yxD/uWJXmAgqhcniBLAa0Skj2fqEz6okf8b4pjWxtRVnu7/nvXOGR
zLFpgIm5WH9UJvDm/dHGeSuIODRhtUckr0WYhyW5k0dPS1fNwkTGOkOsVCsEDcmiHdDm8KHeSSlj
xhj//7KwNxEp0c6C3zPPs//FgTIDnznd88C1kkQOCu1TYM57xggAgb1mx4/pAxKH12yYDB1E0KOo
tfNOj6aWk1CXL36umTUfP/Jrt8Wj244bExV05f3yDofqaPgnvhXvBzFPw+IYZz7eF+TBcn8PsefZ
WtQORcVF9z9znvK41Clk8psH4mX4PJElPyNzYsCmy4hPgydSyspG5tI5uWSSN3uSe9VOqWR6P7hx
IfIUXYDmRpODKZeRAlwtcKVABL7i7NFKlsReS9n7J8xLX2mmDJ58W8vLkMKDhIpDsxE3I9r/Rhqg
Xi/7exuynZjifsF/x2C6IRIarUa//RYPTL6yKyp/NSAX9mWTBh2NFcdux6ZpUfPN5sojBGh7HS54
EXVjVvQ23FPUeeve3IBFtdvDm8cOtre6I7xY+YToS18E1gWj4EAkU2IwhLeuAvMQkThMFxykITXa
NrqJKcHXxCaZwgZZPwDev+ZeUFdVmg46TxqPKOy0ht1KH4Uk8Wyvl9sC+7EfA7MIYM3ef+t68FBJ
l8BQukuo0+G2haitke8kAPI7ID9cmfJGWIpvZCy8IB3OVuEIGu3yuFWMCDjQSy3/PZy2X7fdhRzb
4NLA1HMhyoHSawfhfk/fLlEJh9DGxvnJWghKab68ChB3O4NhwF627qUccxuaMlOPrFnNsEE/vosm
zlSPnogI1//qUKiMgvFx67QH4yUcGRokH1rPXrlQ7eb1iq2J8JFLOfe47f+rALxUxfiB3J9U3RiH
DOvNvdfCSAt5QXQMyj/ESByyMPnXNLmSdBcihfLibL9Nw/drLN3umxGHDAiocuptqRVuhVvnvzfb
49TR5cG+UbhDzBu9F4maKi+NfZFptKqlKDtuIohLoUK5s8x1aqun9lwlH1DhVgJ+wLmR3JjrcRlo
OaIuwwfroDqiK45tYiT1hBeYkH1qLcX8x2FeGYkq5vJLrjP87du/Kr7TS4GuAYGTKosdMPSwMARM
T2btHWtOGvxthHoJc4Lym/EWbkWVR2dOF0xfPSqLj5RSnO2/dvcv8OQnYRvKWjH/AmGphKs1zwFJ
+bOlTEyxY3sDgrdDnNKCWXak8dbKl9gucATWcGuWiJUfELkO1IJzJv37GWvf+kUAz2DDOI1BhH/A
HUx7XD7CnHgRd6mr5tNeNQW3u1cZxH5LVpWajdphrBJYL3vQ6wBikS58uMCBPI18wMKn4YnHrsqi
d7MRaHUSZi0EZx+opVav24ehRFGqveGL4zBw7tv4IYwp/1Su3NgD43fGy8tyGku5/vNzzcFf6rwg
NOxcq9/h69rPfhO1V2lpHjQjjMwSg76GvcTWJ4WbCTr6Dyi0pJJjUS4O7L+D2GRQXJfAmdlswxTW
Kzga60BxkTECWDppECZYdFXBEthhU5ZSmoeIj+nYFPkyqDBJECKx5n0nrVxlJSsfK0mp5tegbs/U
abfMzsByQbHNUEe77FG9d4BjvnXZN8fKGMg4YPAcDdDWS7ifCyOAyVH6Uk7Angh3jhjwYnngAEw0
t/hwUyMAvVOgSIX020OjiwoRetZQOMLDlbSv3SbaGgjpyiy+pMjYW8WOf8ELpNgyOza4+wPbOSv5
gneQ4eIyvH2EKItBcFWa08zcxl4bdg7PURMMoPewlWbUwln6IhxfzIxCA8vOuCxPmoWpSHhcvqq6
fCu2o79LfPUczZYMZrsFlx9AAASZnZPnnwXsYIrrKmoHHzFTuMYJxxOKc4kZRN3OyS6hKbPV11hl
IGsqApg7kl36pw/1B5p1rocd55WA8CVfzXCbhCLpbLascrENdTfi4zZbVLWLIc4NhvwUxXvxNp5O
A04TZ84PcPoVxnsJQ3+0TBp5fZf4c8mNaRA6ooPoP3kHAASBRmN2pk7KACzA8PvBidWS/59vHMhA
+4PafdD5583oMKETnkavNqiN1C5XZ4yY0XoRWHY4GgV8S1FkiAIppHTiH/0M7C0H33VqvV9IBJOq
vHzPlKalPDhLGGZ2eS39G5yWvBEamK2nhKYWuBR6YIzv09mf10djsoUTp5vYju/JdYcvu+ACypvq
pBRA/2pPKlShDtM/vuYfWV8rlwFeuGV0qnzID2mGNKmhrR0G6Av2orzRGBqGGs6KAb5dBgxhF9VJ
+ngZb3mGypkF2oEsryyZOpC7b+XWZ1DeniLVkJpKNFIT7vdLiRqYR2F5caAEo6B1DLKdaSs3ztX2
H8/Dkn4ZiJedn6EmO9zBhC1CYWJcozdZzeT98XvqALjrx3b83MM4Ir6ge9u99gghE3XE3b55gM4i
/Ijw+TJ40E/JcYnREI0JY3AWe0w1aNo0+Ckdd2uG3w5r0R2BEroCa7YKQ7SWjXgmg0d7YkeQEaoe
cxuIbMGJTiQ516Dm3N5nCP2Q3czUe6PfSAX1faNyS9VGwe1Sz45PjyCR9opNTFzWRDOX7q6n6hs0
cYoUAeIOjvWrcMst/wmj4vv8o7VMGIJBCo/YPbA6/hpnVFK00jpJueZ7SMvWlcHR0JvEq4q46rLW
fO40H8C3AccYHTBhkocTIFCD/LHM73PS8psMg1+zFPlFxWO07a85sfRq+GWr7Yi04tas0+324dkT
gR8Wn/gquFDckDywC15yHvNVSnrv/EvMsBzPAu0zGsGkVdo5VHWkPB5z1ErREwSx4uQMAA1gIPAg
t/ACxxhC/wLNe9kZ5iN0emVp66xvvV7PSb92jNwLStA9Mqbs7vc3ZkERcWwO8td+rq26kwj0z4be
eBt8KzKaIH+4HWzWt316Stt0fXyPbW1uTFV2sc4yXoKvG6DlkMxXzs/m0cyDtuFYUl3S5tzCxIRp
KE6Qh7b/dSPXNXK4iex1ttUMqwPY/7h/WNg9C3ZP6DjtpL8+eG4u0EGlMUiYdf6R1/t7EqEE4NK2
1Qzma2HxAzil7GrnUfynfdnDZM5TuDZYafHrBTLxgwmIgieWNv3c3yfo0zJr2N2RIwlJ5yKb0hd5
1wRFybfHqsbL01V2hOl3P/xdsPQ3j3spUwsFYS92xDuJBdwZmAR+wmBbzFss174KcMyc9m1ADacn
HkpnaUTgIN490uUrzYKpddh3E1UzJP94QIiyzI9fKSdgwLod6gLXmLnNHTp1tSEecjOoMIEapO7J
8zClL+7532D3xzPYLwB7nxq8ASzqx7X7Wkdf9sMNlhmhLNoEyuvyjWvDceT6IEG5/DOL6/YVetMm
6jgulfEnUc3ymmRuKJ8+acIFItmKwMaIJW6ZoLb+s1hy3UFtyCgEuDPnXQdIz41+KtgCosyMWiNB
JLjeP64jPqExdZFTCNFCEnnwDh3Ha/aE1XzS6jWMTPaIMK14nMvoMnoOKk4WgqReTlPap63aC0pQ
ttINxgzcPo8DYH+lXiby1VVP3snyvd161rnUV7M8KZqPMHxgNB7D/j3JizAlv1FEszYCgVaYx89r
lkXThPwRx9OwfgMa0lwM89tKEP+wNBNjyFNzwmIuJ49KumxpK3uSAHw4sFT0WWl12iJt+OG+rxzF
ROI8XP3c5ZJjmJnSmSzHIeFv1NefDY6HhsIEaX3PBzQKj2I6mrlpqtRTkZ65sj7WUvBtYc8UEW3e
lETz7k/o40qqiCRk3QZqXL/ZvCYQKYyKu4qnjF0gd2yNjufecVN7kKxkUM6mdHGcOcwU1FdW2csl
5y1mIGqi90m8I5AtUVrY58b78TGmpAuIlsMvZQnD99Qrte4n0ru2/N1SIc56u8Z0692Yg+6lcowa
MdFRX3pcVr/dMUX7ZvcdwW0mjYGaObWmtKFPEMJP8UuKjQyLc8oN29MMNiyIU28iV/YizZTKk4mt
Ai24Zi7r13sqmlzWUUlRRMim/Mq4W/bHDW9VAcF+WJmelhP3arFGR5PgAfgAu9nELyIfr6McfcU6
a7O0MyNGzUiKj7pWjaYFw/e6w8XvsArxtnH0/5SPnRO6z8qp3BUJU1sLYTT7fuFQPUQdRWrAfEud
pCiuXmnZu3OfjM1avNwbGumTRXvFXF9UvBVDIYf/O4CrvebII1eaAwEzqGM6F0pJYmLVVaHJNcDL
zVN+Qb4ac/AfIskEDzdpovQbXj91RGoicDVRX5lqFOWFBVi0CW6kDxS2klSM9FJSlRWfQ/qwC0b0
huRIhkPhHvr17dUmCv/wwTzuzaod019ahsjGFD62Jw7BuSqiaBxOrcvSZKxrvHT2xhJztfZVSdAM
VsERJv+R6FIX/meJ2gzHctY7ToGFCAqJ/9gDqlGJY6EEdvdkmE/akHTbJ6pJ+aqmmPKDwSYIgtBn
cCOYdwIeRUDlVqXNvzRRxbE3Bf9TZXn1NTjku5WE/uNF9d5/rng2AIqrZR2zILTYl9GQI4dOhbPC
ZoKXr2wULSI7lRriV4fKBqNM+lbIT1Jlkk2PaGTCOKu4xbmJPFTTzlVJ7FesA9VmmNVQsI91lqeI
MGJvcRho4kvZjRY6MYDgh/3m1s+7IopUJlEB6nsqU+/cyVT24zQoJcHEWNC+VFXB3WUUrSJb7uGW
06IYmNbZxBCq91GoooA6ZiP8B4rrcUwlM/UcJWs52jLlu8aIsTt4wE4K8BHB8r24AG8hDjDhuSxA
GXpmijhVRMNy1NUo8QcUzSZqirpVUeyD10lkhGQP4qJ1QV7iJ7PP66UH+2rW9MwnkXKHkb/1lsaE
n9W/nsOZMPBT1Y6sMDwHeccyyR1BG7tlB/6sLEWKl8AIsuy22XvmIl6hCyZ3npBATGkpmxyM3JxH
c5E8pu+2tPAKoCLqI9RzQL7BXbH1/5fjAa7qMSRdroQYuFasSmx9zawDiuWEHRIUOnrkbCKlxFou
/Z9jCSEHw7dCfdpgwcdC0jC6RU9MpwvfvotboRI+CzXvyxhcZjI8WzDQ0CX+7RhXjmxB3NTf67QR
1ucntA6P8tBNvFmNOxszp1ncoaa287/S6LRBSmt/vn8EuNvfsqrfmAVBOVLvCLYTviYXfVBqB9P9
6IE+eyeE0D0UlNkrDDjXkCwOuCHjlzSrIrEQiNIfWEPBqhRMRnZOqtp1COYCOrGGR2qvI9gRiUx+
Mi7koSh0z1NcPo24n14xoquHFdPsi2Ws/TtySqmkk9dCOAl2CYfk5vQfRqxpui+bwvSikuy8WmSs
D08xaPVsObStjINXsB5iWp0Ih1WlW9HPL+aGMM6CIh6/NH3D003p8L/V+Muj0uTO1hMuc9kVSDIT
Tk5QxwKh7iF9vcR05kvmcLRaiHGuEKeosWa+z6IsMzye8+bp3X2TVnCfCVxi3wongNcBO04uYi0D
EGKon4mW4Ojwg7xROOQMSsqAq2l12/uQwocSjI6LulV9IJXklaKXDPy1akzDrzRmM9PXBuWeJzUS
+XHGJk9JwAPC4TpBsj9961cdpUvnWVt6Mta7TkjkN9UwgbFJprwI4kXpRA0fWM6Jn/kdfvri0w9g
tSXb5nUIucGwAsF+7x0TJ+mKbR03iQRxSr2kw96+klsfACsZyVZ0STqI3p7R61EkT580KmJeoig8
uWKzoixn0V56JtMa2tTSJEK31V3qQ4acpg/Ga3Y1B7uQ2oToiPyQ1pMH+m3gMLVvclrymCNVmmsd
s/UrfvTZaBMce2GKa7pwCxLCzXd1TMvPxeHVANCM684wi9NTG+blgNg6SkmFn29IXf1dLBi7HeLt
fuS03SncLiYQkAXQp7XLl3BdoUXq514EMSXs+rNktP2cC2i+4MaEwfClMYBu4VzO96plcaTAbU8w
TtiX3P6ae9jdrZQ1M7xTVAXX8Vyrt84loPfJhUcJ6Tt+cfkBYzrXzhMwc0vs/3Czjolgz08/UAhY
sqJ8c7bSvUxZgoMilOQVvwEyP+Qkh6IMJWYbv7amaNLk8f6L8g77oVH6u/KcCkl4VlK+JGg8bznu
jQr4kTpVOZhmZ2PJsvW54CF6leFaEOELFxC2fk4Le8N0JMgyamyEbW5xDisifNGH381lxNBaUH77
ZtwRoW0pQBoQ/sWnst2BIMN5Np6DlvZvxZpb172tJyvckq41eJNpXrP3hAiXNQyslE6pUmTPtCrJ
GxqJW+ETDwp1QuvwKLG59b159aqEEFk6jO4LVChM1175a3tRQB3hzgAa/OVp8uNwQrsdHN1orFet
z7JSRyuTEa9ERnbINEAp7aspE5KJJoI0MnIYMLwe4iFTWbbHaKpalwtcvacKvDR2GtvuZrDzSwCb
TKo1shC5epUwJRfyM5k7gGg+e8Gmos662UFUrJEGHGKKaOGj6TYIRsBKQRIw7T6SCd542Hr5ORXK
EI2kTLSSYsNfBCIblXa62djJT4HjgAdoaSk/rGFdj0LzQl5OKFsiVh0py13q+PdmLtcpvbmhs7J6
HZry+z7rN3BoKL4nhgT91HmPkGZghJzv+oOBx+kovG4JtZC9C1DhdzDt2E52AfDnp1eRbCenaWYN
U4cwCqzCtdDwbKBHiH5CPI/kAvgthIYUBNq/NQSfSwvCxB7wNMvF4cLlw6u3SSPcsdS8xzqTSHxR
sVZuZ5pl1dmkMofyZOXjwZD4IEiTCn3NHbC8SdE5rAmCamcoYQXBzksda9aLg3jICzCWoNAcrckY
jexEs0Dnm/TPTelpVkznm848aM4sKJa4NJfIvwT5dvWdelrH+G64tjLWsuoOxH0keWSKFVCNFTUc
9D+vzaLiYInm/TqW+dOngNaJTHjNlvf8E6BgNDY7+EQB6qgRDaNphbJQiCZyxpNdpTsmCVmM7qFl
3bf5te76lTz5m5D+06ZyjC/xwwhtrumzLmk5NUqopK13RCb/ugYdNi4beMwWcuNj/jhB0eqhkqwN
ABXsIGHiYDQ3wx06QJ6myDyFdLgMeBxspKS1oWZe+SWzSwNCpy8xXm4RUL51gu0m8HgivWXunJhL
pWfzGo70vnzQpBDoFEtVO48YRyQv74DMpGoT2Q93pLW8B44kALL4XxYc7XSZNC77K0wNFwf+vb0h
Fpx4RpYEeB3YhF3Vhj1hvjIq7iEpVDBEM2ujYe9d2ItsOrkqNrSroN0BSBq82wmYhSIsiqWvkP5q
2lU7kBa0gUmVWQxKSsyrlLniZDJXf4HLOz8wbeHTJmukzIsabuxWT9gBjOzBMDRzN8rbcZlJFC0R
UU23vT7d8E0X8JJYMy0I1mYQu3QmO8cwpcieNiY+3gFGBQNReK3ozcZShkoxMHRWuq4Ff7zI7l0y
+fpL6bpUQvP8KwzpOMgKwLvvNn9sEPmBTBixfQjRcW8VZLgMPA4OI0f6pcrbLzIMnsP8iury4aPg
CrsVFTYXODSD8lklbzM5b8y5DOuVtwP/rxI+kkAaABO6xC6+5ZR66gUYZCgeqOuYwunJdsiLLh50
TzwGp1jX1kAgbof+h5H27FZtqKHU8JZZTafH+6ahc6GEmJxMzWsScgY+JqrkTfeW+FhihIhTmwjr
RwEjnYWW/MYIhkORIb35OiR+mtfBYrGJX8RcMIEa8dMe+XIfTSTJcknf9bIk561mjr+Ir4Ayg07O
Au03Hph2369D/PoirNx0N2qUo5xcWxQOqkPyl8tdWN707zXOGSc/a0YAzJXjEX5/j0I/QQmjhMkL
ecnQFICbA+i0O7fPi+bvir3cXHBT7TtqMEXU+0umDbYllIjl1hux4xVlKEIlUKWjcH6PLo/eFafh
dRxZemOQtsgBfNHND+Or/z1t//8hSp/jHw8KH5h3EehziGqnOUSKFc1DSYpt8Iji68xQh3h2OiWf
zqw86I+JutMx5NNb6gJrGurk9ZjC0xwno1imTxeOSxe/o6/X5ZrHD7/AgdJz+UR7b/MGpZwUJLQj
mq73UKYdTqSfVVtnJefrC+0NDx7svKCVoaVpbAeKrhVLghQrbOy4APXIRsyOflU7T0YXlyl9jigI
bi8LOiRe8KNxvCAmRVMdMgQV1sBV3VuWGoDwbc7ld0WIs2//vd9MpSQ5n/somaRZFIJTMRiYl8xn
JJdo+9hHuEyjFexVTyTcyQBeebA2QAy2TAQgP5YA/Z3QUEoQFyW49SFREs4wa6+n8XYIWm7wPmSX
JQGIp2+0XESXOLoYzdMI0a+BsE3vJ+IxDq5t8tdnqgOTmmhH6qAJua5rGUFsDMqqJpSt7XgtdNlb
u7cUGuckGXuH1g88D7Krfj0/B95dnTn66U2/IqEkdpGLXJtqDgH2xVkgLf6+5UqfPf8xQo84m2qA
UGkXmK8n9m1ti8LUtaQi7q579+F8La7/O3NRch6B/NNEZKIwlPnpM8Yz0K2Yq0yNHvDe4BWck4ZT
V/CHbVIsWQGtojYUQbQ3pBEPUdFiKI+w3mf1GsArGPaswWp2W7zQFbQB+In1c8K2qWXgfdSwBezr
BThGQ0E71Vz+50tCDuh7esqJq1thNG+KUKLiN0XZ3DTKc9mc2KLbNb3wDJ4oqkqtmu7k5UgbMflP
uzdVdEyfMlKb0CDXJ/3MoRhjtjKpZbkJM96ZKCyXhGZGkO6jgyi8Sf4nl6IkEAGhX52qE4usVvjx
QU2fgJRcgxUM88kddoxCM+Sxx4/BnrDI8R+qC8T7V+r+qnQMFYabWPbiMNpPy5hfD9j7emYQ2di3
Y8ZxUazSKB7vI+quhD5sTsjLlgjw4Ve8RG4AESbzg57izfnKOz/Ru9DodDWBoidGwFrAs+L84Ufb
/F+mZN9WeuKEa/B6wtQxeXGbztVVU5fR2V03LcZDrnaA6JVLkK1cUh7oP1M0zT7Fa8Bd+Y+GTRnm
S8cl+9jnu3eLp5JE37hiDNSCAFewbFP/DrsrLiU4lJ/9jlr/Fpyp4wTSAM5N1QVlWLMk7lKITjho
CR2JvjRu9X7tm5gZVESfrHuKdYNG+NJb7F04iURLinPV5cfLzYHp1w/FY+ol7my1LhvrN3sWsXRv
RAWhOmxvAKkLmVWbleiVw6BuIRfe1+rI5Y46PvGiFJEEjmgAJL7DvPD2T9o6xVAYlz5PH0XK9HGQ
o/xDDtvCBnQ2fEL7FGronU97O/VYZbtb05jsAkFTnlUrLWzL3tkV6GgyvfwZsx4UYT9wQZvmBHPO
oInZLd7pQMARj8kc2iVJR1qBUr4jm9UcT2u5xVyckFJoRcpWJnFEbP6rw91FTARIMQUu31Gn/nGM
SUUnsOzhps7i3o20xk7y/FY7xdam+4/INiP5Fy97yOMZGrbat5dqnhvhj+if8Qn5Zl2OKjDMqXqf
8R+B2VtkDiKvKNV8AZgiSJLMSko4xmwObuRlDQwV9UG0D4q9lor4GDK486escIx7Gznmpfni8NtO
s1Vbg8XY4uZ1lV1mHNs6L66MyB+nJXe4I/K+yEiaD6fMsDvkDJ0UJshrnWsBu/TBIxVvxBUPQVR5
qcsOVJkRAnXHBot9bH1sv8hTSGVd+bd/+GWdEtiU6YkefnW/IvMdA7o+7qwUcWZtcnamU6+1LJEb
dNdqeAqrer6t8pN6kqpm0XIzd/CAbv3Z5CmVyKyyLxR1tzcsmq3IxF8vzH9i+I/UvVr0a+ZSM/SU
gTm8a3BATXyoOtfmJ0dUIUGAUvOxDJWXeJor0atlCP/JsXXfDCBWJRnxmf+lAjrvdOjp+Z4cSl3D
qM97XqO+wXsdheWurtk+6X4B4SMZAhB5ZbAOEp/HYakl+SlzHuguFloemO7t4oRDnLxpB0sm71KD
whDfzIpWWYYHiu1APBO6far4tX8DvHsqwVs4PoZ1qSl6wAPdAH/n80B3FZ8yWScOJ19J3prgZX61
bIhrGoHzXrtlL8VUjWe5k/dbimIlqs3e2tkuCPlqVh7ClZXxTk19nLT14WLF7vsXIjKxyhX9RfL5
bXX03JO+D9pob4KX3+O3Y+ddwy+fCQCBG5OWJe1nPfM7mC626e6e2824G3MDb8IC3HQDV/OejwzS
bvmJpbCPqwotsSibH0yzkuB0LbXXPF7Pdg7rZqA/+1nQswWiwqgf5lRanqNG/890zxWxqr0wqnyC
7bpeOxQTRmBYFFsVc5A8lL0qjnPg70m2S0g7Mrt1PT5EzLtAnJ0JqfSQlorfpYTHDkeohuuYjNm3
hMGrncMR5zuw3+JX01LWfRvRFDLWlW7v1aHMEEWi5eGQbNnMP1tP8p9s/uJ8/1R9K0SxdfSf4Pti
752+7nQGCjiMajQYNhE2whhWvCHUj0DpV1wZbQ/G2axsQRHJMV6cjBbCQkQ7z1QbFiAR1UcVU9Gx
11nozMi0D51G070r+HIcs/Egahdg0Z4YGnf9yxGbgBTJVMwmLvEZ+dbxgmrQc8S0YZsOh3QovIgN
M7qFOZw8lqtm4s8rZcxiNBMJeqhqD2Ngmeu3NhPxWMuXDXQ6ArJUbn50nnsJDAshVu+6j6cJEpom
AaSqKCGzVp3LWu4u85HUp0k7L0AJpp41ZP6BVsqLeNAgF7dkg9FTx+xSfr7I6in9vJ6hRi53mBqs
TRRvp4iTbd4tsEHph9ETUZK5si6mVG6KxAzn1YT/5WhsNO7kZDvY1ctzopf8cyQWe07sctK7YVKn
LXABIa75L91nTxF9s4zp2pM1NJFXSV0On0EHUmmIt+ggKS9QwR6EmC8NnzjDZiLexJmHDkyOOb6S
7fh1IPrMrh5AdnXZ3nBNP/AEgDC+OHoW0uj7rEZLp82ZslN8gfLLtIcEpap+5FduZYCGRB3SyqwK
ta9OpYBEHVmfOX4g/iWFFRJMJfVR5TeLSXaQHfdVasJiifFramR00Xmlw22rkt9jcl9RWy9AT0xv
0xvvxHz1kl16SjOHscnPekNzlEAiceBbqU7ez5rphHI/JnxveCsoWXQZNOyHWfKw9qnbGFr1/6sl
PzQdgQxzwiKusIFk+kjIy4bNd+/tZokPhfE2yPQHbLYIyttjtPLN2NxlZ7qBOxf88p6TDgSaZTHS
NHqwmdIKPraPmNhJ8t+FTDepO1i4ggwT6OHpOkCML18gq0RpJGTZYGYl9HBmYG4cCn/jcON3+/ql
c7sTdxRnpAqgTpf9SlC0QadOnYwWSqdCnc1NDt9hhZYWiKvfM3S7RRfQBqMihkac0lIfBOBj+IOb
uZvyWLexQQsp1BlQCZbwE4LS+9dDSkiFr7j7O7Gqadk3N12JIT+YGJt9N/u10B5uQnXSDNRKWWBj
fepbcOVOIPvn/0e2KsC0vB7HwB0/Kt/P8TmUaDKj1I5Jc712ZUAs+6UGe2+sbGoZ1PTnwrXuTP1F
o1iymYdvE4fnZr+OeOS/6jcYwSU+yKeccEMRD9D6inH21zLgYW/Lup+oj17tGpM38aNNxKmDlFV5
Kt/RIZMqvIEooJ0U2RBfj1ImD6Zk6OyBIjb39NppT+8UuC0Omr1tbG+WLXebc2YXQZght5cCA9j1
kkAB8EdnUx8lPYmSVIJxIzLfD19vGPZp5V/5Y51VXBUv8wfkCpZjegvIeVhex3M4q9IFem7n31x+
rIFTpWTXqk2mRkt2ARsoKEF5PypwlpGXUsfIfqiFfVgju73CXqtbsUWcm46D/KuqSZdQ7WehQ6DT
UPInqZlJmsdsxS2jk/yJ1wZWLdyKG3H57JJXF7GXTFtvLmkb/ZE8gJ5FP9lvQ26FfYyhSB/71L7x
MOFKbI8Qs0F/3QGm7IBGerit6/oqATXHqgv7R3pR5b/hYLCdTAjtSfAQycmnY+peY/EwJNZhoK0S
rIPN9Bc2egcc8EVjIWDTm9jzkIHLReEfNzfcNvKq/dOtZtRI7lPlQ5OcwfHpbqCusmvKY822iYmi
WzVyVfTLdbUZ7mTbSv7xdGZgMryI6cSWjqIcKBI5wTcqbUMlOa72SMFI3STrfkDQ7I93Xyjbwgeo
Plyq9Ow5q9rMDQfF19+BoXRU+fxVMi9AOB4CVEONVQ8D8a+9ZeN67ZWkTJFO8givk2FLvtSGINXv
exdQT36BSGKpJ2Ow/EREYlXqEfxKr0WodzjQLKTNScDZ+qfLDeJJCZohjpTptqXRuer61wTqOYTx
vDZCQbI3dX+JBCCsHPaXra3rf0fvbhaIm6IDcQpwBkWJNXd9QBVSMtZgz9EVn82+BYfVeYJk88b2
g8nSCg8YeVsbt2oLkj0dOftfYlJLIlWkSK2wgD9BGmiEN7PEjvKeAAZTkIMsTNwLGa0lMZtYJeJJ
BBQ5PcWhArqYoME/9U2dJAznNG5ikVQO1+0307/TFW4xm1jl9Gts0Gu+55RjCHHUQF7BVkQDpkGp
MKD+t76gzqPJL6OPoGz7TEbbOHko0dTbJTUYb6McPDThEHpmwf74UGcKoagcOoiCURxwDzYfUUML
KsZm/R+PPXz8N0gPbayYUSDNGgsFu52clDX+A0SjZyV+B3ontpEd6MKs8R8cSP9Ic9EyUH/vO1aS
lB+T9YKV4RVklFL2kXZzl9ay9B0xBcFI17v5S55ldYbzQnREltdMNFr4Um48WiFbXVIQ9iMEDvm+
YOpy+lU1hX2T0ZTyHOt5CHLwVwot+Op4tOFwLJGoMpuDB+Er1A5uRaHNxjZZk+LsfCQajUydFcS0
/p/RPERNNu8d2gjrFTVNAmxuT0GwQQO1/hapAByMc64gJGqi9mOzhDk8fUsSYDfgaXLrwUFHUbfE
xCUCPQQvgS/bpLpx51dtyUzY2fJ3ZuyhDDBXeuLvjH576u02K+UsheqsPVUj60tOp/cII6BkhUs9
IbFnpwZdlXeSuXj36461jkSBTVHwWo3NlUwhwaBBHt3nn1i80YQ5ZzOjOVYlmRTg/N+2QZQ5Ci7a
b8IoB6Kj0aOW4sopkU0lxyyrGVkHFWEuIYDFUspROQ/PZKMGUylgjD2nZT5/f8A6xdyjoDKnxvwy
YJT0wJBOa/g/qMM9O8ICukzdmA0ef6kYitIastVChB54RY9+2L9E+ORMNJcVDaSzNte8BtRPSbJR
rFwx1irZU5OfYVqZr1oiHSJUm4Kqz9T8iI1mreOu/U5THDaVNRkobEj0QG4e5n7/YIYUi6jbXdD1
0QLn1UeiI3Y6bns2zx2iY0S1s1mPtcLPCjZKH4M1Ylz1KfQ4kQmNaMUDx8LxmK/XNmflZO82f+Gf
rYBuJndLUcimiPzoUrWC+1gfZdC+5VsaqzVNnKI4tDmibF/pSIR3U4NUKj1RRPgCxi56VyiL992H
Y4W886sCYrF10wcMlDd35R9gI6w4vTD3iRFoTgGymcuogqaOoquLrwkHFY1XG8cSixUl9D2AVyXw
EfgYpCEBYgpn7z5kT9kSVU34XLIJNqSjv4zkyZFnxlVXCvE0B054m+PbvL2Lb0xLM+QBSAZqOrmm
/+2ChEfBrFDCfaKqXl3fkfuX0JpN+Yxf4+5ZMEV4Az8N1jQc5AzfBMNEzJvLC5mBoB780MVJPou9
VuRPtljZ2tBXe0QmkuL0vGRw/Jn6VCwtj8I0lMJ4v1OTl+ZfMZEhVq/cgktE1r3IknoUs+tGv4Gl
92aB1K6EiL+VsxxOQlsmOKQDRP6vMTBAw/i/bEZJA80mQ9ibOT+uS669/wy4BbDJuAtujTiS4CB2
4rpimwD8HV5OJ0Fp0iChtkLHvY7csw6mB12bwDXl4drxDi0vlpeIirabh7eoymx1hxP6pkstxukQ
+Omr/WgfTXx5PdqunxTAF04JiO2pQwv/vfte7wiax3zMWu9PryLbnCiE1N9/97fdQXxgBE4zzOuY
jMqpPlhZ4u2baZjJZt9DNBaxtvANOg0lcAN8Mo5T7JRsJRVDuyWzMbrlXeC8sH35emTqRU5nM6eq
CkZvxrGajNsDygahSERv/lKh0E5kJ+E49gAFmfDiBNjHp9BAFm00BNWfthSKSIWVQKS9t5LQ49RD
jKOYKRBuDYX65dZ9PSwca+ZJHuMPBy1OCoguZASfnY8o8tKALzev3QgEugWCvtS/B9YeY+1tZele
F3qagS5JwNM2Br7wtsqyCMaDAe9PlyTMU8OXbGYriIuvvVB3B1T+qfojF/XXHcgDcEK3hJKr0gXz
+bX2jc6BvgKRt6EOvw9o6EUGv4cVxiPCBtSF80WakBCvmJkqL8yf+M5f+sPLYH8nc4UghlPrrKFm
2EWanw0CDtABEBx8gs43KKhIOGpmh5CoA+wd/zykBpjUz/ivh2417bNxoWzBec6cSlanh4hThw1k
/5PPyLReagH65LN3MINCXeVj08s/cOuLg+SM972Ql5jliZLdsA+MuGaVYHjXbL7wcYo16YVGK1Dt
hOF6kTw/iMYzwg1oh4xs+22S+eJmLJ+5jdGKkgV4g5MAvRf1wyRwjbcX1vDTz/F99vG0r2eGU5JR
aMWaB2THoLOBw4w081lWNQwxp2Zyg6FTEAAO34XwQrwjzG/Git5ZRMJUBBGolfu/Ti2d2rvSY/s4
76B7cNP/Qptw88jkDVU77SoCcrbQkFVoJKeNrRGiiQGPHPX/70OzzgerKbRerSa1l2m9wz+sY5ol
2g6zasN8EJyB8XQ+EmNJukh5poo41Ytq2VTyVw5lFDlR7BvZ9xUHw1kR1Mm9g5fOsu0scc5iuG6r
f3XrETqG5s0ixPvLMgbRvnj4CHElxsia6YtPgDM7RmKwsZScXKYUnPKQ33b9SXodoUrsLat0846i
pvCO7dMqaeSJdWB3pPf4XCSDoPGdSlyLswHkPl7KmQlLJG46ONAHas5cbLhtIbQrzX9nu57n6r43
DfrXv/sgeWKVmhEI8jPX6GDQJVo+e1YCweqnl7FGtX7CVa2+mTXqLxSXXjGo/XWg9y0rw/XcHoE+
sJbU1AyuxUDzqSGDyil0kwGiqfAw0Ge83KQdc+ItOebvRvhw5ck6IN6bwjY/K5kUbTp1D0yeFyfZ
a3JzuefjCLWTHL66RMg9BlhoRwgdIRnTMwolgVgWCXK+VbjMFeeSg1eRT8c55lHKtrg+4rMDLNa0
uGz6jBBGLs51ulRDIpXiCbvv/XsGdAvD5zZVcG+HHZ/+R73m7/u8LI4HNhMnvcHy73VeqV39Df5y
bcGxyUKLuOs2jECqzztD4N7EdMRrsYDzakSCkeyWlucohYFSdrGEOi1G+ZSecVjtTBZxxXOVzc5Y
6X8lCxjZHn4VL549hXRSIeKCHIBOIiKmb+bPDe6mYvUoWHihY9QFL0G1MFIIQCAS9S1M2A66flax
pzqxH/eNZ6dX3wbH2vzF5fa/o5RnAXWxCuvXLW3qp0GnUbmZysm3WiwDikDoZ47EalPvn2irH63R
sar4KW6x+NJJt2XnctuejHfmxSs1yMAWwQoCLlsZLkbKQTFCX+HzngdfUapzPgC0BRgXy5Z08aV1
RSWjHySERY+OiGTnpre6dhORBXCVXEt+57ODeivvOt6uW5+O/adFzzC+raZK8+XIeNNztZuZLi1s
r9G9CvnMR2FZxrxI/KwRm7Ft3PmTZifAtJPsO4iYZmUek0ON/TGWrmaE91f4RF4hQ3EydFHSnoW3
VC+4ZgK9dfUaSMQXG0QFMU7y111h0cx2zFuNX5NycrcgpU0Dcfz4D2U3fG9RSjiM128cid/sg/YD
/uC1tunjASz7FmWGeLIUesHEQltfdQk92oUpcAq/KBdtHk3HeyauzEfwECOlRTTwstvLThuJS2n/
ksjcIr3UwzV7SgcEdbsFATMMGkhIAyd4CvXIqd3z65sYGqgxdVkubDb5D1zTq+t8Me2SjhXbZrNV
iRwE2WFO5zA+Hl6K1yH+xpz2xj3tn06oaMabzc3kGQnOWePsrHAHRrUIuBh3byOdM+eo63yVDbdO
QFjcMHWL8VM+XSUEULxVqRcwkS+lNiZdD1vFaFVx84O/c8/+TtwXqHL71R3qjrW4cMtIQ0NnJ2FT
lYeVUkUYMhbGBzGGNmx+kt1l/ADjzIt0RxTvK3/e+EWiGSPl36u2m9d5+nen7IIRHijzJc4Y+7YU
+gGnH4unSNiZJpAHfkFZ7FrJcMRIV+9VYvvNC769w7tKKWl0HVvvwEfAJFIuaq/fmqsBz4j8b9US
wlc+bZEjEvIXtcipo5UxqyUaV7NImZOr8BD6EfbGhxJK2GGtqK6q8/yVwZrBtAzcXUR5hGPA8Ibe
ZEeVQSX39g8bRufWoqRPfjIlvkRM+hudM+fHfbpZii4CNgHU19hjsYwNNY7tvHt18oODhHkMFEKs
MXaEwMT7QVroboUVii0+pKYZxRn3RcQ1iu3ueasHW5piaXT2q50Hi5s8mxjtVdhp3B8q3HbhIqEH
vjzv+NDHb0jI6CYhIhJ37lexysjkQSqrKY+rk42WXZ8CjpjPhzMikHzkCPVZKksBBqWqp83kKuWC
tfiixBBUiV/px7WqsfIhwT3t/7H3oc3WQ6CJYweW0ESq/DRxQyE/uWNrTmR92uqn3YUVzjR2vojP
qnQJUyMhXiZ9uMS1iCC81yr8hxIGZBWz0+/Bbpg3FkNx5Uu84rzxhGVGqlGYeTQa2hJCHfYK+T5M
7G/dCzoKO3t6bo7MQG834nhlyYBcDPsk2MlFGPWnLqfPY5Czj9eBru2CsYPtlj9ZCvuagqheV1Ex
C3Ufh+RjxJdWpHEl8Eb7KtoL/79cPuRdTNqTAQ03aoesKmzF5gOuZsP9OSOb5Kffm5hZRCqk8k7k
scOJeHGRiw4M1BG3AqJheICbeAoMzvQD+JgOZrHruGVxXtXrfasE1EhExYDbtUhSsNCMq9LmJZ/Z
dQmd6HPbjL2nuxNZC/7nxbJ5rjgdWA/X++vMFWC/QubNO7+zH0iB7/whk4+w49OAc0j9pvw0NhR8
lHgECZ0AfcqCxEe0xxqlYajb6pqnJ70Fn06I89obBPHrn8LYxQVzE1ihAZv1l9ErGi3yyS5Ubd9V
6VlGYR7OJ78mYx+qfLuWPg+YdDUT+FtKuVihJ6CjNv+hBnqR71nvsJwWn7lpyGEAQpC1b7gCWK+X
aWUgvETSHR+bwmJ97rVyOZUG3QXlckWskb2jQJ35sVQpJFTC0DSj36YdF35Xun0BDiYJ0MRtvve8
0U+SP6nCmUpytL7+yztjnJ05F9PWn7i3pCdPalK9xl7kA8rxXFyLw/TV3VeJW8rOAF0dg6od61aX
neXCZPxYD6GmBcuVSqinoWkVaTs2pMKu3mtbmqF4/ZklwGvxvJfRRxobbeTRE25P1k1e8Pqxa/1P
8UdJzhaaVUSQwzL784pUd3bqQ1PBWHWCda+IQBzsSv4piwxe8qDS8s6tNaSQRr7buZGeXPRplzyY
kUCzdIsQiLb/4oJhf6O5UbsOORA5/29gYXqZ7v3+OCphoBkBx8lOXPDvdk3zMvYaoAanIO1Jhlp6
TsQAN4xhhM1FeWmxXm8VLyX8+WOyZmsyKSBCnklhZRPp1beReEn+op/oKoGOz5sMARyShAEdAuun
lQFWpfhvH9JdWgZ89bJftG2Rocm6qF0VBZK2sYektEABMaUzIEp0tjmkbCfXm1ZuaydI1YVdaFdi
zCIxOCkF7hYa1FFZN9s/cWZiacmG+Zh3Kt0jhh2GjJ0jMbB/GskJQTzZEdtEiBYM6iLgCb2P8n+q
5VpeiAw89kSLNdVeuKyElTt1x454wJjZxczg8QHjvnDXJpzk2qn/O3ukvNg913riain1JxF0epTn
70mHaNdW82ix21sQb5WeeW5lroSOeH07WHEQPp4SDy7xeNQDMkNoGTEmiKXhsjyS7nO1+sz2i+8z
40QVqWlwxXD7c53X/Z7ZDlGo2WGUp2RRMRKTnt8y9jTeuBehIAsqn+fs0ya4L0Gjwdv1mft7JuVa
9LftL8K/Hhqpvy0IRyLTpfCIKh73I0DOT+2qOvJB+xGNZLvJ7mVYCzIWq0M6Nil0hl4ZYy3y1d3F
1eHiuHVSiJO964aBQQ1JYIBTgX0kY2ZSdBNDyJVn7QSx+r5jpNu8shwRtHaYM5ipFdUzCGf2pg9C
ddyXFwt2wbKff/nj3RWaSLU+X2aEsbBX4B6Er0ByuVoO+Nq2Melq9WnPK0PzT0YeNYqTvV4tp//C
I9ls0r+L/9saowEZBEDthr0gIYPKyvZBVfPfoGmAxfTAZ8WPUf5+1EGRHSX1vokGzLhvLuOMgaH2
YqF9FaDhHy99JqU3OgUolKxdTHN/swjZ4sPu/GUeHRnqHp/P2iPu5//TWGevIAO9SmJ8MWy5WoRU
5Gv/+UU6l60Pldw6LDns4FfPG2UtlkUwewDQkLsQJnGLfNsypSRXRupG+1FixMfkOV6RokVJZKUm
C2XpRy8T8RjdB7S+lzbhVH1147RKFnJ0VCvrCFj17BCwsZMjlQL15mn8b7AnSueE5TisUBGPT0Am
RobjQXwTRgD0cl3E786d7UcvKSrT263feD/VXo8oMjpd1lJq92iunl/2+yKd7+G52D5oYVEF1gXH
9Mdp3PW9sHZ/lBsVC3ZifTTW9fELNreDeVMintepagSeQNQfHB0Dt6W/7+W//xyyNh9GG6DEtuXc
12qA12TDDIZuoBKZnwjgszDsEjaXVGWuLuUagrDZrXozGIiDn2ZsdIB4IeueIPWO6cJhbiyUaVSP
KQzxK6AyjqLHls9QzqkUQQz4Va7h8JPADNXg8ZmxeR7Sqs0HpwNPEi1mJ4dDEb5fpfkd2YErAz1C
oRBZRcIbvsHLUeLvcz4m8ML3wAPWhKcEyx98Jn+DoGeIhFE/SPTvrzinxMAN/9c89O/EGSIipuss
Z3ofHGQXjAtmjuMuZ6/DFynoc1nZ8hPZjkhBQcxOkN8mMoZw4cVbrK1H5owpvnPFDvKhxCRytsai
tdjr4RmZQr1l8v7t9f4XDmOsTsm+AEdN3/cBJdMtJKTUvh+OroxcZcV8uikt9GoKkyjmxSVy8Y/Q
5L1xoux2W49ause+wawS4Z0r/RbqYxrPHJkM1lyOLvXwzxSUeAbQ6LR2gGGEH0CIaLL3bqOIvG6N
3/F2Q5rCdlxL49wwlFpb59zoQciXEFZN1e0RKqXg18VkaCu/tDXNyOrp46iYzOQLJxPmYiPYwRDL
9/oMiiqi/WF0TAmHBoK0g9McTcknmH0+GNBfyya3oPLV3VIJPkEfE+cdSxP866VhjRS8arSgybgg
auDeA/ueYGSbHq/oKU/Yh6ZyEGDgayYnc+23WT3e9RSE2vcV7U3Mqk4Eo9J7yxhDraB94JR+cKXc
gI/Ug19oQOWYfQpj5NDB5LsGWGWGLnj6WMGlp5oMVDSVXaig6LQ4/FK2MpjWPMKjDTAssSn0fvnw
f3pQZAXwJ6fBA9r0NGChMPW+NK5mI2kPn3JAZgNngzutwbwFHY1tb38mMludvGAxKTiOyTBhHOF5
mXktR+VuWHdJ55LM5MRKv5HgzNHWv1+OMvIB7ukxtV44PUsTyULZswQ6h9Tin4J7gIXGgdytrjO2
DuTGfXHTZv1nZK7j6c4nZBlyUiMc94CFy/xUJvw4cOw1+z+4IkrnEO/04zvw0bWvmqNcQjkbdNZA
R3tkJhnb5N7YJGMTRbwF/6iM3kHmjtgh5tL2ldkHKBoIgJDFVRwYlDM1507kbyL2NI0fKa2PtEqI
mVIh7zSIX2LaYHfH7Se4p4HlbwW8HWW7U8WLu3QkBh538UjN/cvd6Q1Yr+53tSiHS1huLd5umAj3
V6Hu7hqE2UnvL02dqytnkDgu7bUH9hBrpMa9iauF99qklBGPVqY/aKl99Rj1edWZGDQwBqUZmU8g
lYfJ1eJ7QJ7rKvhnJ4kC2YlUuadRIytYnLo54M4FgG4xHoIvMFIvABj2AZXY0hqkfLske5oI/A/D
z46W6LYNZ0foHp5ekO/60uil9d4GNfqeDzkY1A4PThN8e77CNzRE9+Txupe5I+1uAc5NOYiExDRv
WltXManIJJiQpsBJktO3fB+mgibDXYdptfXPuamUH/Ilxx6mowYRM/gMMhIQxRfxksITx4fhiZy9
O6CgitnBeLVLWbxl9QVreGuI0WKGSW5pUoLrVMVInEqCl95o+gIO7OK0G/sQeCudV4107Qxn9rrs
YnaEJ51JnsV+PAd9SfVFgc2EA9BaI11tCI2ylfllXFX39BvkR7yx5EeRCmWIo6+yaycf08V9YREk
Mw2cvMsw7YrkoD3GauR3IEwnt78+NvdpIM4pouByJh+Paoqt9xEBU5G3dRgW8vHkOcuSllWssIXJ
D7z/p+1djr3ul+OD1xSEhXd40FvuTnsKxZsOD1FmcMGKNDIxGohu5UvXk5V5Yg1ONI5LZbNp/mza
0NkQoxlqau3gNqLGDZnPDDQvuPR9ObMbVI8gLKg4ntHVZ4iVjAwwC6kkOeJVuR1JCrhGdHtDS8jS
uRMluRFdzpwuq/7tI+cLqy+vCShRSUw2cxAqqmE7ZYQA6CSfey0PBCMLjLck+mXxCDoZHhgIIjpg
ziN4I9S4KXKzE27b7FZ/tqPngO46H9t5Gbgg8eFsRqiDocONPX7xGP/p3AT5yyCNcTbOaqBttB6H
ofBWUHqwJi9hTbsVOUefqhQKPiBq4bSvascjyEFPknE7xpk9Z7qltnaBOjlGGj/Y87EeQCF+uY3I
3h7wZKjVVJ0kiGO+y5gYUB4cJprzTf/3nZbO+0ERE4PocVGXCJ/nM4uecER/m1aydOnLwRegzodz
6JhfXOZSvjTcpsIrYNiy+NPilRVm7jZkXd9+ZMNmbTu4y5T15oUxMwnnkwgTKvCT/HpBaaulgCdl
Fl2T0k22odBSqcjYGDhy43EiVBDgrlc+J6rU8nJxcXLxexObCHjmTQj2WK6yX2sQSbnxvChUMJ0o
t7IAX1A5OV+jRFJFyjiDhvZAvACCVk74WnltWL3ERGRYBBZxVeFpoXUbWVz7oJvi84XcGOR/OP5g
kfa0lEAZ2NHVq9Ul5ewARAOHDcHlGbfHWhKni6O0Q/Yl6qEy5ptrkEApkd5+VlziTlnTRFlTFYrT
hWyjwMP4Up3YYily7ykKpcCulODimT+rqDLR3sY9ARkGaqaP/fvw103pz9kdcT23fnpnTOMRxTHH
t/LSvFxDXHt680UbCz0xZbAbLn0J+O36hlpjEiLyNpdv8AdjpAOa8lDcw/hkMsi5gLnwiyHPtQnF
vQ/EiMDiouWKgLQe2NrkakbmDWmMCfdblMj13QrWn8PEiGnjufZa+in2bgAtP+C1IID0HCGKALVn
8tC+HDM5aow6ysm9CITvUBcDP4/zOMkdW5wD3ICB9KJai9Up0RDHf83oJq0390rxwUz5WECA64Tb
rzm0EIrChD3914kaBuzHX5fWHgd7lK5GiNJH47wE92B12Or7zsvD+U9sFB4oiMOSK2CXrKaM087i
KPVjB62nXQ7j8uRjf+wwsgs+7JQqcCfTMdA7QCwvWkl7Bs1j9fBpstDl8MW9ZdgyqRE8ofSYDywF
MVtiVp/LMpIJIXTuh/wOql3xQA3VAqABlS7baR/c5Vjpx1SUpNfFsWxfqIdCk11RxjbOfvuqgswE
MpauWiZGIdkZLgkuiM5CjAKI9zyJlm7t8/miLUxH3uUzb24aBowSYG68COTNsKXDhlnFcg7W42Yu
WFx/Phaw6RCJlUMCmto5I0zhk2YshFkCPa4rXf0L4KzhV+RqBFrl+udvemXyS0s2jJh3ODcPEbpF
71uqpu/CzQ9XgqCC+2y7bKKS4R2G2lUIjYxPTmbYiSp4poEsNjWWUzFq6y5r7tk36RjeZZEICmKT
n7VZADG8HCmnI3HowwC2XWNC1eTuWuc13tNZZO5IEViUSgkA9gUNPHKStMwXceNRK54CeIbKBqsU
or2/3RYFLIrMyIPnN+31YDH6Jd6CC3Ado3yOxSZc1Z+NNchkAJ8/ZN7RtJn53Ex4mVFjiNsYAGj6
mI6hO2+/JT29skAzJJ8az8VqcSYYRs7vC5yfqInp3Iu8ncxRG0/RJWPaIHry+ZX5Ynav4MXwl6En
fjbCFGzAh4uANKUlpcEt08fw96eGjtEmKzkGIHf3R1X/N/HWiTPHyhgnv/5sL3w10E9PSYccUNlz
CyM59af/GG+9r1dwpz02q2s/GnbSW7pRHpIELfNO0cFRA5Ejx4Jup448qtGwtLYoEGdg2k09HT0Y
AUJ5yAKxDZWFqYlgCpUk6iEXUEJMeagDRAHO7vtCYrZyewvkYWEIWG6H51CQHoH15IviV0SKR+Z5
y6SkvRXwxj9xQq7ylruWNRUUuaDlkaaAyuByAs7In2bmukayU7wopmn2dGG2u4w6me42vO1Rsy/2
MoqrumWRgIo5jx7LzxUr/DOXSci/07l6tNFSUH8L7Ym5XqHaKFV95Nb3Py1LancYZucI9jq3lKOz
U1pFMX8OsIXGjASYSKA2TCaFtrRd2e55Hz6Alu4qW0ZtT/lVe3L4apSpWs3kWfUL+geCpgWao96o
woSeEVne1w4ao3EYrYhcPRmVcvSJTDakW6XtstmvXdptcg/PhHI1b7zWQj1yKJAnWweqM0k99Uwh
kNUB/2xqbbyeCf8OcAgarmarVV96NZlXhxEBvyIJoaU10X09OMELd9IidKBAAjm0/F211wAZHGii
tCpSA9ivif/VwMfOEtMbt5hZwoqEc0oGZ/FtiQUjhDTZ4dMTyrm2awGIzDQd9MkQ7PMxVTc32TIr
RkQYtKSZOgIlWKeHiWHaT3PmGiWxPE1gXiVxlR70URfI0hLbaYFLjhzzACuC73E5yoxZu0BFiEpK
ecq41ZM8lYa0Kb0/iCtl1WgwKqrpgR5Vy7+gTat9pqDnkbzouXZut2dsxU4J+leB8yTFWu7eo95b
YnoJ9pKX162rPuc91veQkFCi2ihyGRUPgybnIXoOypK8b87mA6oM2RVd54ehjKtg7yJAf2KmAbFy
QeWiygNe6h6vEceoeMj2x9c1L+p+JrOMwHmtc3ZG0dhrmNBpd/CmVjOTytAhTqXd7JHqFNGaTV9E
Y03B0oW5PTslA0UpsnlJtl1sSBXH4Xz0U6SCE7f8hCc5RO/MgWNGPURuKtP9hAUlrTnuk8EAOfJ8
d1f+h7PVOYsJPIDHULpxU5Hyo7xVltRl1U8MfHP5+HAXCh92gAcB0Qv/bv9tIZePiRyZWermbyqo
RU8b48+C9auggDkGhGddDJDmez3kQatfJf4W4z+n1dHKdtIJw2hlMEAYHsBR1JK4X5U2ReHLNyT1
YiBsYEa5CZ0ehe2B5hN4KffzMf6OvfuJxe/0fEBcgxK5MWB1k5nd8Iy0lqOLhEoiFdEqbq09UYQa
RHizrgGtvWePRI7ib9EkDQ87Hz3H2ycz1NyhFn7EBAs+Xf6wWhSgsTb19C718eW7z1S1Cw7Yx2jp
AhLvW+1xE4BnWdGdT0fftElZSSLyqWtkufrQbCY/+eu7Hf/cVi2VL6Yp0HK9Hz+zHmj+LFkQlJf6
uOe6wF9IzGZC7sxX2IZ3H52gSrSm08+WZ5YWhh9vpe9i+/uryAykwSMMIykdffj/Yw0SqqpT/TkR
UQcWTbENWu1bZjzMPSZ+hfha7rtgI7LmEjhcOiEr/aGTpPQuVh499lajBFYR2XX5sbyi2xWzh/hx
bO4xWlKJVGD64oeip79AsoxNkHmka+1wjE7oUn77O3Qmrfhd9mylxrN+F3BR5XfLbeboOSW8COMA
ubfApjdqSD0uySJJTY+er+Ir9TNNhWijUMKGybs9hIZhEzH/53X/I3tc+1hBq58V07JWPZMTDdJB
gnQGlSGDlHfCjWNEQD+N+hTvlM1mLGT6Y75vW3wzY0AccKgRMmE02619nkT/mQw8amzUzBu6q5OK
raH4UVlFbjDAANkbKsWKBCokT0h7ooUVg9PCaRtzCjY2+/sN6oZvRdLjodHBYwqMaVpW1AC7n84H
HhFJ7WdkmE4og975zVS6HQ2myTjZvMB7MhHUnajvxgP4IQ3qJE885YEVUmF3C4aDvEytaPpFn5m7
+hDOBruM1OcUhAor1kjgqd4nyRLGSbU7oq5aNQEjgin1aO0P41G8NyZyTIR6UykYBt2KhnDZ8Bra
kg9pCW57mKz2iXyMDRti72LehGSt6T2MYmbi18WBFZHi9BJp/OvjW6OHJWR5BKALLndjrEINLdu/
O2aA+RDeLPB9rt/w1hhDi7yz7L65D5H4vAxsygdoXF+aTSB47NUzK0CZKdGO3/T/K+4TIsxCeKEr
9Aw7SnIYR+NMVsyMTE3MbF/IqGO5wZrf/LLcJkGGXs2lJwPXd8cseOy6BgPeHZH4ES16OxLsNBJI
TgsNXiDLJ4MSDKZtTbTLn2+R0bfjhZY/vyVc+YKVMv+R0ySoqjpyAXlL5gupQVIECJOgPUdJZttH
Clv/njsBR6RTliMQjPqRvnfAUqUSm88Q59Gfpr8AgkdHqwqhhlpQFdrzjt5odLQq9HRIs+1WrfLT
DyqBtpQLGdO5rhO0HLukZxyN8JKT+WvDhbKYC3OMF2WhKQe4nD4z+3Xdf2SKRmK5V+oxUdduWC0/
HFGCgzIu8XunpoPmkInRc9gQ1RBzkE8hQVfZe9Q+Ny7JwFxYFvCNJATvC3vI8uFDiANwWTaK2KDF
TJ+sPePOjqbbDsSndbnfuAqnuiRNEnBVH+rcWBSDDkdxDFh7OL8qWqJRAlhWVnCzU/ORWYMtDpDa
TXAQ4+aDslTUMjjOAev+F48RF0I0+XohObJpDrx2w5LCO9nFMDhu3FX8vjDoZoMg2nIpdYIOP0J6
5AmGWWAy4QDgdHePlEUTaL/7LoBiv+zdziVXzUV7TZaUG4MRWpHB0pl9MW5Q4QKLmzTteGcwMWlZ
oX7BjdLIG00LiuDb+strw/s7opk2Q2qcYH84UzSXfK1gb+kyS3qhmk8jGJTKiWP7AjgHbXTOYBH8
MRvuP1A53GnTdNM+q+awjw0hGfKJ96V3JnmqjeQn+S93LvrNTEpcUpaQ0HQ3CQESFuuQHJ3cvixk
nEYSC8/g1G2UI6c1isNe7YyodmrYWJ58OL8pnw7Q1ZlwOa5UUxOhQm3xVCyOzXnWZN9fGX2bOkob
r2KjuL8xgIYhtqOTEwwHys3yfDVHUuSaE0s//9noEiireHROUrTHufnzwnbQI5MnkoC5gVvnN8yx
lkLMsrIHzGFPhEMQaqxfSPxvl0yB/6WPwlvcHkmY4aH41ykfBItlEFfnWbugSupcdWUEcuezw04j
TazN9MdVzHtL1rjXdv9LSZyw1fVlssLgRgp6MTd+6tDaBxtKuVY7zNtmaTU7zD+Te9nFJ6r91vKA
xKH90QkQNVmc/RDewKcVlV1zd8CnT9e9rMOdTUnbm0Fg4JyE30TiRZ/NZ1WO2P4Nf4n4qOk0vUB+
BhSe7LiN0OS5k/5IPv3KOl16/WZ7S9cICcb2xh2iHC1opWLYSFp+rqbEsj7jdUNIkEZP0HuyP1Mw
DDdMqLJYakq3LHNX/Iw0vw2mux9rHL57UXNBLKH3i3/+MGRq8L4hnZGCyVLntXOYmrxYSdwdyf8w
K1pvYuzKLFtYOkp5t5COb8RDaBbevsXQPnDJ1CLZ6ixlWTg2wiRWRaCkJzRH7yeC8m3Lzp2dKAps
5s/pCAURpyJgl6MbvPWeQKoxI5B8DKuDvZ40khbkDSfOolzgKMsk2LozgE97xvpwT4YnzrBt+YpF
VCza8WUbhLFK1pVsh1xMze4oBIA6iTLHwwX0cBrQxo/vCli46kuyxVSNookkaUOACyft8eoOwB6E
n5MLm56P4ImVTSbQ0BnBxkWD6h9AB+IpUMcsgvAiR4ecPZZEGRayxfbaRPqkwXOFB90H4xs4bL2w
uOC/YGXyiCP9hEk4I0d9lU1ek/7xcTDJjnf6XWiTU9F1J6AHmlOTeyUFGOGwyZRbFL0Z2rN4vgvY
r2XPOd6vLhbju+xwsnOFVHphEy6Ov9kx5NQfehY1DLAEzEmfSZnndkD3VAOeI5pNL4hHLA+7Uepz
Sj9ck2YOzpthQ3Q24GzOxRT+V2yn5bkeYJOU6e8a8QBIR48JUCxejb0Rfg/mKW1/2umUkmFIG0f6
OXBPcX3kjc+fNp7tnxxCbsKMr50R5Fynz73ONriQVtrfqZf8cGISGdtculbCowyVZlY4f6Qzzncl
UhG+9KOlCzl7Zgap4UsCbUX6mCUK+U7gYldcN8KbrQWPgXDIfM+v5Dz+YODPxmYdgWHI5O28T5xF
703u0Xsdcw1F10iu4ljubef135W/VSUxx3AgMKExZpmUsnlNuD+50NBgwZTNd7Yz1/2G4XP3+jXt
dKSx3hLfXgV7yNx/1zQnBkOTsOuviY+QSluXLZad8FrcR899QTabGj63B+l4eWHE8wofMsCMBahj
6E2UV8Prn4+Fs/+KZxIqDb9DvCJJV8lh4XhIUvut6vkYDjqawm64LfirjLlo89fz2fwAxe7xWHrT
3gapBrJ1ZBAKCoNH73obW4zx1iDPDajj6/NowUbXEk+TXGYWMzedNMo0b0InxgNo4EV/IBCCX9qG
21XYRlr1wwp8kjQH+Hkp3ZxA8NNSlggB++gSL3E5WukGNIH/V5saUPSjxd75DEBUAPCQw0clq0nx
XCpdmYmDaKOpuDnbBAah1eHBnVoHW1Fd/GCYWJU6w+ItBdjx5R2iTUCFdLEVyDo0SeX2d8rFV+ck
78Z0an65S5eBSthMYT3tnPMbDcBf/h2Voa0WyDJYIK24hEk8xqwKrLyac8JlErQ/DryVrZCYuLum
XCPMXthxc9lNe9Z9WvGI2CMLqROEjexrTnYp+oZo8DY7XqFe+lELkmXkUxnDgfuvu7aJ/OGOR4pj
qkBsN6qqZSWtEAzhe9+EFe2YrWFacEm/ijC8PneMdiv3ZQhYSrFYVZzXIE8+j3rrTbe3iw2rErGF
paJQC2ke+3iHYFKMdk+Cveq64JzXHdmx+Lhf10dBGNv7WCexEW9YhHt72Buvj5wIRc6osCIeHIbF
AxnBI6NduojYV9eQhiWdHmzCYMAxYYkUvTcSY+c+Y2HSaBfRi0Oq0f4fa4nJcbTrhLv9kj7z4IWg
zEYxO/MK8shE5mQLM3rWAbbhWuokRAWDViwuUhB0tNQDdKSvZ3XEpwQslzVGW363pDcMVyeRKL+O
nA6NXN+5gPV+Gly3wQEKA5Q15Y5K0CpWMfuH4ibICXy+I9bIMdmSLQxM05BTqGseiDW44Cc5xyra
BjycK6gMS7zyU+so1nDI2IIiKR7JNQD2yWk15V5iivd2qEpRITMQMUiXwJnCL5dXy5GTjab7XVQT
qNjQF3IPteYImCRnD1M5o/cqhN7qxWpHXbj0s/H1GZGi1ILELvn3EDkKm5I3v6wFH0OIvidzbieT
rIu53MBI0SqsKsADD2Bj24hpJoI5hnJ1+PkuZ8Q3WzD4TUEirWD6q4sqcPBwteMZlw1zUqaq9Z+w
dIx9J1tRbF5N4jfkDuX5aN3daIFJqd6qPKse0AH6lsczHy+HXjLiEvmP4VdtV/WquIiA91zVJjZl
eu8O0lNTab80Wm02AzwEC7FgtObisc0lFTf8o5z1rdCmzurdtsi8khb4T8IBbmz7V6kIZe33IYwM
zXeFGQwdhsH+rBHt/TZYKzkGoGkaDsrJBAZfnaQnmpcC8A3awpUJv59DToz1ZWmXtfZITApOSOgP
vBiSW7OixymSkyGsw+Io17nzubmufxDjZLJP3Xv3gtGRJZA3w7ttLPCQjhmbCHq2SYUDUJF5PVMl
MjNrOZELMmefG7VEegsjxdrYTX7ajX3LZw4z4Pzm/yLQNLFf8IgbU1AakCKzZ0i4JiVUr9tM3jLv
sLVB7qPOlBTBdD6a2K9a3arU33zTWCaJcAd5v8W5reAEKfZ0M5LxXFlZ10Xm6uc23qFIJ3r1dTUP
Mn/UgHWlkOrg9uBLoHktX1vqSOEf1KNN3om8NCq5xf5ZuAYAK2bCH1n3iAmOMzTBl09wKYf30Mw0
4zoXZSY4Tg5bZlBXqYCDDlsmfSJpenoFG4EuG59fkHTAmsdOj8qe+f2aJzq/cp0k8LwWGQdb85St
r9ERY37hfcEcD77v6LIdOPjKBa4PHpRT2EI3MqcKaRVqlgsLn+oQZ3gBjPTzmGhB9XwzLpMU0BPX
6SHUwLdD5jhLB6KSp38WuGCPF7NQMaOUcyYR63x4GUAiM8oEgoV8CR0IG99/8q14MJR5paY7zKoP
mfmvisPUrLFzrOTA5SEONZ/q+iR1s18yeL0m/4tgFa7kytmcc3B7qjb+JR5PxEzwYnICRV5345ON
Y7S82gI0iQbECG4RHU14st3abWm1uaoF/kipdfopvLoO8BUn9yE7s6ThIxKEvVSSKEsbueO4uYv6
6LyE/8PTSmaUTMBIKoOVfdQ/h7nuhMHHZqK1zlkzdXprCOTzm6K79E7FDSUM4ZdLMQscZm/sasUW
PFlVZ5GfdIdECYvdAcNv6KsZnQ3K4kpLJFKq6fMFh5j4heiaOb2U3O3lfcqu34VkL7Fc3+uaw7zj
NucA6qUEQAz2FXuS9/EkY66eRgXoPn4r4DUDR9N28lR3KFdsrU/NXBT0sDYLn+gpDsPhaEoCCoyX
v7dnk9kRvBmg/Scnipm5uAn8MmOAYcB+gtDwXSfbFAV9P4RPy1bZAj8hbqqmwiB4VkOVLCoKTN20
F3BjqQWkspuebfYglskYU5uAuSnd4B/Z2OyNx4KtIY1oTJDjoHUAcTQZRRwk0uG1Whr8l4LCS+Og
1lUSI157JV4wpF581ZR0Cixis2S0pMpLfCUt1d7sAyvgrhOi/EMOH48WZxlXD7YtMl+JDnWY5kww
ImB4DWEj/CiYikEkQqtuTEsmFm2tawbg/V3etpD5k2p6DELtpAeYrGbmbkl8ObrjuwHPhmps3ONW
bDg1tKTUZGYmvH2nHHps+VnHa68vRd3bHTMo8VwjW3XVQCJiYisBGx2PiS1vDISOrJIkIzm7+dlr
UkZ6DyaRn+Oo2ytippDW4N6tOnS1vu4YlL6iB3YfC4o4C2fhzRD3WVzze5VDEM1tb5Op1MqAniFg
JOA2NjVrC5F5pdwscKRplEZbKAg+mSLgkG6Q6AJI59ZU+vIjGS4OwntFOquRrDu4zJrj4MSNmhSU
XvhrdryRZG2PuJymbAlKtvwLTWV4o9Mact28JlkoqLbHB3zHsPDpJ5e7ziYv4WHLHssOj6+QI5uB
WIla/pU+C7b9uW0g2nCasTIY6DzJxqip0OvIVxcm73sNvf5F5LAjE8u8WJPE9UuajwboCPCeD+S4
g1a9r8FaOSVJfIOa5LkAfY71hUe4TkRpWEQLEY8CxXn67UOgrCdh8lVqAxN1qFICCsprk/BP9xqa
F0O4V8foSjSYBM7M0PjnyE6CKdoYla/w69YUJ/KdABlD7OjfFWgWDXrDoW82uI39SubLZQoMvlQ2
fe2fKJmzbh7cnBwnOhSOnnp2n4QAdBHZdllq0TR4HIT9R5wQhEmjGjsDDyfAoDi3W9xfVplGr7qr
74Ixo0fB2NukfGY9XiQwwrP1cgzcwvXGiaxOXtyTleUxS5UltZoUS0mG3wBo7h56IJSAS+3TTddO
Lrly8WrFZEZkSZmX+f18g85FryqYfRddsvNyfgz/5FX0t2mchZXH1+hE/hakwvzWIgnClLboKkeP
YNBSC4QkziOOMwUBN50UjnoKSVGr24XFwIUhtrjnon4CUFUrF9/gn50N7HZ+oyUMS/X/d10oYTvz
uhj5diXqXDBYuQjJYAKevQuZ/e7/oAAN0hZY2vot2ubNMX9YFIKSuC7FpHFey4z1N/3FzsRszo95
QjxYa91DZLvK4oQtYOaJf01IJ1LQdhvBE2Pf4d7ZoNx0mtBcJMGzuufD1ShgxGoZ47LI60jJBejJ
7dv5BO3FAsgUUOD3pTuPuemsp/dFC3tCRNGiH5eGQ+rMZBCGYeYFtR9vnd8M0i5IYv+4fVyO7ufh
7VeNFWtBD6QzbZpjpqn7U7vnAvL6dR7prDA+T8DmzyS5cOPmpXJ6HJXK/8SxFaZz+yErb+9vmqsl
cNAK0y0KZ3YjxjqVUlGzj/0rYn7xBLLu+5MHr424dGf8VveJhwFs8zIRZClq6UVbP5dVygGjv3nb
jsDT357RPKOQh0pNiYRBs5P6CbXwS1FOQWOioOqHvPcbmeB3LZlW6QROrl12gnT5O4c8sUwRCBVv
imSeigwBeYZsH9/6ymN/Dws5TYoDr3YpXHDGAptTTrzGqkr8vDSXjnM8jvIbveVoxq22ssoiA+VI
1nEv5yNJSIdNkDaCsn+lGFsW1J1IyA9z8FuVCfC1j0ebwj4Dt5pOMhHJef630yBRhcNoKUhJCM5G
TXFHUdT0JSX4PY5xyEta6OpW2MqLabuVLHgiTnt2j2+CLqP94nDQjEku6CQ33jVlWluHKcVS+3vY
x/B0MbuAI/edab7rEyE5XBuds7AiER6RZDIW5rVI10ixiFwJunjdQXW7R+e6Uhr5xYPcvGvtAhmf
4WfV49OqAtYpvyuOw1c3EWxqMUiN08Kmm+0v5BhBwsc+03GMyczqC1DTgI6/uNDE3NNPjKjAEwBd
q+Zawrf+3cSkh5bktHnbloOx4XL2UN2HLjc8D8tBbvPijU2fTRglLngUi894Rl9VLKr4bz8MKKsz
rTmQF9Bxw7cogZhbXicpem9btCBxj7ZoM0sOKpLwBsleFFCRxwnf5EFpS0CvzpCudtfkzx/4e26Z
/hup5dthcX2anUoI8r06dFNDuy06dm7JUjjUpzr965GW9yiPdQj8ROfZLnNz+iLHyvTvPq9ghkyJ
S5qKcwzcqLyye+mHd+NQw9lU5hJn1PbAilDYo0cA5Sr7OuAFDSfbzERq+n6ugBbJ5pwiD3aT4rwB
jnWuzsQ0C8yiNwss1pECMjQ1j9flO5jsoPhZ9HrOikdUTBQZ7DB6U4lT/kSaiM37U3y1plHKX6QU
/dp5rTnAIFwbqdXei8Bv8vXnb3eU8WfMO6K2IAW//YXlYZr8ajfiP9nPeRFqMqlKbszaPZMyk85C
/WKJj4aq29FITRDN8J5AuhXvOg12euxhzIIbfn2ce/lyQvEsPhTbGlr462SMUSsJoOcpMr7i8DSP
4dLoLWMfTCjYYNrfBM6ca14awVfcxgYVr0kOGVJKk4DcitMLK4w+ujIZXtlJgMRDrmpGo+J1s0n7
gHTYRd1FY23pWRjZOvXOEg1xVo4wGVTV+MaxQ/MWqI7PTLhwRvh+lnS+1P/sVy7O+2qyNYly5F82
c4G3Xt9UZbVHT1lbkby0lfXiZsJec2pfku0atkCL7SGO3UCSRjXPYV7RFCRVFD5W/zTLwPw6Eck+
LThlsPbze9DlbvG3weK9U3LVN+vuKlkBsnDrhp5uDdu1xiI2w0ewHA2gh+d5HeOP0sGExihXwRVf
cHGGXx5eCwEOaJ9k0g/0SlsrKD/0Lxx4Hm5BHAMAs+BuMz3etA1ECXTEKQ830E9+GsD3rsCr69g5
gFpbXVWqjPz/U5V8j/rMT472ypbWDpFZ1mRWd/b8XF9KmUq4WLfrfSj0WIbdmZcyjnl/XKIFupU+
rRL4tzwlfqGyb5gDE4j43LQ9pkoRMfq5kww6GMowP/vKlf3tiDtIneKZVcZ7ae3HucQY4RoRaunY
QHkR3TiHgZ1xW/fw3TSN9libmYR3ougAtzji0zJ8YlWO+6yAOb87aPwzP/nqxQFR3sxXfuTxTmBC
mxtCZO2HhF3+3FprykDq29CkZkmD1hMy7gOeWC9wmTj2vHpbeS4jmURguyk79avMTTbEN8A6AmRp
5+SYMmqAwsquY3TykBKhXmcnPliXvwufHjlZaby1Xuw/xgVgL7ctEnoEFNXDL/+8rHyOJ0UBkjGU
jOpYySlbJBlnKx6L1rrCb1QNVhGNLZo9tAcizRhMPNt9lNRPPu5/YQMPiPtNnjvWu6o8OKLowFOy
Yd8V2GVkEPbauUxjYPd7W3E0+j9mXZWRVA1pRqCk9XNcTsUG4uEPV9T1cvC6EVhSaGi2ytz0ugI6
TXIBkbfqcqbrjS2442odWZVZpwUx2nFPu2sQBWosda9AK7HZnvaNb+5dd9GN7Qf9OPNll2NzLDAr
XCIwGRQyaic/IHs7dISf5Thk8JZjQVjwBnn4Ubf3ZaC8b2UQtbbU3K/Rk478GTgDk73nxGBA4PgG
Ck+3nTKyz0pJ9owZ0ioGin3Hy81Pq+Ef5I9C74MMsB3Ex2weiWpKlUVFOqLkFV0vrTjMf3JAPjWw
Qfl6PxFBaXhD2Iv7HL11F3+rFlbjQtmre/uCEdVpC8vsws/WxxjoanY9lEo76paQqHocaqaexmO0
7mjTfCbjlj2hOM++rdJoI/B6FMs5yz/+JAPuDhrwXQ3gA0egx674j7gdquvbrh5PBjIqWjemu2Rn
vq3dmOP3jaKUQGafchQwY4IPqUueV/90SnPvMjbs6GWpOiJUrmz+Mj8m3uYQ/IwSvhrB4LCRxpSV
1nhgTCJGQWEO995mg/LgFHXIYwtXM5IlajyETBuBEhecyyRP1+6LXlR+HVEFBSkqpDb0FxpmUxtG
zxIP1/Zr3oInyQeHz34ZiM/nttuMco8Etn7sl7a2IX5NlDgczJsAlCXOTGJbysV0AkjUP8/52oad
0m8m3sg6Q9s7uR0tO9cMO/O8EIrj18zGalOMw+HMpXn31dblYFcl0dr+3nVB6w7CbCOPMhYZ07OO
WQ1HiefL/oPHSxa77Hjo8ya+/LwAdLQJfzYgp4uCu7NMEYYKN2vVOdNggBrQyRZgnHcW8HZpjJQl
oSd93N/6jBMRIdBc4VOYlLpEv4qbv2nvW200+dT5W/aiITgb7QM84q6n2zCZLyyY7pMmSFQSmWmt
lOBYRuEuBFRYKKgjRKuGz0jn3jwhxvxXdd68J7UsLpJSgRIjg5MSn6tUg3JdcAE6R7dEN8A3xNB3
nERpkWRh8LDwaDlwv6oI/9RjdIJlDh+SYICRgU8I/ol0CRTwnHPtukfnC8wCeyAzcj3tRQReN4Qw
65mWDjB6MRG6b8qLm0Rv5OzpeCHSJeFDSdwshKigb/CAeFUpGgW8MSpKZscFrLb46kyNTeKT0Zs4
zk3KW/NMep60LS6cKe6r9EN/3g80uRHqzOQcoLAmWXOOtKKK3MsTyhMzt7QXwxAwniWSoWybLF/G
NaOko8epFPGf3lapQIOPiFZQYzBDUqcAfgG22GXKjyESKXkIrCidhlwzAVOEQzjlpHamPXBrrqaF
emmWiBOtE9RqkArcl7NQmZNN/rnDHjy2VOiw6s8DDWyvhNpbu3Lgjjo2HN7d+Hpwzzk+YK5D0r5j
zQsig53Ruq7FDMwU2ry+Xf8hUaBR5boZqoq4CdGPD8dqX56ZwjmatPN3fPlAVQPuY2alSfxWIpWL
/FNkm65vgQ5fbhzrhRhLw7nyiAJMr5K9u2kQN1TNzXcDJBiucwcrsvj+0bjkVueiEh+8ILcRXyiv
aQzZC/diFhRcRLenGTsRZn6h/TrhzgL1+2IBs1olEwsRZO/msg0YdlCExc4N81G6dIsiwNMlT50c
cOEcS4QTTkeoE6Fe/1NS2WuVGQ+DhUiRRO3NKHULnS6todeiwISN+CMMxQJVXu37hAvLhWDR+BD9
t3ubny07gvOhYfzV8fld//jRS8N+Scoi7VDoa5Yxk/YHW8de9N6s6I8hRyWckFS5Rbg7lt8jhZhn
OqTT6TTH7xlhf8iSU71IXuYrkJ72tJaNOrQyRh24kSFCrTAHeZCUAId3oaeC1cvaihroFOgkT9I3
XTeMTZw27i9Eh0bUZoqbB999UAhW/u2ip8Xk6lwvv3P+XUkspqcy4rGqe8XdZlxO4czJhyIopgZb
AfmawCDoPmNwQR+2dDAS0lhY7U+kNvQNpl+lrSUaFAdhWODyzpLQVaFLIhbO1xRxK4/iQOY4jvB+
kbdj613NcAwswUgkL1lSfPxiFsjtuvZN3G6+692kbrEv9VC8QlDdIEc3kiksJjgeGlO1bhmaLsFf
YcmJ6OXl7ZoYVdqgUzh7g6wjCutrCAR2AeTOMu2g4XnBwoT+zKrq3a9gQIkfmgnuc8/oDkjj5xuZ
LloR/r8diMP9ykpaA/bkRaBEGrzd7/bJWciwRaq++3M1d4ckqTbExBo6n8wlm3P7LXyVv45c3L8m
wZNbg4kSRijHewiFFqGJJ/ZqVjwfATk6w84ihbD+HiKE2s49+Tpsf4EheuaLOTg3Quq7/5aP58O6
qirmYYcYLpcFky3imnU4z/T207K3rl6r4cmuiNgESJ/DMV7l385H2dWE2Wqrdm7z+78sfTNGIjvr
ytqZrFNoemZDVnFTQGy/H9t2FXTpRBzHC38SYO+cTv8dHkPD4oQ4xW3T3UDV3aOE38cT7Z3Jg/IH
eR9Yi9qf+CD576wAb+oh3jLqurPIA/k1/0+6Xg/ohwPlg6Yq0Ss22POZoHMI0zCQx/3/GvnRDT1j
4WyvESTKVyJreF2/D1ljT2SJ9zTtf9QDN0ZicgDUak0Sgy0E5CnisFHFeCaAuR8HwRRpCqsnPuzI
yGW2NF+DHbvRLZjxs3wk92BgAq/ga8YGIBiWT5uumYMdtcEKL2X2+cSBr8haCQoBnHqMUlkKQLiL
Fdhws/2dnA2/IxeRrJoxr7HahyuK7xk6uTMLcdwAfTPT7xFT9hSKVsPDq7jntf2pQvHqKQoy2YNc
BFNDZDrFiGIdkuoWb1th4jR7+4hN6BIW6VtmF4wwlux2AzvAq7aC3BC/QLioow7klHyBeo7KiiRk
fAIzkRGx3muGwPlDPPSkIbmWgoHAJYjPHjRlcLa5dHFcrQ2IcR9X7DILo9Nedngp0WrZY8AYY65L
Zv6ov0C/M/PruUoftrd9XVDL7WKV6f0keiTWc+sCvCrtEldNDcLsUy+YLCxMomGLo9t6ORqfgS5w
z+Sk5TbFIIdm0vr9h61G+KG1xbgya+qNWU6c+0WuxRH49ior2amFpCHPBvMOjq+NSkOF3grNf9FU
ZsBNj9eDYcA3MErWTOjWis02oNHdVnMnIHwiEC9VEARYmEXDNsmxNtpb1ziJOC1tGpa4zE+IcQA6
mgsfPzyaObUqCsg8KgrtDdMwyeaW/V5EW+B+Gm6bPtRWIqkruKpKQRWx5tFjujVqF6FGCD3b7vXi
sE70IINUyUEiWV15yYFNr6fv4btk3T6RAa6ckM34s3K/MWORCanSOTF7JHChtUocfL+jBkRLoIlq
3VTlLqBbrhzDRVBj+ye66mGQFUHUIbnbHb9aNjpfjdAmiwGKffwt5HNagPOcACPbMga4YFqYfbtK
nbHhUOZWMVPGeTSDTwRA5jxjv47Hld+8gSt5kKnWQHxdSNdM6co6hW2UxK9T/BPGXxrU1lG0Fx1d
AOfz4CZUh/2TLWDh0RLMtjhEXwnQmr0nxYSOOGrrtRE/rOWcG+LAsh7XWtSEJfq9nSrTb0Zz7cIl
tELBomGnjpwCURyOOY1oMLEGknvCEd1u5tPY00moyjYAbHfblg9j7s/vfb09nyvZTAU52ZrcSUyK
atBR0Y2nFxPjKLn54gZcsYJuzyItLDHbqdCWC4rpi4hYDVvAdQTobSLPbc4Zs35o0osT5oGckAxI
iZCT7hCKTExGIudAjqMmEGTQH/CC+z28q8uGNmls2e8lh3QKTIlpScMR09oP55wFjaWLcmbQd/bf
PiqbqfqGIo70vmdSXZs4sYcqmm9e/7d5pg3br9VShrayv1lYJaweP0RdtVPrS+qDrZf/Q+v51wQj
+DebySAoH3phq2DTHPGJf7/Hr+Lx287MidOxjqhgzWZ+29Tyub4v68mvrTv3y7LAbdv0IeKbBLBz
1MiPhmVvOv1wqM2C4BHVtkMiEVVH7TKiY2NOtwkYsgdox8oswlUS5tzECEZ9kkIA9/yGhG1oo3e+
lvWX0+osv5fRC5wbEy8XTkiDq7cF/fG1D2jXxMcRd+pFC9Kx/uPEpiNuKHAdTHh3xhziGFqzSNVk
2K0wZeV89oPLKBCLJBibDEB/3AqoSM6vqkeXnX7U1ERn/Ba2QKGM0ea+48/bzb/Lt5vuzQqAeWb9
m8CsjQav1B6pzEzuBon9U3Q5mC8CMuMgH8Clbu2pSNtui5NVNiPEatBIzfMdY/GXCJg78wndyt74
yeTdrdLW2Nt6g0dFfvEl/LuafobvsxTzLxrNJJ0Q6c7NP/ZNGzSlmbWA1CeG6dHnN5Gh0wLGTKQk
aWHweXFxrftF5rcWRysutuWZ9HRLpTTC51life2Ns3pU8URl2ofIP/F2gRn408itlPRkrad378xL
SNboBooVooWqEuGfEOTuMOTRaOgtEmX6WcYsfUjs1z+NZ1s9DP21ATHOkxVI2SF6qhevxdk9yTAJ
XuTBnU9gjDEu5o9tZrM1QwwyESPXEa1iXW4IVt/Kmao/+Ntd9hg4JR2YEt/XP0eK4A+Vrp5FdvRj
+4WdIoQ6s5TyElBtW+qk4nYZEkKSVOzoZT53qGsvkC+nAR/1R/Zqwg9ZPcTpeBBDS71fmCroRfva
5MOLewWGSzaVD37UPxBtn8vOE0zhcPzpPyDLHk3lUY48CqLMCLkDrtdZC/1GYjOF69VD0vuPQ3LV
8kl0mALRfyqefuXHoGzrdD3EbWZafTC1SnUoIeeV0YWsMylTZ6XVbqPLRn/K2PYdi2UgKkAc+SC1
J+zLd0X5WzkC3X5L4HTMufZtuhGzb2uBovU22ucT1zDeNCHeyNSRWNQXZaTIam1YmnyatkcKn55c
bv7wil+dTUynluKX5Ey7t3XL9s0ahWjZehHrsAoK5GQnws4Y7qviwGMElGxYNIBQG7l7rMuEbtFi
6oVZAJ3vHxq4EVzWX3x2TH6bRa3j3XhRaPDZrnO4o1hbqShWoKFAiWymh8CSX0dWUQj5viXwqbi4
9m08/7eBfgpcYJpud/025X3ZDftqRC7BG5Q6Qn4D3r4fY3ETtHnUFImk0q+JG4xmJlE3UxzkNFNp
syo8mCNnXPBd92n+Oz1B7fxR+CbEIk7Pww9+ltyiVXx4tSsvU1cgfKVpyotAI46BsIbm4OMkJ3L7
sgGnvo2ae/Zsvc9YaRXZN5tQB5Vldc4CunlSx88499SXu8KLWOStnhx4D/RagmTGwkjKBXX7M65W
WWg9urbUy0vhBe6zRSrb2tTcI6kNAlJlMNzdiL9vtvkhzDrkcAfFC5QqwwFUR28q1ebOBt2pz1T2
z2qpMhLLl3DLQLCaEvkTm9xKL+FKJaCvMlvQKYXmrq5YKmxKcQdcGZWyyHjQoIarbQJnJ3nTbVW4
ZOdzsGG30wXbbQed2Br7nuaSiQRJSyrLDkJ0mlrMiruTZF1/fAfeGUbABXaLAQxe2EBsDb/KcOz4
BsEzpBfD5L/qNeosfL/1vcH6IvOhXeLvST25G2We0CHJhlrrBtvHQRNfsVsISo2Yp2sz6Puh9ONU
Im+jaz0CjsG8Tk80mZQAEQDOJuwVzXEgadP+GeEvQ7dtQHx15S1NZEKtI7COYMTb6WkCDg0rU1YR
EybVQQV9yT52bW2WkKGnJyfs2JIRE9TKASzc4ECc5WxnSHjTugwGOwnYQkJHmwRm9tZp5zm35eQW
o3fz1PO6xKH79jX3Wl9dPtcKDpbAArgdiTALLqgPa5GGTNBnttamUFU0iU1w1Q8DGif8KsA6oQwY
MkKMtw87YUDzHNbR5iVi7YosuobKTWzWB2uM0YwZ4ansDvat6ONeUqoe9i+V9MNM0plzoEl0jE4M
wDmqLCfrbWYxMUwSQM42ekaakWd57BFZcCbGIPnusaPdITCzBMyJ+l7M/hBGQ4mLctRf7+2+4WCx
8z91PyX7xYOlkZXN4eNjAOMWjZuzzRN25tz2x7piIN72n/FX4f74ivzKknZCCsE2exsJAOy6Gc6Q
c5OHfqvjGpLx168+ecuPrDQGTofyWKlSH+MMQLK/tCXjscFnFVhwn4BMWHwRh1B0atjKHtXjOrv6
w5bQvqay6Q0OE75m/O47oZwyQ8Np1I5KJtjCnnhEolnELMR9eAFe2MDzTMz7cklv/OUIEn4Knm1S
bXJj9bisSTtfNVSBOoCgTVEl9z9fHdytpkgFTBG8uOz248UWaB1tTc6tHGmFn8J8S5gY8jaEINjM
woO3RJwt4/Vz41sMFtO8gZhJ2Z4L/zGx5yG3oq8qjNNuCuNb6OOjAAHD+IajJ9FE7qEB5v+BqA1P
2ZBXZDok1UsDXx6sAbkB9b0/4oAba6D0KrN4fCLV2kM3BIOLGdHVeC2Px/Xw2ZCfwBy+41xBX1ga
rE6k9PLV2nt+88j8jJh1bvs/aQIh/1y4ZvhGRP8EoeDSdlBb9NUCnkr3IuMiIHJEL9m2JpYQH3p4
UExDM4AFeMZefxvhVdu8obQ+fa8jdFm84h/Dd92YwWUZN7D5n5/LrG30eZ3T4kIzfw/8XqIT5Op3
GBsNqiSEF5eYa970TcmFHacRshJNIWguAIw666wZkSH7IX0uljrDTA92CRfy0zCmBmqapqUleUCr
jDIlMefGq1Cef372wltK3XvS7sZDvRnG7oc6q9YNRetHCzPl1u8i/vkhtXQgvo9g21CSukUzE3PU
xOwvdOPER7l0EWB9YFbXWeRaAaMmo1qL97wIh0Ipf4dP5CxKFVtclMfCy+TUoSk8BT3UD/HMRCG8
jl1Zk2deIQ6WfQX7TgxTa9+uhje6qbEAI2fWp//cxomkUcOqJF0tgiPKujThi6VOce2oR/MgfMBt
EPGStiAIe6KCYMfyLm2QjckW/nTjgCdLi8jATEfrMEtxL8ysxfVUVm9W/FIc+cGSegMSXU0MJ0dw
AxdvNBE14urf5ZZPoLkwvmU2AlaN5MUHuquMUn5viw2Yxr4Kpa2D7oWV4lhoGs69G1JntWnYJiJW
9mOk56oMyg8IJLyCyGxAwJvVac3LjFLJemGPYB5s40WnpHVDYenR0cX3JOrxwSc47bEqnSaRaqP+
87fhZg0yrHTcWkEUU6UmT3dPosiDZG8m3FlMsAyoBrYz+e8QhrbQnfd+O748PR+72YShH34nL2aA
SuVm7orL1TCV7sD1sBaB3w2yHhjL3X7lTeoaraW2hh9+m4BpP15WBQ6Q6jWG080LbvBzUHQ8ND7s
qQSzLwXQqbOdtQ3yOyYfMoQOJfkhAZLA/DtKHjhFE7gg9Ju6FH8/MMSxt16qXrXKywIt4FqKFzNi
jtgMk2W8MFG9Z2w/cjnZ25iik2stIQLa2KsUe43nbOr9pL3fmt8cdu67+evDVrntP9JPfScot7/L
8oMs0A3nrAb/N01dDgjGoJ3c6lWfJ4lM82D7UcmNNmiYBmiuROxS9lvKLoQJ0OXAeIu2SnHCCELE
k3d0q4WqbOBrz9lL5QCLewmgAt7fuVhFMDFu0+bqoulT0xkqwKefU3dBp/AD5aFSt/1fMP645YnS
XQyRbQZImKcJmbpM5okXNv4bpM6xGu1RYW3IZ+Nf20EbHRVZcPuviLh/xRzDWbzjnpSKh63R5VMG
Nx8eJL+Uk9IRukTTqVop7AoDdnMR4t6cpaDXNYZH9ec+10FJzTuupCF9kbUrDGHgZQ8Bu0zYgr6c
B4pRvn4F/PMzb/A+S6TriLSzTR95SzuOSc4Is6qnLygBrlsoBiKfwEdf83muY96AYoZo0jIfckJp
luL8zv3KksuEWySC/vMsTcI2chYi+Z1eypqJWV/6k58JlEEKEuJTCbqBgS3Ykd3Diw/iBTEdfAHE
WvZ2gS61rBzNfoCiBebihxLeObJG6vcUI4UsXFhFqDAF6vW7Zg2M7HMvJvQEc5Pm+xsXaZEULsed
Wfj9q0sOB837rK6Do9V/Pyy039eQLot31yE+nCTDyU+AeUPOpsk7LSvW3gbDqwkLBd5eJhDlvGhc
h8VqrBBeaq5q0CvFQenYMhE5WQpuC7kZxnDBsRMDionW5hV9ltQ1LhyqzGnSR31hhwFYsAFG7d3D
H3aGy1uTTfe6871wF4bbViycKYS6XgTqgk+2pwXHmNQqZiL5zEvdbnurIsOZlVW+GnVEZz8T4kUG
3T/lMuj9yU8mo/WM4oh8O96qv+5GsZrSnwYos8fOoiTQtOdnIv/5MD2Ar4x0xMQgT/H7wE9DUJMu
qoUs4Ucnen+WWpllNGujHNqKQuxcTG7QLK6rCq0TkX4ibM8hjlIAMWPBBVW8/iiAGJ8L3A9uW2HB
yO21b+ZluvboMdW4fCQA0Xf4T6SSc7VGL7+OuDgfTWL8/xj/bxMv9Fs9peuBygK7FUlWPgEwO0Ks
m0j+xfeLkv6GH3M9BeXtJvraX68GwX7tKlymckj1x8e96GwOE/T7Poqs3Yy9Ypvax6TeUmRPWNTy
NSlIgyZiw/cfPwSlLzINyyB2wHs55dQcHA1lu4WjPdnMtCdCq9uHz56xCXzr7Ct15LulKVcj41CQ
M6HKCX8iCiadHBvShLe1Yu6gC9ExMqAI4DuoG8qAHIVJ7C5zRuTJWcnvdN/9RyJ8ClFNmTzoXgrY
16BKcrIwPIyaKBgWb9SZXy2Wa0yeE9XeX9ESiXxDvqOpToL0C6KGBG8zhhPqar85cdc4kdIIHWWS
ZDvi7C0EEs3+6WUv4j9bE+/Ad5m8M/Eas1ztEzqnxdirbj8CcgwvYvJlpGrNR05/licCapsRpWKr
vWxXJwg99RXh/bsaA1tTX03o3gfm4wmjjJE0b5+dwnAAy4+ysvi07uIow5EG/Gws/F8fJ5vCZGfV
AmlK2fBnq6tUl2/XVnjqswl/L6xsARFfLhK59zLLeE+5Ick6X0X4mMefKrnQvYqIANYnC6iaKwDe
C022jePsMynATgsVuHQtYL3GG3A/+sndnDNvdSRH520t0gSrx6KRGa4SbvH5OvjwMND72x3dM9uL
CtM8xiKQD4bC0Pdf7qIuvre0843vT0ZL7J2jl1Hh+xMxaQfYgF9U2P3f7jVOgzetRoRvSmdPRglk
lsF11/tRRTHKKI36YoDhWc8HS6j7rsRDUpp2GLwx3w0U0v8azkyb4jWtgTM7jfmdGTCMluuOenUH
Jc1GVYLiPi3rnZBmZ1AcX6tC2h8Mo+UvuEK3gV3Puh6JwSXYLm28gjx0lNmaYMeUGLXDRVLcTnpc
rO+N3P3eisxWz8WHldWPxpJZiSkbTyX3mHsR5jl4m3QTqrqhuXFSY+PkQI600Nv2KAG9N/+NHEvY
HxqQxKoX7iesOUeVXhqVD+gYB3o3UImk8UcxVx/jRoIYMNMIlHOu5C19pPxzA5TnQlw1wbALuQlV
8eHk9XEsIp/1aIwlnQ6K3CfUXDrZen/Rb10JwE0hCinKdztg2BPKrwDIwO+PPdbStQ3yMW3vdtIO
EUUgpFfEJ9xjo+j0DimBunmY9XHngQkgWa35l9Bmjwsks5ZORWj/QbQCt0y1hYEXYAFY7gfKpg+3
JlqR75bHE5V9iU1V08W0bvlpOgXz4iG7DLBFLVfS3cTQIUV7uVtMxQ96Apd8eNNoBnzARoBPgvpT
MLdeqZY5Ib9My9TqIfe8pyqgK7eja47xicZC+1AFbabBVpq9YgIUluKQzr5ZH5Wll2z9PZp2vntl
PCzYmy0tle99CSGtCN5GQMYNtfR/QD62XvrOFzyMghpwxm2jqfLrgQ2ACsUaEvJjyrHqIGxAxXx6
gJz5boPBqVSSnRZ0lYYgu+g4pL88ToFMOyxCDy60EEvcRU0KHzbX7IsxdTvvAYGWd0ahsyY9LWQF
LGCazjJfjnILPd4eVR1psr3ZUdJBld0PlUmOfgfgpM3E7sF0h6EovoFWZ+QbS9MQyHRBwTuvu3f0
zxnCTs8ff9rU1z4ZmeMTQ0OkltLYa6y3v0LNIGlVwFg1BV7fteJDZy5vok54kN6Z//xQf2OtjmTc
p2WBr9c9Zo7g7RkKuKrKG0Ualihn+WaB/lFelCByk+2J1sM6fLrPsUaJPRfalRknrtv9lsBih/FS
pjC8yGCdLFyObbvP+uOJ2724csGGgFS9iLlsV9A9iBNoUD0Vtg3GvFxjeIWMbs7cWUUby/mH1iS6
jGQfxCpUQLTAYfIkUOBGPzUVBmeiMvoKC5u0RA6/Ki7yVnMZ/ZbcE++e5FKS/bbi9VJCYeWFbW8B
Gu9JjVsjbuQ2neqaf+bOlKVS30uClvlEUbncQMvANPaRP+6bixPRQV54WAUW0hGBsPzGmAt8ZLGP
df4U/a7qvWhFfPOUxUdovjDhhoV2Ev1rlQC74xrJpoQtUGn8p0qJWAaY6vCZ7rg/1T5JvQwWsJpV
xaUlsKEIUGAsjGkWsNoOxBkecYuP++s7t3cjsmu5plDwa36I6RX9RSVDlfYe43sXW2b+LODCq50I
D86YJ8oz1+yX1XYL5ZvCWjV5ObFv7Riwv8xi9sv1G6lIHUXVOQ1Q9w9UlIO8DAKBRbQCkfLRHaXj
yYJqzu3iHdk3R/zX2+9x75izTLurdHf8YMAVR/nDG/xd7yrDenLkmyIutX5UiXr9wYzbzkQGZWtC
Lkb/Nm71DrkqBDtVzCza876PmKfqUILIJ716+T6ZJkMutcP0kMT+eN7kKN9f/B0v+nBjduhEmV3M
AHuaXhZsupsAc8JG1chCJcRkAwSU/IcaATWtO546uwTIG/1lHDrwXxLJFN/rMTWpnTgjTfTJEemI
64clXK2pPZO4Cz4IoYaNYGyf6ijghNNDOxz5r1beXEokGL4D5hHjQ+a1ioEYC9KaZIAT85XmubyW
wXM2v4CZMen6gjXxZcGWfmCoxIUsKPCFEM5qCwkOYCEMxayHV5yCy/RUl6CB3YQQOsGRL3gK66mv
MkrwNPEersF9iugI0Sb/UzzxJ9LWOnIqF9EEvSlvMwh8oblysYot7RVGyLO2GjLVcg/eQh1+id3X
Y12/c/iKoHavT22ZZi8EXzHUJz0p8ex8XwwldTZ/o9bdcW5lyr+t1RBy06iH1r8dY/CLHFBXKDja
OrbQvma3303Z+EPt4X/I1nJ9JpYr/bSHl+UFouFpqOiw6cntqi7+Lct8sbE8ElfMxpG0oD2NWyu9
UtnAt1Ogm0jra3qq1cPzYWmkHfEwcSTn1g7ZzgoUD1fywQ9TgKIDjGHwwYBqwT5DlNRSxRjic8Rx
E7a8k51IpsXInkUOPmtubMAJFYugoRP28LrbSEuZau+zdFraK1xwYeeU6bsv6MBmgCAEMCHhqOeT
cz/zyfx2bwWBQHUMq78gHq5fkVGKXU3f8JRwi4bli2xUGyk84jns3scR1nNCUTbqbedOv4lFd+Q7
8lNsSibr9yZnP4zD+jvacjobaryYzDgahNS6r2vLpRYvJY0G8VfbIHX8C8cF5b4Q7wb0dZvCSB1d
rPVfFiQznJB2eL+UX1plB5YALYPyLIhy4rf2Uyx3AicY1OAh8iquoYh3B2b/kMhIRzTFIlmYYaAL
zI39gHISi2AIGTEmMePqp8LoRfANoMp6de+LSDI//SEhDJaPy1GtGZmycBZbDmYJojTxZZwrvcQu
/N+y8AmlKmrJ8VXoZi97fDd/iQcsjtdeLvFfOIVi/S5b5JxyX3A9D2Kmbci5i+F3jkJxE64YX+Jr
e6aUFA9N/xAj+AbszMYdjrIlYdk9AA4XD7mrMSQHHh4BkY08B8PvbFUDkaO67clBX5wGbelDE3tz
Ok52rbdH5U8ulvwj8HYEqBpMwT0GFGfcS1hT23j654Xj4LN/KLbmvdKwc8T7xiPjU2SoJ3ifZiRP
CK4x3g/OpgSBL16ltZJWaDJRD3XLeq69Hf61X59qPn8ESf/14rIBtJjjp3aokRfilgEGYU06W1Dk
pIAvTnVAHDPgb7gn3Q1HUL+7ZiWOZgKnt9bHlrAmCxs93Bqnhusnus0Ci04kpWABOJYu31F5KdCz
i7leAqe1ZdAa0vgvTk97zy+S2fbqF/oF1Ouf+J9iE3VIbe5AO2fTam7GUDGB7nICX2KRvjpLgzQS
qyxbOIVXdaVRRoFsGLfnwWnqpGsHYbqumigFb4ViMMt9sLDEOy1zyqiDp0MpzvS/KnGpJ2kvW2RL
O0B3G1GizIFs7T6lArOwIHSmIJthudSyC+juLgrl1FbyY3JChf2d143O9uHara+rML50+IdFjtwG
WU3EO1LYYkMzET2l6bBBo0SkNs3gl+3MeBZfI47k1JLu+s7FgGLb3HnY6FrHIXuSxs0YHZtNBM12
0IdyplOJZH41ieranKrSClqlyQ7oB+wUTWjuEeUOFfU8jxt19x0TNwRdHluJCgVHIME9R53SSaOp
tcWsZobB7U7fe8K5J8YJCENKTUf+vOcHWFDCWIe9h8XJEkYx0stuaj5fW1KNxFjfAieG9SKxk/wb
ymGCUe0SHoXLaXruayfIAVPy+PNRSPinaF4/hIl340SX8UIt6Fq4aWZSxBZBEEZmMpWlteNuSMU6
0CHnUwBGaDO+/6KQQQCP2VQPuEVmfCxGhbd12LIpzFmuOXubi5i+DQveLlVrL8raBf9G3O0b0SgM
MV87bSE3nZLh8b8d4BG4/zQEDgZkStq8sctNYmtVi7ZmMuVV37I2gBW0ASd3DYedNewun9gvpOt8
k9HAatUOqlBAhZRC7djhDTvq8lz14tvOXKb86GqbFGXYDFQWuqnYIHW3gy23P7kH9Rdcvoa+UacW
2djJyoIRr2LHTg7Jeo+AF1/5fFcbATQ/dsAnXX913xiH/vgG9k3GFMzcLzWNZu5xfMxL/E2ajgoM
gqcOgamJT3PLGyS8mxwBBl+zgghFoQaizIfcyYz5mZ0bhlxC8bi6cHFTr/MJ3zFN+p6UqLTE+BgT
AKTu/q9cIIP0SExgc8w9qcGBRnljIBsL4lV/eLJy1KeeDlEXRjRgxJDmcwnAG5PA3lxGkfiwFU5W
7tBQLOe71Te1hVUMffFFnlkiODY0JRJadj2NkDbPFDi1DBu2mtLCsxclpf0K0noh1YzR4gttr7kU
2Or0XmmJyDdpw7lwoy1c7sWfU6wr1gA+3SiqZg9SKaw6txRvj8nfFqFvAaEl/KcjQVtAbP6DcSt5
XBO8Fgp1Q9xrkSf03K2KYxKCo4KuNc0uh0grQ9Kfhh1tyYH8/WWM0wxm+r+4odOzH5c+EXbGbtjM
mfE16i/Dil137bJZuws+U96YLJyqQ2g24JHIDkwoUTcLr+dp/vEQ1uilctXKeYQ+MXaUC0JphdhA
MzE8tnXOcjmvEB3+14/aXPeIDYbXPNTd2Mq0RQVEF639RWb2UZi0nDCqJHD2pE25NgoZswMxeicT
LJ29DWozMeVoVBGHhQuPUsfLWItO4hg1cV5ZEjtfgIPjgxTyQQuB95H5nhiy3mRjcK+F5YK7Yr7y
jNBxK1EqHYQIwV8otDxlS+mEeiY33FX3ge4GEVUrhppLP7hnjE+t7E4KiZyoNkJMwvjpdzqe3sPU
OLznimH709/E4jMvjJtZ33LJz/dux73DLAJmlv3GERc3Ldm44XQc2xTJGE/8i92A0u0f1DL+bIHB
iRs0CWNkAVUw0lheVzk9SDujGGcf4H67EYMHxKy3/1iAoZ0G1CYYIE4h/rDOXooD8lD62nd3H8Fl
3NXbcSM/1Fjwl14p+XVSvPIBHwyOjtb6f2bpg0Voonwr9V7nz7cQGQjgcPRgXmBHsqHigBb+a4jG
tfHUuyOjZMlUIxAno6gsP7dAUfvJYusLWEAs+GL5hPsDYW2bKQ3Js4rYu6AehNIkZs0oZ0rP1Bxi
W0bxaKe3lDpIEicvwXtAoIVBnFPZA5ctju0kC0oODEbW09Nhv2E6GDMkHdMHgnFvSsd9+v/rtXDL
XGiC+hvgGbNGx0hvEdM93234O77Vvie60tQxkfcX0KOGqjE+1DbaQadN4a/vZvtS8hicRjQErLLo
BQymdnNLCnUiKutkI2Z7/sJzCnlgsIAiCQMuZ0uwH8hs2PFPgkCnFWxW0fQv0K4Dym1RJXfCtVPx
0PPZMYr6lyp/S+yThka7ifmAe25rAZdAE7d34jMB5C7YuDtM0P9NH9NhWByyCRFT8vPHHmt8Qp8S
U4f/X7w2cgkOs+k45yb1TLlFKYhNm653UcYs44sX6EbUiMCCVtE5HaH2n5nyF1dMa2nLHfDpoA6n
/a+ey+Ght+AunfyBfGmMyDSPEk9Vc2LxJMGoz7uEK1MeLuAPOY8VqsK1k+0iyvDeRl/vfCBJDpwv
eO+J8Q+YKaJCBiJWszmbjrhkX4sU5hUNojVbvw2P2UrItaGi06Le/AGHxoi8L6gvk/7ob2vuw0W+
g8rsbVRO+En4+ab84q23etiO3XLNZO1istrAcTfIqd+Tuos5mVwuWh7/DWWaL0obBBBQ7G4wLT44
9ZT8S9rkbjUa92tovY4aKOGg+ffhOoZ4YSP6y3yFn+AK6+8hNrIGmtu1RUckThEJZqgIh8WZxlB4
6nxOq7n8dHdDSTXg4U4oCFZsxS2u6Z5h16oxtpUNImP57K7m38ejrWDt4ESONb+XbG9T/FfCJ9VD
A9m2tBc41mV81CFRdLS3c0WKzlT37MBkDvTYUlpLTfVK/kfJdNXP8PmvhRERvd4Y9HCyUnKpzdEw
ra/oj2NrmEnB4ZKuwAz2n0ARh4QHnUS9IwfT6E+7yesppqZgy/PBjlAwFLEbE+z3vVGgGOGrppLA
Eu5CYtftEizNKYgSysUAXjwrA2JkfJ0fbco/sK7lZeiPID7KelgDhTXbiwgCLzUYDp/IkOcodc2L
v5684KGXpAqg8nCO5pkE6H/uddEA5N610leAkaCEb5k5NDWCWFQijNiW8DqT2AoZ/PYmYSr8eeZQ
3wBRpKAhTna87HfHDIAg2Pk972+/K569sy+9TeZJI0vr/tAxYgP/TH3K1g2Zcl62pjcZfMioOrTR
xJdaDhvtYuDfov73f4oj41MzGEp5G+I9bUE8phubR8ycxx0drEeCMkUkFMwBvoJs9WO0nbwnWGir
bt4z3CP/8i27wHxMSuRCCPGuFsW7MLhtq6eGfwBG5yuK2eNLIauU89z/6xRo1ADW9DFUiMSgMw0J
Rffv1x+KziAAu2hchhuebOaoMCR+U6JEP7xx8uT9GyYaSC2dLToegrJZjEYzO2rPT4xOsAsRaO7j
DlTwsYy/P0mH5AoRW95H9IGvbVq6cE29YIy5ax5GC9xLLAnrXx8SIpdOZVvj9E808DawXpuYI+Q6
5uXXn0Bnpe8QeyzJu0MwTM35D3pW0LpSA6bjRHwoPo7qgsJ1NF5LWtCyu+ynfSmau7wwhMFijeJI
1P9cygfqBjCOS38Bwm1cHBIz6DUXSjU03VihIekExpbqb0J7PD+00CkJU1s9vYJNcbPzl8DArz4p
BsUs/NfZBn/3ovcYElsmVB9TqSGg+hw6fsAFHanfAEVb2PU0RxUaESS0M5HUp9MUQ/ifE9mPsLqz
Kp5atXu+/wddt751KwoddBLzZaHI+WvvjDZCzr390tCezGZoGlTCk/QdfRy7K+gG3c6NyjHbMpzH
wG5aCiQcL3b7D+QO8zGnjgP5j+8gz7GSKZd+VzNXoWBOuHcvDCvf9YdanNRQCVuoA5PzQv+eZDVL
ptycPMsn6bSnaIErlYvRwYuAWLUiAlT8lKJUIBST/QKRBirP/tH0KfBzUP/9qUvgQM4IEd3f4G5C
GpSL076VQLhGgPqATpHs9HTlZ8UBWjyQSoVJJmDpu9dcxVfKhMQjhr10gCOdtr8u5qJgB2Akz002
qw31KypBGw66kCu4EJBhqlHd6NjMD2fB60tbXck6W24CDRFMgyi9zegR7zZwhKI9556yUUW/RXcy
OymGF5Uava2uZCA+ZBCt3Akp74/0qRlTDx9oD/i6Q7//IX9fXBsRec2dWmXJWDLEEpIWtV4MA6hm
8hDCg0s+7AoUAb19Cr4BCdPJHvYEODXFvN53TWzrP0a05kkpwPjnPugvVPcjD93aau3+I2Ofkz0F
GeLYadsQzQncBiVt5MG4gf8hctDYI7sefEzM8GOwxs/v71s5Ra+PI4rbnVvQmhCDpbwSEmV1ffHi
e/L8hCUuSvVz13Ije1OPujPCiQhVFQplLUx1zoH1/7em2gk5soiAuN1XIQ30VhBLaQZffoBzR9dE
waBiFSc7IitRKGbEAJy12p0Z1zaIjxW0toJc0cC5/ueeJKfZvs68GDybg4Sd5i6US1+CrRj/YHGC
ty6cXPpdF6fxzbT/0H8VH8iAhM/ZLUJRc20Kz+0Y/RborqqKL8x/9j0caJLuUUms6qlwlO1tlsRd
43Fqzcoo1dOiWygVUz4StBb0ndjtywHfDqs+gn1bJSk3iy5VwY7oVhkeRKKx9o95NsCfJyOH2R1h
Rr0hu/a9THwbOwa9biQrMFe4kwNdXXqtE+ul8qa2W8RIHmiyscBPgasBmdzzINs9fn8Ab+ghSY+b
hit19ThFapHz/EmsxNLjljal3oXsEv/IIXd5QvRDdwPB7MF+kgs7U/qcVvKboiM+N0qNy6ihwQDK
wh0iPxUTyw4WQYqe/BYCw4z/eJMkYtjxseec8JkqvM2YfSlG4RH05qOvgDCxJppMRAWxilCwyEea
xbMhXB8R6jXt2EW8bUp+MmGMWdV1yVdDdwEf3rTRzcsYMP+ZnESqC11j0G/DIIP8cDA5qoOvARiV
jNgHCm4EbIAHCJB6q2wZoS8/UXxgWXYVPmRR6fR28P8uicTCJMtgL+B1cMSNKwCHzgIakpL978HP
5cdeE3NeS8gpvHjWA29urUbBr1pfcqsglYcSgDhSWjghyywC4AfY0tUGHt3M+onX2lm78SWWsJ+m
uR4puk2+cU3x+iuhivKPP+xvtAPFOGKpuITI+hulEbLXexTlS4ovLhe0BQFtnYW+o/RMmKF7ThQW
CUSy78xm/sDO+JsqkJn5dHy0tJb5HFBTBrL63FMwh+wub6NfZzB3fbNY+byUIqLU96728d+7bXg7
G84kIqS0yuZczOrUYAyBFxOuJUwKf/55SBMWmhA+5ee/l78Fkl+F2xLZhw2xZ9yd5zeSTsQwqsNi
eKq7SMV5w/2t1Mq1zWNIE/nK8hQXsEUCl1E501/vsThecuX/40XOM94oDTcYBkp1kfkF2TLyKQRk
iDZZa+Pw3rrsNCufKj/RQhSxcndpnqBVmL6hSh7P+Q+nEHTEaYJtmnjAL1Vv6ZzPWIWXkikguP6t
GdfDg41FSPImdg+zzyGI6Y2vnfx/7n3kfQtWFbCRgY7D8h4ttn9josPvjsdijtNaRsZtcoA0XIzo
DbEoISVYnFcj32BK/62sS+O2Rw3svFa6j5XvaR0z022zD0Ia45ZeMnjL6fOcZDAnvSEsoiavxCO6
Wy14FkTepz0Y7w8aWt4qVoDvxG4qsNhm01l78yKpsM8+nI+Q2qekAdaHtsNvk4pX8PRK5Dk+FwAe
ElCsHkkJiZfS15W8IXKJt6Y3FlqAttJ89G+drZeunYvzRncvRCQdNX8Hh3mVVVcEyULr5ocuv1sv
aeI+HEnayUfgKTpQUVS4xDr6j2QeGXaFT79apwomWuRxZAzBJNsDB8VC5p6ighSrjPbTvOMmK68r
fwkQppygamXqNpm6tOIzOOOsoVXmqWgI4mJNmXjlhQKbIiT+HDXPrkpOFKa/Sl6unaSLEUph081Z
c9qVVxOAl1ogONC6+k2G6PdIz3GwhbvSkUzDOl4NpYARvW6/rtaj5CYOniujRLH+e9H3Jd7KX/dX
Q1dyMh00aUj4/deFvTuys7oS48vmFxu4l61CTTfo98ZiK1JIsHj4bxMDLvrEgUR4K5/TQWb3VmpH
Y809Jbj1cmhdooyUFnydrDEZmwVzyg7Me3+wlEZ+Y/9YjXwXeFL2wa7EORT5a8bKNU4NBQFWd8jR
bW/+033pUpLtSl/kq6DjqSw/fFSM0bhNx4p9KfOjAEYWuLDHh5G38dwwEe1eo3JuLXwRwGX4oty7
daYpklWmZpAaGrupQ+vA3ZrdhQvHQxBuN+aLw4HfTNY+cEILlAL3ElYyOe5LQbptWVNjFt+gL6lX
y8lzGG/KWJtWYfP/lZoCvjgTudLal9MVS/WiaI6wk1WGDLRItdeKaj5MQUuCpFv/kvHOjY7u+0X1
MRSwomxUWHh9ACI6nVD/aaG5rkIpyA5mAGDgWiHC8//RlK7h5yQMswuKFu6BkCq7JYHN9qBq3NCp
pacmu4o2TxU8daFGLW2tywgHWK6KWQiOSX116mEa5OCQ5eglpYk92lYZwjBvJ30J7P6aMSWF5aoO
XB2jXVZoyslqbHhKXxBhBrO/ER8gIa2nVPN/t0iEFF/IRSEVtBmiLPm0qj5c2QG59BQ6gt9Hywwm
X3XgtjKUImbwRHcgsjnFGTN2h06YmjVF1stUXZuboWKbZylRMpyEwxiyywBKSWU4LCmmIawcjB8T
uQ32whRXVsUGvstlJAREiwBKLlY3dScxzC0mj3OCneRmrj4LpXJvezGbNOLXudZa1ARQ87vCqKv5
l0t7QhawrMXLPejl3KBrdnFgbuFtFLuLJsqs0szvze9e5DS1znamizx/TfdiCdiw9GPisG2/lKta
t7fvuMe0TJEbD3ZDZx8Ry5w8tZhgBjou1oByh3DuQxhzO/oiaWONr1Kp1ebzWQFPtK2h5Vd1GJ2A
m3YCKjEsoNlefUPoC07mj0C4giQcRKv2DTXD887iP1TvR2bSQP5VNKe96KxKXlDpHJ2QElkwMebb
7esh2JijA5hGtWC/PI5szezAOKTJuQBBg2pVx7v1qSgN+RGkl//Odw59zdKy6LyAwRp2jeq6y/UZ
C0aVWjm/uGldCZG0oHK594Qn1GM6Y6loSclZmQTaVk4WVmCr3CrwDMELnEYfbs5jstJ6EbcxcePo
cQ0DqM1vJOdJQd4pSXwD/xq8vnohFY0nXwg/Nzb68++2d7HQdNgyntYxkEwNm4jtLv6NBQQsnX9W
mB1TJHZHESRq+ufTnKrH3YG2ZIb+GfnPBhPVAtfwRJTy2zeLlfZ4wUzB4k7/ir9Rk2h8m/kw5HAn
PEe95PhWJOU6kKOSfh8dznPQLqEKwyrLFqtZacPA5+HSmsHQoNBd/dJJ2W6m+zySwqo36xesNX5a
TDcggHZcCZ+5Q2PmMIaxjkleCIGT5HUOSPkV7U5hLfQ6W+VY6BvVizzcUZiW2jxUbvGyWydqJ+Yc
v1jHj2HDXsUD/PnuIiRtjXoN8hbQ6b6VgGa06U86lxRFS0xLaTZ+YlwRXwNwKk92ry70yBfR7f5k
yCRXqM5NA3f0R6NXEO917GNKYH8GZV8ZEvWAt5rKLcOAgBSl2MGwnpRORMWAlHRUzzJxsGnAmA+e
PVlpY+CfZorez5PAq8NmfUuJGUo0z9Rejz2MsO0++Ct8UAM4O0HJ4t//iHB/D9b8Tp3Bg5FkTPId
lSRRY/Iev8wl6BrxBJ/K5UzbmnpHfU9l2z5gHLIYP8AH1htqZTPUgWcc/kMemIC0lvz5JMNVzrXL
x/YBm/xLL3LvsaowvMlIRip7araP/IWIt5DPrYpHJf9gAz3A6iB0e3FDF/qOlXXi/UNz3VniaFdJ
lvYEn+CkORaMMOilNuD/OXb+3UxrgccyToxmadJIP99x7LTL+7AiLPt3LOPzMeLNJNN0EYsLMBdy
Ul6bqL4yxAHxCXyHgu4dZJRHY12TspteIF10jF/kx2Ydn1QctUl3d5rN8ctHWTvRl20AmIAvvsHl
uK+vzqa1AyvMJTJQumrbeh0LoS9bVik7b6IhVRrTAyiXZ3i6OivR+7TlUps7IPJUDQ/qG5Y8IJfP
5lOtWpINfglhz7QFz+LW4WuRh0fZrQtfzntCqeDyVjJFLspn3yZWQVjWGVZi5UK1egpAAi9r37ER
2Pu0bZTswHLW/Vq6aMb08BjV103fjATv/foOeLk8JdvLFkg0W9ib0hbXNE26P/y+uZ5Q0GVu61qO
K2GG+yTjMRtHjm1YAVj49gU3qM8rSwmST3j2z9ry3xI9gad548BeSXXV5kqfzunjbXkcX7sWPG0J
DCTYoSNk80IK3KfUgTAUhgP9FwgwzP2oH1hZPMEyYWeRDRDxoaApTxM3mNydJBuNY22dGrCX6Tp8
gkK4NCI3K8csU21e3FAJ5J+WjKMthTzRgcjxL1/q62VodkHM/IV6mzXXmoMA5K+B+Z6z5RY0Ojq9
xH3cRvRf4nemPFjiaHD5kB46oLBs516D0Fc9RFx5xtkSfe6ULZpI7Srg5RfmmkPz0wfXgOB+plES
7wLkQ4yoJQIrCdGp/SOgZDqItvieI8ExXECrV/xa6fxydFQTunvKzOiZ64KFnJMzNLzDSEH1+LRO
ETedBwDA/+FLUKFfEBWBJJ54x6GfIE1KXgdiYI5/cDdGXHhRpU5Tl35k+a4iRlx0ZXFbkTa5D1KK
5PoZMWdtt/KuxJ0vNJbE5WFatsQrQH//brnRZus3qOAAqb0uiK8JL2c1nd19TTpLmlZlVxI+jg6t
RJxO8u0u7Fcw5/NIjxznfQNEc23On9ZjDNPjytwZXUoigQ+guWlEkKa7TvrIQAWGSl5dRmM7jBjc
akPraY2K1AhE6Xm4rxKMJYFk2UJ8qU9jvBIwPAMAXQY5dGHPs6ZhMIYOANb38ofH+6Gig6jriiWP
Oeel2HdbGCQpRfFjONEF7DKz+B0+ld/SELe7nodHT9IOfcA/rOXjKSvPHTPLpwMSNnblDa3faoHS
7Ldj5sqHLD6ZqprkQSxfwZD9LpsGIUrGx+npyXMwnxr3ixqIQ0P+xTKpBTdSIIPayQXFAa+8fEtQ
nqZtkEbjbNCK6tMVGX6n9hElvAbxcL+xSh4upCzfz8LsF5uidIH1/YXa9+B6eDW4Q0YzRS/rmbxU
iVD56ZJIu+nS66vP5bWfSCFgvQSvFPYgX3ESn/prVeCRsTnAi110kw3EC6hoSjmt9FtwXkFxYOeu
UY4XIt3Domg3b6WGv7j+OvEBzhAXf7mj80/YG/tkeG/dnw94Z9nnsyDJL+1XRk/nYFdBP7EHdB0O
/ZxoCWn88ZMFvwtMnoOZYJqxje94v5fpKAGA9jkf8Kv9HvGuiZPTqE2L35o0STVivUPGRdjaZ6+p
bVBg5zB1cQhrS56Glu56ktfw+iXj97LfTWcdSHLI8depvGSfme96OMmhTauuEx5iOkvmt3UWWzV+
E9xINbG3dVsmDNupdaRelfzrwmThWNTnVAooB47tpd/Bx0MsCyrUf/RBs75sc3M9VsrXRk24qo+Y
UA+2N43jE/XRkr8sHyQKXgyI5RAXgdNT3ycND3XFzSzvs9bJpA5jLy7ZgdDxGtLluJseDlwoTzSF
Jgt97p91a4t7CMl7rs1Jtpx+Y6GZ2RFDNfodq8XBNgWyBRJFygEFs3HDP1Y33FUkZMkLX5gP66WC
2FLRTKCoHc6gb6FPenVzHOtfw+dUqXBFMcvHS0hEvg2HFj3iyIO5vlCxWmcvDl6H+jMeNnGA6ccY
5wtPcyenvrokvYXyIe1hJ2hbze7srLikobL+U+hKFhRZY1u4p2cphcsQaY76DNs1qvIwWo2ueHc8
B+dIYvQ+UyA9slpZE2RP2uLUdmC+WO28gRy8WD2Q7BaQ4A8rEmKTBfgqtbbv7JlZbhgPPsZ+gTsP
1I4S5TYcEGCVWTDp/h9ecPt5ETvxIye6i4THpn/bivDE05V9ALjz2ZQKAMn/hdekOffKAWLYWd9M
ZRfUdRXDLrWrRoB8KJm7LAV3j7t+1/xpNIIiZtG533n+qTWHVCTuLlfatvj1PQu8ic+c9LqTgcta
6uW3zy2NcQVXnIom2phw4wcP9JSb8e1jE1ePiNNsQmKviSARst8yAvKNNKik3E2/adl0d6ELo25i
eId9viJlg159XNdkxaQjD+8AcCSbeUJ8sOZ274B5oCjbEu9dUpVUiODbcX3jBW08QtNEFUjg9Ns2
JuUEKB2KlcZxWnF4EkrEeaz8QlQ3r3s0DyUhJ1KUmqIWBNkemJmll3o82R4185nfk5PfB/eUwUuX
T9hkdNqiESsGK9bB87xkAHbiiHU1/GDn2VpAN02tFI8M7LgCowfXpu3qnc1spGFwWewHpoC3HmuM
LSw8RH0uy5+88PU20OsH+0PeJ/PyDnZ3HMnZXpyeemol+Er2ftbKMQ5sLK+FKxZ4iDMdidZLI385
bmaQ9PFqNM7WM4YrVzgEf/KWH/hRzkUNKyMOjbBPXKljIVgAS0T7hi6BeP3ze6ISoM3nY/mc1cpS
U0wv1vrZoeVDyTzaCpwtWBFC8tix5DpJJ6UwryA1ZMVnv/MXfd/4gqp16kM6ua1bvYEImcwM81Td
zVcR+7n4Bb1twtaSBH0ff36c9slU2i/zn41DIh3C8/3CDwM1fsPuaHSOQu96qB1c1IBGbRh8Gchq
2k7BsaDydEl6QyPnazk4mpIv5f+sHpbt5R6x3Gis2JzscFLSinSqat4oi0GOKOSopt8NQ7T+sIxJ
67SoDdQcNuNAA93LyFsRR8LJL3OeXtTAL8RUfrgp2v/pUl3AS4JzyU/wy7ZSSY7drSeSSSPQkJUl
SA14is9IDZ1FAfZKHPeVajxTl2DMoG1S9j+nF8eIGApq2a9qca7sKP5tcYZ9eqdon7jNjQjhz1PY
RXURwuykuwc9qFXpsrQ3y0h6Gmc+Q5ngzEp1IzoxTgf+FQXBNxRHWY/tpS6a/0AAwO0UEGZGr/8T
OiWTQF6R8kiVk7dvtX4rduksQTMYlO95mpyR9g+8qIiJUMEPHABHSV1jDcFDIXo8FGwixf1+yXE0
QJu6ev/EHgiA6g+sKliZA0UxigdgSSRnx0xztscyWs+xMT5J4FMm67Q+OuEEUhozr/7/JipFMYUs
uoQg4oX809M6bF6uM/4AuGRRxCTdfOc0fkXYW3qLqZ24duUbyODSlogwyH1ml4IAZ9SJVzs42R9j
UEiflAxdyTAkXDMTLb7RxV8H6dcTzeaRXOhUpnZpeZkfmm8kQY4QoefjLhvwXS0k10FMelkYxiIY
VkZCf6K3u1MOlJq2c2WKMd1ogaqKKgTFRxklHFmiBclOvMse2XCpt6RQ1xMUdCpsjomLn0L0Y7Ta
83aR1L5X8Y/e6WPVSbUp1VhIFYIis0BwZmotbKpIwRybMwMEekjbv+QqxJFfzd5Bczmac9MfpgsQ
9omePawxZSpcBFwMF1J5NmLXV88560oFjD9KkJQdKNmAzfNM30QfGNCARH/Q2p+kVxArqdjtIfu8
tOHoRYatNHxSotKMtMEwIu9491bUtcparPbiGIcHS+eU1JBLNEt70pfMI+2w48uZwLi8QSsLhTZd
ziNfjnNKqHUqV+RDx/3SBte8iTa2Js+AkIF43O/Ra6OaEtqlre0mUfCIoBuMS4TmL9XQ3NQg/d9b
b7gjEV0khpxISbyxdh8e4CHrT2ViHpUG9DafnQhZvvaffstCIOqPxe/XBJFDpPBUJ+p7Jbj/MaGS
h3/zn+ia6f8ougnnzmmZ+gh2yNNNfJqzb9YXgFRuK0ekYwej/fAs7B8uU4gpscP/vNxixp9WXUeA
eeHDeMwr8wmZDeQJMO+PxJa08eIkStRCAUyRUntVmKvgqWZ4m/isnCfzhVvaJw2eqb4ASkA6iR3L
dbFbKEwn0kJ+8C/6zT7CrNuR4VUnDHqQVO1kDg2Z9iL/LD2kGYK0wg/iUmvqLlS0AAIAo406x0tl
bYRftU4q9n74Ln54RCwpHeUz9xzRT5KHO8c8p4apS6FknniNQeqig2sBDuZ+HuWcxlXqFzgV2nQi
gGb9nA9O1CdAogn4/mdSY1/MFVAjYbeFUXwhxJbH9ocmpQl+cuHs09hTN+TQJQynQAivVw0pzlfG
tT8Uj0K+f6D88BjI3P4Zh6MXob7OxmDiRHutB7+S04LfwWKjx4A5USNDac6mIdjO5NfmoxBsAU8E
2LuB1TC8g8bGaG6iJYQ6YyI9ho2xL+zmncIsrUQqrDZGRzByt4gFhMgeBoAuAuGM/6K3qyS3QUGI
nCA51JFFN71PI0urYmAwbQPH0ZO5PX2McxWIDP5SdWid32HR1tcPN7T4wqM2zb9n57sqnfbAaxMl
c76pVtNgzRytRPAM5/ueGU32mIuZOlqMQskDobhpJxoMOD430zwLpnOpRC7CtZWerPNmYd128/F1
RKe7NjyrSEMTM6VnDgi7ioSwPOkU3pBS8eFims9AzCV2xZbMjgSRzj1HAhC3lsxmjzLgmJJQq7Co
D4knj08vJjbDmyxbggqjdfB5isiNcb4TryjL57BP5MFiW+fL3yvbgcCiE0WTno+cE4TQPD5R+H14
a9t+zMvj0PtbQknDoxr0MeFWRLO50PvRiPiaDLm7AV+PmyvjLaGPuh9Me5BzBVTPIiJzmm1ocHCW
tVp9tu+DqEFx90j6AR5lMCc2oQNhOr17wAO1Pldbctk5vgimPvD7Z2Pjf+HA+DYXSUUnKns+K7UU
Uv4Kmy2XyVX6YPZl9BuMpgwWR00SGvpTSefzKgVnBN7J4JeVjomtfhmPL9a0LstNuZK+zpEdvEu1
Q+LKkIpg542JZ2eO8ZvSdPVSL4XCLapxIYjsH4xOl5PNEBXms1eNedcQKoDuJy4J5IZMHf+s23OP
mG1d83w0q0sJBMU3ue75upcdB5Yrcb3uU/fTcjCXjc3KqloMBUbtyAUgIKNvHhHhm8awUUFRiU/g
GiTPqa/8Sow5pvaTrq8xen+SVwO3Nusjz5Z+1QJTWO4I+HZGI8fcz1Kno523K7AJfvy+VelIHS7C
By5qHTs4GIX5SBV+Rpy9V2r0PgcJeHu0I131jFiAMcTo+N1MB86R/9xHpY+SQAwUazuwYoyz8l2D
G4KhuC8bev1cEiC2Pxcxqf2yGnmZPrkRrl5xb5qGdlV61fv/Ove0WJydbRT50sYpqPvio1z36zuq
/YBDPTW+gpxlPS7huODyEoF5SJ4lXYVrR3iCHyi6bUiLoxboZ0RanOINFGozFNk3ObmcvZeBcazk
7Sc4jJ+yaXhlwcnk/m0ttgWFqinmBt23g/d4zY+oyqCJPakuz5yvo/Y3NQbCKzXncWgmSVGBax7d
zyvJbLZZ+2ruyLjuwrEb+iCiHV18DwQFx3b+hzbZ5jJYoBhBmD5nctXKyWZmrBXLMvtfigcp33qI
rpR20rYK8hTQuiBO6FD0u3IslFkd1FHSEyFLiKiMJ2Uaa9xBMEXwa2Tbdx+cldBYWqqDE6lz9ro/
BcdRUE6d8P2dqon6d2In6JWzLM7xRYLzAnUoFo1/nj7S92qaAks1sz+0p0pRv3tTk0Ay/fvlxmKF
l3Zauc92bPUEvSSp3+INPG95Fr+XILXsYTUbpn7MNI91ceE+5ozaUuwgsvLrdxjCppULyuu3RUNl
b8aXtjGQSb9fSpN6wb+AuCaZ04Wwc+cWQjCNpKWpSazSZRKiZ7Ji4V9Tr8SswhE5I3hRmP5psi22
GO+bzATAbZ9CqMRTxHEWhzpCGYtF9OnFjPXPoQF/cbdaT8eVSkZAiT6dtfOXsJvPZ3RQuttZ8Tml
d/P0h8HzLcHaJbro34xLZx2NYpsqmd1Y6VfUrm0t028LTA93ZVIGqjETF4/tWS9PXrWaHjLL1Qkj
Hs5ONVVev5ByWJioeMwEp22J4PpvEK/vrfE0yv1pZ/rrTI5kWKH+l4VCP2f4e75Vg11LpZxWmnOq
3JzvhLyNvyo7n/d7KhPN0S4PdsBtzEhV40roeBd96D2xe9Nx5qfGzQVoOC97FPkSv6yYIFJPn+Os
IwY58CaZAsiuN1lT+kUbhgSY022LkUs37HxMRX8a1lRwFiF2+h9nHIj3ooyv1uLbdKwddLcDFZus
+nZHS7zL1YygxpVZMaDsf8Vk48kdeWw6dIXHrrJKCpX2f/WdOEqJUlJN7RcyqEd8e4jL+9gINyvR
ULr4JR05u2LLpJ4cAc4mikgYySBrsnnqHpwfXm+AejZMGuFzw782bb+qMCWbct6OtUA3YewU8Ius
JfDEXpznxaatiQZF6Q7CTveBhDFNqKfGVr2wzvb4B17yNpJI6G7mAjrD96BRcrwii+X2ZXOhqXqx
toe74Lgj8JPOCdMimsAahgGuwvrmED3lmsHBYebmOP+ZJ01DVhuKMpzruiQccPW2C3EzDoVAzBkX
j02JxjwKHmu3xKx31AJRGSFte/mXg0mPMRui7xLuiX+XvQmJaVImMOfh1w935LxXZICL3CG+rWe2
yGBydcEwpWM9UTb2P6DSFKKYo9cAyEACKRhZtQ86RNf9l+vBroST0SGfjWHaVwR/53Ie0lzz3s/j
c8r1NLL7oCRVW0MDdwHyNhmVz+3STH5zxMhnD1D2cNs/kgdfYgGy2haxj7qP1ohWr7vf++sMhTWT
hMUoH3UEOqOsj2PuhUTERhcyRJ3YwO+hQjIO81JZS2dx0ktaECsidPbzJIrAb9Ck4nRNnV53p9V7
w0SI4zucdB7i90jSVZoLwZ2wcVFRIxP1MBUcmcJmwee0cN9mGSpyGlfQdAWIdGzcYtvDNLMI/BQ7
LngTHyn/OFayawPuRaC79vSqhvDsXD5hyH3NRPTU5fIFivpPhFh26GpUCRKkhMnBujCv1l26gVD5
wHkg3wxCTmn+r9xMulgAKXY6tpNrvY+xhWcY6NxI6NpvjVeAX2vCrgXFiJzQueCsckyDZ66Fyx6B
t5yTVJ1CjJCNMTq+lbcA+KhQP2OFI+kUn8kEWQK4T6rXSbpuKUI10r88emSxzpT3ybh8qb0EW+jI
Ubuu/kyx47KufdSk8Iyr28Z7xClV/ecmZb4PLk2IjwnrAEyMuGeU+D6oHDLq6AKqaAqxRGiAJRm/
KucylbKBHAfRhmNFyzNSQ8IcMlmnqtOjNU3EfkVP9t9K92W+61SCQqS57PibQIbVrGVN+pV6r/4J
HO/vT8PXcsx3MmF4ppXNcnKK+uu1/Y96ERyBuTrTmDye8x2R27Il8ddE+cYnsE5dzmhJCzgQziLw
aXFTCmO4zt8NoNjSzWrjTD0eFHkaPKe8LwGC+t52J3BX7Tep6wOhx8XQgBQDsP0GCYy0i1oOlE9v
0tvBWuB/UeAtGEerPfTtymEG/TngLr3AxhyoLA7TwgVsLnOZfbxp3JH28IreFgzODcGWteNDKT2N
F7AGuFr8VmC5NbrviPbP1RS42lYzCahTI5K1Z2/qawO40p7SDeOzxbT0GJRdWD5RAYvcxhL2mRjg
oJW2flz/4b9KH80fK0EJ+UYZrAFiCjtlOfYtG5+0JO0pqMRCGtJ8RL3yaxJ48HonFqnKYoSige36
quJRo2LGT04HH7BhzJPU6pLeP0v8QC6vDuLH5gHVCx07paCA+LeXbV8tcxYyJGItP43t8uvU9JTT
XXn9WMGs++5nmJee6ouBE1cFxZlIMrWZf1G3cE9T2Be7/ZFwp1vdQqMLXAk9tYPw4hQTMqUTgAKy
mAxscjt5oodKhwjcvIt2qrM9oNdcUr6fUHWj3i7oN3DAB5toissQEvI9inPPsSwjuBiT9N+gSH6m
5K1qbka5ivwfUSTO05d+fXMY42SXJGFHUhEh2IhePfx8sQ/0GN5tgFxbcxzkCt9TycrbSk4bPEyv
4p0hM3ZfTUjB2wdtxi+WbJSF4szPLKBfw1hcJLuFdzO12SwEX0+m+szbC5HxUuYTRfEUMrRiUTMC
EYZrz+FrABl9rXZs+aZdnqIUkIBKodbr3s2+oBojqAHUAjS/tvAStR5jV2J+YlDt7lZAMsE+cReV
EnrXK2S77AWvpv/iapDcLoj6c0XKxBM3dwtrhCo3yBZ0+DLJPrIChGGdB096IQ3UziDpmEZgVib+
5/jhpybZi3hww1fgwyR1n1vxn01WdgdK7kNueD9kpZkBnRLXI7pZ9XaqWgwPYPgksATsYqeBr8zi
z3BiKKZwh7cT9ShNzPnwSrI3zMJNC+FkldOjEnmqamX2rpruDRvzBKC3VrCbLwYIKftED19HqTnv
Gx6KDt088lqOe1V05/hzGsR/1QspgjdTfXHmCQtGsHygeyomBM9hjz81vkMUbe9Gv6UCf2cQYuxD
O4x80NBkrf/mWuaspEglNBXAjQzwG7+eHWIPMzmvRrPD9GSeqnsjRTv1ij7rCum9/D1nDontiUtg
Ec0yiA70yzcrFmn6uNbJLLqwajhwPMNZZh+Ihm6goNCwOVKkjN4qE9luNu3+jODL88YusXgJ6gIX
MJS87Th3rjeKtwpiFd44jR3SKrtJJw3D5L7/tmobk3RUKbAwpuWkDwpPjnt/lXDZ0U1Ker7znMip
vKDfBxQn1wkERefegVASNQebhraZwvJEIXPkyVGu01/vMtTBFGylhN8S0d4VacXYHXg8aFG84oh4
bjr0msT495AutuZf9hlrJ/OJB8QLgXztVHGLGG9Qvj9199HxjxCng5jntDcuGwX+1ZU6PLjQvXGY
oVipJpM6jH+IWqkyRKp3G8jtoUFZ5zCFSaVDq866XoTCIVi4Zp0/8zSYa0N1o71mvISuiIGAHb/X
C58DEXv7dlPKrm/QuXhlOZKhNg5NNy29k28Kc8CxuKR6Rsp8cthqdAhZMYZ8c9N4GPejVnIrpD6T
SOjiPJmW/Otl6wbTiPTppKdBTWlvWzdwRKg0z0lnIKs9h5XLINavLDctChSQo7EUlARNcYgU88zM
xr0WPagZqKkyJu0IEm8/C41Q/6lPQyXID5Z58Kfhfe2Ryw6+HHOZEJY8BzaL75avkH9xPqBxsn4W
dvnK51nWDqj6jlYep6M07UpTxHeIiRJRo4bsDlctoYlfyO0jEnqFE2YbVRPtFvcK2foRDyI9BoD9
H4J5vblGZDos5pSt8LdND5zCawJJtTOokjv40ZHc0MuLO1h2NAB586Cb8RaLkePvQWJnoWsR9eEn
mVKGeMtIqQZ9f32RDOM+qR37dxob6klgapHt3CnXhu4zQZEhSgfhplQMfuzLcFDCR7d+8ozFnxtW
j05LXgDXg9C7j7ZSnqCYBavByoK4vhepoZZlc4r+lJ+d0miKEenVQKw7dpQA6F0ab/ENgZjNqF1Y
TD0t1P+Pym0PCjvyYOpNTFJvKKF/+LH0w+2ocz8/F9Av3WNRjqutoXxDlwkL0po3tD5cxoQHRS7k
NY5BS6lqqF/E2Bxs9/jjOOPfUyPN+j5ahbW423Tsy2RsRVv5rYWTacgmKuMnAHTSuXfehGgmH5WU
D6NYVh6ncfWt7Rxwx/A95CG6p3U6K9lhv6nvsxJSeR3ay6XosO4T4RPcneNozkctzw96j+yzr96v
lO0bg48lZO1K5Tr741I+dWyFhENr/dieIg5xWPIQjgxqTuXURaB7JFK187yipmIyIki9f/Kk5xJC
ujKcnxrg1SGh5WROzMxcujRXkCeV8blBTuXreiqH63GvpdO6bbF9ovcSyFiLe7CEE2vPVebNNNAK
pxEjv1KGdGQIeYJ7xrU9+1jWgdpksjfwscGo7kinpRBHY38RlpnuS8WaeGvaGJ8oDpPYPltBrBef
hIY4CEkR50B+EAUks6Y9gk6DJw9m8YdpeJEhlLh1HuvMmuJ2z+LI0oV/II1SlVKISZqrPDNTd5fp
fsM7FGKZfxxvPpvOA/umyo3NeKO5HyOCYng2XHJRyQwZM2PPKuhgmAYQH9GppGOEwAS+rfsfESQl
HqnWIbh/EZPl6IGtBG7RQ3lJD1kCOfRMPSdgpX4rrd1Wm67VYBudV9IwVWvmqtdZvB8vVHigpYDg
bvw0RvknrE2WxE79NNXsosDL8Qz1BCmqLRL9Y3nS05VAJuQb4iDZlPpglq4bIgRfbqTRZk3vKz8D
7sHRn//SFGDIi7bEdFkMfO9iABXKgo4TPPU1tPDbC3ARPttPSG9qXT0Ac1GtpfD6x7rYSN8tROYf
qMb2Fq6+tTErujjazwrV0zcz2Us3sYKDwndXKJFRGijYUgLFFRXWd1qLliR8HUAwi7XINuvgg7no
Egh0ytZkHnPQZklTDMWCRRtAP+qoJAXLQqajdSd0Xmcoyk2kV5dWzri7Lohe4FL0+Bzv9YoChHQD
HzkpROKMA1HRnH8LTVzjmFLqnZVdW8crAURsy8+/+iqzs2CZyhPfaNVP16Sz51cyLD1W+gqgfgXl
UWESTufPRpbBXosoETTKnIzvUJQLHP/5dIvYMUHBO92Am+0HXIuyQc8ScAZAg9ccnLgi6zNEkby/
Kgyjz9EjlBAcLumrjxiGjGGSzU56pn3IdA3tAuDykjTPHdDeCQIwJgvFW962G3UFyHG6ob0Hxlel
VhKfCdOGAbLP98RfoFTu4EoqxZqg7Nz8sewedZBydSsJSgbVJrxO8RnnvniCAt+8pboQAwTWAbhi
mo54soZDR1OZ89lzLZW/8D0ntlxi2tVDkovFMxHnbqilsLBjnk679daTJEQuuSUeyqyltC7PUkde
bKHuv41fcfMHMUS762pPjMZ3X4B64CCykQbHpj+S5DzPmhiOO+KxrHAaHCvk3OxQj2QBV9hcuNN5
Hp7s76Zukp4FAE6a4//EEVj18yJWE8jQ1pFeGsETljjRDduAhv7Zkk3vqMvO9GOLdZ0dvmwvd0Et
MQGyYQh8i3yYvHCF00adMuYhp2HDuGuq/ZTva1TMPDMvmweferLPY2aqrIPXp98nO2hX3940Hczl
8xvzeow6b5kXXi9MmczBAr+tuy8Pz7OGM4xBV5AjVgGELzCeUgsEv889S/cncdWJlHJZ/LYPqas4
YvPol/B0m3S0GtbjcFZ7ytuMCUz8lLz8kojqNgqj7CiF0AHiXkR7ZOl6Xm6/IP+0h+gyi+t97bIn
GgIbEEzkBCbmqKxC/uWmM9sM8DrqPqoMqKn/xbNvunBwqV3G+zGHyXGsTbISV9+r7vaWE7PDB13c
A/aRiVRsc3viXd1tbrNp7FEyRW0/YjXMidKejFXCiUhagKQlE0/rxWqTRvhtwz6VJ590G0MydmNc
/jq2x//mxaMdhYLBYu2gSSbyMggfQMNO7zAfeMfwDyGs85CT1E60CFusMHwwsd9CJRiY8xcsEYeH
mW1UWirao3OKjyX1xTKPR9whMw/UlF+wh5aegjAGjHLPnfFyH0q2Kml8xTe7jAWGpOhXJ0EHBdR7
YW95I04jMUI9DoNus4lrYswhvk4DuTVA0okrDzP0odDMi6Ezrgcni8dSXVdG8GJOs+thEk6/U0SE
rwkfywbHxYcUfbs4ypuyybN0/A1/wGgephQdCoN84hdufUVbUxLHhaHIqNWxQrjT2x5iu+mcpBET
dIc8Xr0xJvsCKIUu46ywDrfjrWFHs2Y07o8f4DbWvkXn27OhVGhP7e0zuq+OCpdI34S0NztLHPBp
2l3KWvmSKN7/fUpipnLIvOlK5VJXcm072qwCxTkrtCJ5vAmjNyLiSdvB6PLzdQsWty1+XEOA0iT2
lMh6f+nKzhAe/1g8WSAkgr8H8mRDIbHUauaniXXPEcfrIxzJhyQGoArTp8B8REv7uvlmm7bq3ahs
xykbiWEjV1ZBiQX5HQ7PG4dJzZ6au0sCY7k+TMdXuhw7CL2jrzY/RtMUaZBqICQqE31q3YvHd8Fp
WID7/jBHtT2D9bSuaJQARIziy0EqxijE4LF0YmVAHX/tDenFOe12zm0PzrOvUP1KY/t9dJs1TvXn
j8vE4m0Zl0hJ9pElGkn2P1MkXyynOT9dZRGC0LZPEgrUGv1yY/9tyFpbm628C+XqcAswKlmPThAS
xzSHLXokVH4ob+gDgmdSM4RiHVDhPO2H2gNXfxhECyWfvE3JP6QgNENKft15KbXNp2tZs2PoWaJ9
X4y65c83rNVU8U/vZJK2FjJXilLXcBKqVOl3CleRkgD3Nh4iQHJPosakpXmGm2XNGHTTHZHseKi7
m5AfopOrcWe/ntc5/ZaV9ZOXmiswjAiQohTfjcaUN5MQteVXGYWDZEGUtueZ99uDHVYYfDaBOZkt
MVayzBB9iOaJbIKWoj5lKKAV0AvUaXL4sysPolvH02pxbztQ0rtZbv4aAd+vrUruLASD1hGhbm27
HJgheBS0L73kQircD9aR2WP3VFuoVMN8l8bof2+YUPYIrp09Q398+FfUMnM4N+LtYeeOTty7vxl2
jN4t444hOfKbCxTX8ClteOWDKlZRjG0smZySrvG/irPR5el2QIDTWEZgAoe54DoJupoEpG0xM0WH
16VPA2KwZvsoXTTHvHFdS4KkLsAMzmyXQwoauAIxWgTPKRq6AvJtWlTRLYt7EYOyzQQ5e7WpQ244
9UchZdocrkYDVjuPbqA8S9N7oHWQAxtjoiX85Kcawz4FaZW1RhJu6d6YVL6DA7KZ3S7cpaLRO/KT
abGI3rFPKskokklPfHMiUYxr9OLKMf58rmaM+XqrE45qG/VUHvOnn48KGWl5bSPEFBT5XFtR0K5u
bxaKXJE4kRMdgxfrFKToccxYK53dwXGX+celbwjAbXfmbeSlJRyJenITOFk8c29UvDxRWtJvDs4i
1jGut2rPg05ZAre2afIJ/gZ3x7UA+MgQ0S3jxIhL+qpvAY9y0fIn4tTV/EEUduNaYGl9ZTODLJ3G
jG7UYp7kQLqA/81mLmKyETVU4907brzfeLyRkcFzX8BxE7qraq/7BKxdUJmZyPVzSZIu/zicityg
3xTrcCZ1qVbMo8GimC6CJ07PpIjgbQpCOXaM0crGurEpEVTFUtfZGkcqa3zoi3KSjx9/SdzOtLri
33TmamW0+R+NN/pZMO+DxPN6njc3launsHHrO+g+9HAHqWT6iWH8IredD6Fhi44tbVZjWCdD48uk
8JNYUOlgS1Wkuy+tqWfsoQkkQureY6ivzEY4VJ4rqQajuXFpWcHP0KVMlX4HM2Zi4dOeIaY12tjC
An6JsuZjOJNyx5ijxivdmuGaEHEsiVYiFZf6TzQc3qbdjX7JY9xEek64TO1zv4KUuY+qxSt0rWkd
eG8cGDRftrxR4cyKQQUDWoD35B3SqExK8zELXZ6QUjTx2iP4N0mK0ypzZRqvEDJou4bctxq2Y8Vf
TMTksc9LM7i3ZxS966AhaPqULNR+S+k9WyiJ0YUTE3IjSWq4DYrU8ryIajJIZQDUw2CpfZratmuH
iwF4+dyy72ynvez56n0WYDksE+9bhE/AxrZUeCeCwehd8c+6GEA43Un+/vHitYVrEY9c9etSaeJJ
Og6XULhzL5XR8llB/cbHtuIO7o5HyWdnYPRcWL/nqV/mGiDfg5Kccw8ZwOGX8x4hKjCw2c9Jel/a
XbYukQZpfZXQyCVnKjVRDX93rQV1emRII8iygUPX932PLLNVCATjl5PVCQ8dKD01AM8yDFZQoWj1
DpURpH55IW9XhQTNgQrn1Ai9dTLiFMumczDyGq1iHGUL4ItHnYM4LbMFifvk22UMPuAZVoHtO/Xf
D+lOHM+/4bHyEmKewLpQF2S6Qo/7q7gyvafMr8xZ4EgdTyxoDazVQXkWBHYhDCItVfBtItCfZjMj
2y5cvngwEKcA2HBMx/5GK4WNDUgFG8kJGMqLOnhSCTtqUrfUkXWD47xLeQupxoqGhc38UJxGjelW
Nhqsps0Jp7tyHYF3dHlpd/bUT2YaQ4mOYnxRPAAqjfI8zdQfJiw15JE42L1J7LpYCW8z+N4yjwEV
QcOlaC4SZVB3m11brQqYxh3sJKFPBKP1ZqGRbLaBRYPFD8xFvHwicQva4RebHYJfYuMwTZI0rnGZ
8cdO6Y836IEaYn5J02OrG075M3LL6h1hjGmHOQ5KFXqKF5k+c8M5jd71w5ccBTg2TS/C0xOd2/vb
otgkPAtcaIJT8uRcD5vw4Q5wgl93Xk5g3gubD1DoGXgcifXmpPOY2DISAe7ud4enrTZnTvMv3Tun
lv2iEeAXsOFzPoCERDrt2rL6PaWAnB288iH5PQ2BXviXufYwTg7R3TDUsxFSU/B4e52hIW7pkpBL
VW8ZwySVu4jYO4UcJDMPHdI1qDumF5L5SBSLmWStpwKHK5IkfGru8oHl5Lw1Anz5pQ22hMbQYPkx
WGqLoXkdzyfc/NEP3KTE1k8M7xtjRntB8QoZvapv0B5fBENb3DDsUtK57qIPRfZgwTQip9ZzXnQR
0sherIeVkcvTUD+fPvcc1XCTb6vqqVtlFJvkl1NIH95AQhoARIZ86kfLm9Kdf6skvGkbTzM5Kaee
BUdgGQC//8cUC2wK1xD0K+H74jYy95hyjsQB4QiZUSEdEAaUiWCGkjobCnjyQpxTKndJplxQoiyc
9pgCR7yaFXwB5evKVDxMUa7/B/TnphueXXIauszwIVhC59+QG9ISe2pHN+6c8fSsAPv81l9Q4zxc
U37SMdFDQUdjMcfR7+OlVEtibnOuoAlwSb1FSNNGTjKaU1yda113rvVQglAGUnwQvAmJWjvcAH9b
OeMk7wU6+ljbgl451v0WDUJNpl4kpGvhYA/SJ3zi5tpANgKE7PL1PIvCBu+IJlqkhRs/9t2j/AY2
q8671/MT3qJZfhAOTlUCm+aVMebxXvA4tJVz4V9Pp6n7NAUqr4Q/AmAfd+iqe6oLmjXQn/Ww7I17
34gSN1GoO0MergWI0MA7oD/KUPyQeSNzYGl/vzTCapqS8Uu68RnFZ3WL3G5ItcUWGLsHfAdbBxgd
/yHqTTwP6iyPEbM69oRUQPoEgfjcY6eg5Tcu/H2/QedpDPVIGvW1+rtDM8/wOtFds1icCM3letzW
rM46W8zWR+23+rBuYJm3bUXk1Hz9Qh+cEnk7H5u0mG+NeuynQYOwZrCQfUMGfP5eaf1cV5YSxIaT
hwMSzBw9eBvpwU0K7ie302hIllx3V1ztUPUwFn+A/+ZXDfJ8ocKeV63+Z9LuafrOybMJzy+Kd7Cb
jfly4jvVlh1cDAiuzdd1iZdD7/FN0S3m039nKi+L7J5F1Z6ulrKH6YDAI6SCQgX/m0okluvbBCrB
uSbe5y6O46Nmj7Jop5SnCPfIpquLiLx0MmWLjQc7qFaM9Aq25GvaCgfNkMxcHZa6ZbgZjuvPC2jW
qYadK0yfo94u8IjH3d1vJwLrbrgeW92bJH91/0n/1ZLg8awJdgbo19MbNDOOVRVsF2NOh8sYXIiM
asnwl4MsN1Ss1g9uHQ3DaujEugCyZjYlsbgHisZqe6WoOHdY3E2r2tfrnvGiQbpDdvMWF+xDVJFm
dApZLJEbWqVI3ABZyEOoytdWDdP303pvfLTEC1wWvCq/JUS7h0WMSJBTfi9CmZI+DkAaoJFCvad+
KOXns0VNaY8gTTQ5MkKdNJcIKX5nZsKI+1ar0mPgxGmaOR2qzu5HX9oL5YomUb0+JVW8MKtx913E
TZTFJQtXaPCDQvbEICF0hKGe6RtxpNjy2BlQPD0nzG5AU28vUf7e9T7bLvAkBZFX4ykQHeQbjT6M
VCvqJD/fCWMuiDZi8mO+L7S17MThw1/+lG4Orp3uZKao5uW0lEBdNZnt1U35I8rr6dshEJekYIYD
eiZYhzW0Iv7oTElDiVE9NG3bS72Ipuyf9YVNosg3w2Wybw7EshEGsYbA20r2s/qwrQChOE23G5ru
+0wZxWLrcS5IrXLPcyF97gnGIqLARjNkFEUpXhll6XyQ4plX6OlTosq2gXhjeFZ7ZAdQRlIlvLOP
PfzrU2mgkkMpSNkUyVtR3kMdD9XqZXwC3lezc1QP1Dm6Rte8eTjOnzHM3FGE0nwL2sGmjveDaXpc
zhdqeomTA50zEHOpK1oCgESipT3hCJLFpaJIt67nVR2Q67s9B7ELaGZeNHxnXSCZuBBmglJmRJw/
iOSGeN7MITM05Z7LA04BJGQWFp0uLxsWDXkrSJSzYHqLGGb3U3HUUL++p8BqCvufSD8Z/D/0BJwO
K53fR9vY2Ukvpym4Z9C8SUt0eQDZjFpsgcVmNFjAbK6mtFPwxchA8HImRBExbhrXxr4lpCH+iloG
FE0VsagMFvdaLWAEwAsAhI8/22wzMslke3bv8Bo3frW6knz1C1udGtNSF5Q3o5PPrBW53/UemHcH
o1RXNnfU+nyRdWiV/zXWp2exmhI1xM2VZ6LHlUQ6iCqD0P1Z5rZ8l/TroQmYi52YxQkYGvz8HI0U
JKkxwv6QvI8YEdztj0WIfk+XvuwHw6tGtfNCTb7z38JYUMf8R9LMH+fyp2C9RRv9DNhRVpxv3pzL
V/5zrIFdzheA+3SZUdcKjPY7yk6nmG7vJexmF3t48tpGtaa50RL7WZerfE6fZPBrsdjDL06LPGE1
7ApnIqH/fwhjNXxTKLGOxQp8oLVN/i0Vz0q3dgQs/+ldrQn4DX5X4irbLvPSbMOSeZ3i2CWn0Niw
5kiAQaX75xNISsLPHRMjWGhGGdr8lxyrbD9btpEjXqofNh64HE7AmEVXfhII7TEHT9HrI4QqZQff
qRT46c0UuyAfS4vATINpagWFolaoFDvUWBv79q+R8UZum3rFuxGC238h2ny036oM/51Uy/xjz5Oc
PojGUgpv13fFR+QALioMQmtg2igchBy7m6zAp3WWwHtje1ECZnmckLfE4cNG309nds7Os9XRSDrC
0tYZRMvzKgdJM+CYitxjXoGvpOJ9GjFtyX6CG2YbMCkEL1JVsfmmUTihW00qUyaKh0pHRKlPhdZ8
YFvYCHCma88GRuWwn9eKL51IHHnXSze2YlOMuBLYTHyuDsoZ7vbWbwatTGXAbF6MNIoxo0NA7i9b
FdWO/8+BUm0mT8mq6X/HLK+a/1tTuLW9Axv2LW0Dkd5q1BqtJAPBqB8/kPpTNnDqEGaCl3vK98dQ
IwCmtZje3OeZf8hTy63YanWUJESho3K8wAZrxStThB6cycxy1luRFe9r0veAZpdeRRusIRl+7fks
GDniwh78VAtdNQhbGeTzGABllmahMW+cIjcW3CAtcuwAaxEIuAOnWZjwOsLUcMfxEYIO7qLQ03JU
7zgaN9KOG1q7j4qrh1MsfxY7rKK42m82Z9JvT3Hq9we7KzPHEARCe96FJ4Ytq+CjAZvQGCX1U/9Q
AbfadGw9pUidCZ8sj9taWrScAJOfSNlXvn4zPN9e7ntI2Pe0lOwdibZgoqJcrUi0BNIauvQjetTM
L5+rXm0Xp5gmHUxk27VqJ+bcdQxaw1W/XzhjfntnOGhSEAiXAN5opgJOP4VK2CobSkdss3ZL6sxe
8JjMiDZ1ZHnYVE5zZ+1fSYJoNkxIXI9kOlIOb4IBsns1rIKW+w2poLeBUSa9wyZM2Ps2F8heXY4i
vRiFccBdcqnjICqLn1/PbWzLjZMKAm9b5G4TebfMqErAfH8X5a8Ybb90z+/6lRvAYzelDW9pcqZb
pOHBr+uKvcES70+x4QJiq7qt6neGStyeRn5h6yX2HHb0ihbBfjeOgI0zwZ/0g4Ue0hWVmsjHupZf
EEGu9u7H8PXCrnDgxhyAzjp9+a/BiyM0T3TFIvt2TrOHcYDDX6UP0oRuub7FCiwsESCebTj2M7t7
sn0SuJcfSO1WeeotgJEwpSamAdPLBuEb21A6nHdVUOE/0dWYoJPiGTPp9tx6hdYz4DWkHFPwsxrc
AcvpNp3zaJwvqIEuXXPXVRXWdJT5tOCDBrHHa0jf7WPf2RgnNmaRGkVvNeFxfuQJjG8iQMxBNjbV
EtMRYJDcfoeH/obJUjrLXOGoIjcDjvnK2viaBc6fRfAUVbKlkgNmy9ytb17sBhnEmbiEfKqQoY3q
KJ9+K1j3Uhbb+vWr7g56V3TeO1vET2HKE8JSZw/aU/TBAV4x74vDLy5H1CXWh5Enh3OZIEHVI0ZD
uVwEFYWfKec4HutBoHUzd2fMQBqxHcnKFBWR/jMX/36xlAfdRrNr9A5SoiePai8//4IWZjTgVPUG
hftVBrIpNe9UPrq49wjHXjbJOlVopDph478M8n/YQEXsYbuszrs2kTMgLI5nOZjF/rkM2vnvYxRV
U9DualOx3vDivWTbCi6POGtY1a/TjWYSmDV0fOq2/wseRxv3JXTdUDuk45vbfxwaOKcWW5et03s6
u6cbV8S0tRQyggJ5NdQ0w96l5QKNLIj6+FNnuyIBebL+ejDU2Zgi0WAQAYg/dagjEq7b+d3Zwo4l
h8k72tyvIU9Pkze0DpRqvAHLzHt4CO5vj3ec5UDwSxq0e8hq6q/iMSSSTZIxbFkRvYzUVu0yOaIH
WLgxaZh9ULrAF2HPj/XojG6AYmttxz2wvEylU3pd/4tDiKAqeD6wxg0AEC4O2aPqSKI9Q56o8oFT
DklrXhar/UBzh1z7RdwAqM3NrG/9HcXsA1IfngSYAiN4BSDxRQDwj/MoEBFcIzO7bpQA1oeuKnKr
zDFbAaGslFMuIhnekNaWjM+tkAOK06JzMtSsmUHZAaGc4/NxcuD9nJXg/roGGLS1CrlDhcvhCEpu
Lq29XbT2zIGNKzGBuhPkN3hjUU6KHRSg+brqdIWvKimiZTvR+73oN/ise7+vMafdXozbKZ/k0xjz
iM3Ozk+n7xWjnJAW3E3FEm9dImgcsES7ymNYYJAoh6vHzM79KD/mjMtFp/F/o7Cx9G954U6lzXwx
dFCYUrMcUWGDzVW5AN89uYZxTT1Ly3wwml9ux887wo4X5i5jEgRHaurBMiOUcS/Ej8aDeCdcEA8K
2za0NneZ8RUPK4sFEKr1Q9zEiJXfHVb70mZq86mXOT5NMUfcxRJQ1HcHiGv2gPGq+12KjyU0HNej
Ofo9JcwIrrH2WvHKY9s6K6hhsA85m9LZw+503zDPfNH515SySiDV0GzWqaB/1+QXTJO/wEywi+R4
Lkak6HmwLTz4lUuajLVS9SaLbHvD8F2rRnpu1qSMoascrJKEyKQ66I4zJstehW/v07uiVFTLJSD8
nxLACALU+xXEM7IMRZX3P69GUsdLTNThoHfNnSmxp7N99zYXZQPD+8NW2Pqx6rOIGLBMXtQ5FFEl
7TgOGbS95286FDop6Ot41vPEn6IQfmq7wAM3u7hZtyJzEpgMkjJcFLSItfKCWcLleiBGy7qiTjfb
pSiZ4R5K3JZFCURcsZyxIK1+p/5L4Kr6zTRVhK365kuNT12pT3hmnDYtgXDZKAfnJ7gvxA52dVo4
+x+S3b65ZhRA3kYP3avVLPITFH1hrVugNfDI6QT4ZZk2uOyla/h7avaSouK+fznKo+x0mmAIjYED
c6kV2LGP2qU4i+fZKU0tAfLCFAVDIfzEFoFG8vGAdlIJH7VuIA/h65Ir8r9MTxbik1SXLpC/+6L7
wf44nt2pvy0M+evtI0mliaOCTeurlU9WyBxiRYumPv3PzseuB2gQP/VgVx3SKi8PGFI0rPB244yV
iHHTK1fBEoHWVueO4PQiNkZiu5nHfdTAqrw0xx22nIsoRC9e1Tr/luXvQrsIbQuneCs4XRjcnODh
x9ZjBP6UnfMOA0nexvOz719/CSw3tgXCayDbFW3E7QxkTalGiP6dBGrEn8As5mdP5zGE/TnHJtPo
57sOv7XgIV8ILwveltGUtcwfn5C8q5lNFe1LHtyPmFOJn3olQw5XS7AwoZaYRMLxYvJ5kpndaTEd
JnZJnHdQsHj+kRXiAPAuY69IIYZIqo+CZUHdHyYEzd8smrW+/VsD7NwolV0bYDb52nhkL2KfY8xo
MNw0O21pc1WqUUGNxzfQ3BMe7gsBTIxIaFbr9/lHqOVf4DyUgbqCggEAX/rnwDCiUjaDZMWwgIO7
KkWWHrrS10Hu2T9t2bFA0kxmSvyw45F1CTmE46IJLBcxXb0s/17WpFAQBoX444xSovptdMQ/Zz2B
OIKcaEOhqD2CcQXydvzazZAhcFdcqhmjnh80GV5BdZ0aanpznanAdAepxkzEveUGeaKFEA7MVFLo
wwBp2DKeOLT5pPQrVhILBIskwEOB783QyI4yzUeqWYzS2hwWX93Ytc5BqlrxUS/17+krT3xU496w
LuRSRiimX5FPvXz4PP4AnVr1dg9sYjJUuumx/KP2T04eDYzPRsMEZ/NxprWttr6ZHRpfNdlq2WsN
OV3NbM0Pt4UqU486O1/VIkm5vawNLe550WpMbd79Ou7cJEI17mKquQDf4vr3WsuWgppy9rU7XapE
8oz+cpUyIqVz5sTgjR57JXZMuD0YKCoXmios2Wd6R++PQV5rwipBoS7LO/h/0DnTOutPNIgwtEV6
qqGnYSByWqnsYMEMsjzXm5F+0uBNl/uFBNTRpBhMVAempIuzWLnp3xxR/paE49Pp1InDQXKH64oI
H58zlMMblzlU6vgJzwzZL88VUa5MM2e+CILm/4q4QRbP8l0GrrLLdi1YJvYf5wzbrmCSLoz1JegF
g8u9jVt3tTq1GMzthiXQ8fYC+sSzOsZXFUlMlXgBM+VNSUYl4/FfQSrZO9CfLdZ+BBAb7JCRJLV/
xQJpoC/bWK+3vsmTQvrTcQoZP17KvxGDKVXVNSfys8WxFqJXli3DXD6HOh/zMlpihVAdPE/a2Pba
naQqSjQoyTZv5STDm346HPE3QBxddgJwqKfCqT3N2MVb+6V0ld05p0UQG0zmq6HCCPgYNaXnOZop
xClXsc1P5TbHIYMqEMdt6baWE0G0dWDhw1VktUxfvMwlm/YcLyy6OR5EOpb/MrUF4AO3XaL4KzyE
9a6VEkmDMub86L3kc654KIDRtvYAbCYQsYYWIiUb5yWrvOym7oXbntp5QK6FNIij0plGZLdCrxL5
y/lD8uKWcwS8ys48Ty+2cVnYZR4jajvfyUxbekY0OqSC/5/nIC7BKextu3eJVZU4rwDxhpi8F0yT
Hoe+pZjQeBzaauD43DWzOjOfrRtBzRz6CLSg1gtkCWK9Nyw4+amtQp5a5YZWugaWwuFxuDE9v2Wi
FX+uBwRKXmitWkqt2W6eJFwjQ7ohw9cGlQwcweXaCqNuQ9B5nQHttlyvwGlwwS01YdaaCbcx02nv
Fm9a5izj2yCTqcX/WthRrsgmY65WKUtt2fhGddWzNrAdzWfh26I9UMN0sSntbHwLgLysdmmDJuCl
kO1ksY7F/2RcNuX6KPiEjaGioCd2tXw2T6zB9ZIUFEoAwmHr/oZ+dolEsVGGmKcQhJ+1sBvUtJXw
HNcRC04JksWLkFOvIZsZ1CmZ/I5faGfX+yP4IFRdixbxyrp0wNY/ATdRbU4jS6QRgLmpMWm9ZsgT
85OzGLArqIIJ9mz/0mvg3nkJhuDexWyzxF5Vqow5xZ5UzpA18ePyChTgfSylDxDsHVETBQaDyQ0o
Y5fNU9kEyRm16XiD/1uaKbNvVI34mnNoqFAimaRInch36S2vOETZM0dgUBJtNdiMk75o35WLQkwW
MBZeiHgYHOx5GN8SGCZNbBkHelUaTht1fwmy7r3DOCugYpFiRxocrKJLBL727lU8qDMhfGXd54Wd
TLcSqmcfAF8MG3H4BgSUCaaZlyL2xlaXKRhxOYceYSkTblxKxks4aTsIgcY3A3uGc0u5GKctfJId
boYuIvskQyYXtOUxp1lDp91aS6f4uQT2a+/6smQbVTTVmdshHxlalZKdbNcSr/tWCpQ3ccKCwTrm
+nXIStUAc+FsyzR2QItl9gvUhRfALTazqr4euwtYPMu5IhzxBu7danklPsFuStny01e8N8q5aV9y
Fev+cD6LRzZGf17OKFKrMMhUi9DsfsA87bAcSU2mdTNbguu4ua7YWhzGEDkLz8v2bvgjVgPYi+m6
5bzwX90PlJ0hHHvbYkYPm3GUBWhJgVAw394zUXtS0o+uwZWxBDl5ln+WlReCUOGnr2sz3Vr9V7JT
ncH5sfy4GRZIXG3WF9ade9XDFRjkXgy9sjUJH/yU44zNX4JTpBkvjgjivg5P3RjHZAfAnKlsIN44
Q0IEo4ptYiDAiBWL+7UjZkDESJ9pwKY+6ixsN79WrsTutW4S1/TmMX5nbOhZ5COtxEnbxZRVL32Y
TKB9KO4A9sg93Wws5GzjrAnMCTIlpFlXjj//ECuNIPGIR8VKv3lqpXpU19Lj3tYJNYS5s4jAgc/T
KYS3ub9hTOIIqF8KUkIRz4H4FvO9WjeLx16IdDAAG93YUzSfo6E4m9KYiJ2xLkOO0H05UK7Wj8xq
S9TiC5oie0vGeXYLir48UlswgEPcyLhhjHzYX4lVl+9EHF1pVNn+RUF+jOUK7auiWZQwLHxgn2nn
Uh5WJ8W86tOFZVk2Kjhlrwi/bsqhhCeYuEKeo/1r4MypbKw/LNgVyLclTHiQafjPbTthzdoREGiF
G+Yyh944cG2dqr7aTSLuauRXKAdQlYOSNCyXDeNYM3vkLoQ1ifofa80so21MKPSCazH7aebF/YoB
2+mX+ZGZC6A+ZEwFEmBQra6GB13PLJWGGi3KBLbt8t3me2YzQNdK2kc2AajTANi8lrQ6x8b4FqT2
YZgOMm25roFWoSvcjgWLEBpvxtoMtfwPmcyZWqAK7QlewEgoq5t/VsIz4hsxJEkC1TbA5AjBSLOT
UEUfYPV1EcO4duc4/IFWFgPsv0u6O+WBr+wZ5rmiw4LVn3fSIBNyVObSCJr1QObAosKty0kMBtSt
Wg7L8nwyZeZcG5puVEX4yqYFE2dyrk6fEE7+Oi51WZJmwJai7F87SKQiEeWkhqhXZm2fR2dJFN0U
+cgVHveuc2qa1ZZyB8j+haJMkuy0e27ZgKOz7CiTbDN+PE5amoMRuoaNQxcwrnF0xniXK0iLi/ud
HoOfdI+uQFA6dAQIkMdrcgGt6cJdavk0otHveApS6U8z/mycsqL4JuVHDKGzXk7SnAGcV0akZkdE
/K2HdKsOdarlV0m3K+HaQepMCk34wjoN8KD/tAWmCTsvyosy/H7pinGnoWogDGTQs5VWh7dpfrh9
gV4+6ZQ/+WM9aXHXhP8uWLAsFZqkghhH61aD/Vz5tnPnzXOt/bIv/Sc8nKdgTm0/KKfzfsxZCeFa
Yzt650q+nklTgZbYLjek83Cac0n3oPmQ7O1ggNGg3297HRHDQo7bULzwqkk7rPU1aSdIPijrHXKZ
r3POfzrgYXA5TAa/Nj2dbRvMPDMdK+x8LghTPHfeswSMKEaIEBkcKTMlKuAFBg+A6vi8sojK48Yl
gRbGw7D9d8Cf81QghbJDb33OOaz/P7zBFgzS1cvircdqkqYDH/y9xCsrIsxH0Vm7Nb3gTBnSl9ET
rUBM8MFcbPO33yAfXn2/50FfsoP3BECKMKXxwM5Z+yO6zauPRQMckcDAdCUstQTocaYLZF1g9Pjq
tBoaeyeMd9JEZvwdBiIMnNJdlWJCP0ygo+Xm5lfbv6cmmSRsF6L0p2EoT9LLTZNPPD4SJ/r6Aar6
3AOu2UPBO8OPiVKZTiDDra/pZnqcm4c8JVgBNf4oAGAK/ykX5QrEoHoVHgDoB+Foh5586huyxs0w
1ZMl9R5o/8PDSI5QTKxbCPrtibs/7BRPiVClR+kXd3L6sXDqsynQ3VAttDgAgmYcD0bEdISGSxcn
v+GQshK0khRXgm2Z7WLzd5IoeuH2LPDmDiyxbUlBJkHYEuP+aUGvOrDPaYSgQSy4bwb++fJJi9On
w9jHNcnggbjd+00PW50PidyzArMdgo4wkIwYAn+8wUW+dYF759qyspZdKN7KMCTIrV2yrHoEbGym
b87YjygJVl5yBafgC6ZfCwyqykFSf8qTAXDArEcR4CvG4IcT+TPRAHPyvy78mtMsaYTTXbySmN+D
0x+s/zi9Az5BEJiKdtlI/yUCdtMvAtMWQ3Xv1sDYLm4Yd/GeT/tzm42sETjgNNiADleq/2cfiard
9OMnuJaL3ccmk603gCSMagsF5aTQSRpvkt9gjbTnJ6/Gl/RvAROFLye/JjrYlqsQZV0vHu10Oq5R
44p3E34RD32cCqpotVZYaBE77FmJcChXIq84N60BTcjXlnl6UVeGrD0TDFls2bjbmP0vrwsK41fJ
cl1SdDwNaFV4ewWTOAGUj8yLD9Ret6Yd5yCSktPZ/iIf+ME1OS0iONjzpUW5UOvevBN9vdbWqBo/
gDzl8ISskLS9erYmCzADfU8qkGhh4w4ijYoubruPlrTiKHAtGAmiLikpSQ2hI0rFmSvPiM+cezC7
4s5/1FajcUWAZZiwiTwO9ZtRfwIXbeU83PxQfkoGvlSf8/BRlhnV1mm/lhqdlXSDC6TeQ5+92KQD
FG+1qQuDuuhklFrADsXmYtsVR2QbtnIleZVWqm0fq66/mtWOv0FJcABveQdM46kiYd0CDFIYFW4C
W1WLG5L3aSTHgFJEnh2Xyy16gwaW4OQ8YF2rFPkWGgawBsY7d2y2DepOO/t2FJ9oE4lZny43Qqvr
PFE3Tb/4IYSG/tj5NVC3gsfMjT08AyGqNNJyQh3BXPDsx93opLN2R/cutRXkkOmMd6GJQwtF/S2W
rfg+XsbuuLBGaGFJPyGgew92B0hciIvqn84VEMbwJknFVnrrOL2VPe+CK7Zen1EfPwODWyOnTGJT
2x1bBErZLTeO/myCIVLiGF/9UbLab1/uFN2t3QykDE4UM/GtprMgMRN19wXd3hEhclk0AuuCqXTh
XVbn6qFkIjjoIW3NL3qSgzgZBymgxsF5SQYSOhAYV4uOtd3njJb2d98Ipg6kMw8Zq/h1yAr0k9g+
VrfZF+I4bqhtwAtDD8Y0QBxtjimSYwfIktlVdm6xddGBZgalKehd/YtIIuIdvxMLr1zO/gS9StNw
sJQeyxAh8h71GpQ60Z6oyzNvOeX067QWmMEvYb7DROkCNIZQUyuFAlOvb1lDx1knNH4yd2WaZK8r
r+CkmikoRvzvI4eU/o+jOsvVFSWgrydlGdapIL99qPTQneQcc611Oon/Ab3JGfqeMX1ao+o06umh
8vZGBYpMgKlvfN3niid4OiEjPn24owe4P/wf0BcEtzsUH7lWsUWB94z498es+fxDQnuoDh/nY4gE
ajogxrVEIHqfTctwuMob0UDFrvsIzKwQf41Lv1n0nRBcPxJLM5UJ4FJlZIFS2RYIJdrd7gF+hih8
YTOjIoV2JrfBdD0xK//SdmI0GUXHf8DOIxI5kGMsMA2C3TGy4lOGqx/ul4Vad3YQV9RCGKNSBSmP
swelcc76ZHQsfBv+R3E3Qhj5zVjf/K6AoZcuRmOR8oDZH3kuE+SAguAzah/7ESvKGl/2j2XOqDzR
8iiw4nialt0pWtCS6tkAYDgNFRgBuQ3JSTGYVBXjfuzTxw2isrqagSJPHE99MTW5AL6pXUJymVgE
5paNBZsADMcR1hyMFUpH7GPeGsBLRgE/AKMgA2GARIoaY0qLY7Q2ngQkpZxzDK+JTkB2d9bPAKqB
xP//3NfAVyngOJmT505S7l2pkRJA3zrYI5j1lANxGFxyNlWR9ZV+jIsmSRw08iQNYJKeIVFvFn5l
1qGHvHHovG+z6dzxC01rj9zFwVtlh+QuGUZJ44LULZ8d9NIxqFBTw6hzTFEuL46TS4KITWMTa2iG
iawcNB64KNCr/hxLVwfmEPiO7V96PBbe96vC5j6ZdJ9pZkuDE6tWqujrPd9sPbGbOKfqfCMu1lqr
gnQGK2zc+8TwEh7mbOGCbkbR8rdZ+ejP/5kyj5vlz/VpfsT3EioUydZUsNTWnKPuMXaHjUC3y2/b
GmPmlTvqKIvOTpMd1gLCqFjYWWqhpTrAlg0gDtNHHujuUhV37JUpOgQyqvu2yfL0ys1KBhX+KKzc
fwwwsbhs1XqR56X2EuKNYJNJlfGn0h4d68iUsAfHFhWSxteq/l50Xe9B75wleo0rPLXaLl0cZ4/D
+TtblDQbPjt5GD6CqdaoLwzNDp7sbMuVyDrKgABFbLepWep5iWe3Gx/9AEaAD+qIz0TQtdMLG3Xt
s56GGUY7kKfin1p9z+rCo/yd0eak92VLYq1YxTUoSy/7gKhZBLIovInn1DYeF2RcZSBCqIdzpQJ+
98rQYHmzURIhcv+960/FqHzeLpfZn/4+jZ+K0qq++ARWl56UCMS/tsJWH18ASjhi3yXtTN/dMk8p
hr363JRUnazoPzjnW+sZCU0jaw7fLxTzW6MNxyBoD+X/7zjjs2QTAfKiYAfG04VO3HS8raJF/m49
XxPD/s+Yn+z9K8/o3QiY/hQ2Owp6xlB73PLx/Ldb/KPzdc7AsBfkkQr3xJraAEhegTtvnN8n6oXO
vRF3Rv82uX3wiPSBbdaYW9949zkFf3UcjE8vnGI7jymx5eK+9sj/L/mOK4+TluKQDEqo6yIHAnq0
GhXokouz+YH/biv/1C3pYYmZtYMP46TSbHeTg9Lhu/ryEUFxRs9tGTXErY0InTDpXqBpQf9mHK6P
2jF7bW0saKO+hhkzIRYnsVhMC41X+i1uG0CBOfDFgVwiXx1PXdcUY3Ez4N4DDDaZZ8lgUhbTvAyQ
vaX8ZCRa6AUOrcqYzmY0xNkF2vkalIbqfrKwMkpYQOB+740RvNloTG/JSkfhyn4cBdhsahtu91ea
NNcFiukrOsYLZKcNdJ45Mw2NjqFrOf/v4RBHpRrZh9lgJn/7ua1KojRK9Shb/LC1mdgBwm4ut5qC
IbuNjzS9FRojFqDP03lRHGq2/iEdHIVGJGJ08AW1CU1R+RE/psouENV28DWBBZTGfc97O0HqTwnW
mmdM9wjCsukKN2qX0U6w7ELJHDTzEcQ5PcP6FZVEVoF/J4LzSwcN/07lodkHJjQVOBy09bSBymwP
QIi03OlXCj6VclHKBXXmuRLluQ5iYY+6KbY1FV8ra1GBaJKT0AOSlGoamYWc8oO6xCHOKG7sGpeF
8wCJMwwQ8RJ7jyvvcot+FtgRD22B1nO1yYoWSlyaYksIIDvyyJhSaUOyZcQY4nvJh4mgvZq9WZd9
MPAFAVLirpMKVk06BhngHG87iAJIS4VLaGq4T142hdx6ELiOJ9khhoKcF3yNDGZBnvbwk+gu7J6M
Pb/65XDtDlI12Cnzk5bMFf/GQLhNv6s6MLKvmxj6J5L6KuSr+q/BDVn++YqfxqNImu3kEBDwVBuH
Dd3NiFcUx767NF70AigpY2oH0AC1ZlEq/SGw5vX1bsCM7QfGyshRT9Sc6NBeE/hsEPYj7ILxy4Ms
NDFqF8UK8Xz2RAFmlDgidkRzc+8TGyiT/micX2rDw8NJHyKQcgHDOitN4jL3dPvwmmpcrpckFLGQ
fH1WLGzW9XDZt9DvTmixYAMDT9v2pQiljs3DP8jv6K8yG8SEK/knm6eGOCKXIK3Nbrz31rA0RMjQ
hXPUP6pXE2X0ip4wyYPH+mZVWJbfCum6iggLnX0+IlHo1eSy62FretQ1DKarwuuBIDwT5TFv3o2I
b9wLS7pSHXvZ1Ezg4YlR0fwpS6NGbJUqya1KAEEFau4X5/julyKFyZik8Ymji16aK+ZFB2Q0SkvU
x4TZk7vbIW5+fQaNMU5aZ40/8jjF9mHUwLdb+wbhYbiPCifDEpf8HpUin95IbDmOeUgVLwSMQCg2
if98VusA6LtGOrR6gRvGyr1fgVGJKq5faC7rEWJQfjjoA0dfwUP8VtFCtYNdF9uyCSOUGW3JgHia
QB+aEgcH3S/CsD2251pJYmuUqcJl/UQ3pmj/HoRRHPA8YurEr4364AJZbu9d1W4Ngzhej4Rk1E8j
YFELlaWcBJQBz70sR1QSHA5icHPAc7NNhdfD6kg6v6vdizL1Ke9Fg9E3GciCp08XdjNSQyzJW7ew
1mk/IoOn9NCX4Pg2XFLSni+Ar0wGZjnOvHIYafxt5Qu4JADtchbzzQT22asOMpAP8IGbBtuj4ZCL
cPZq19fb6qMemofTQ5dyIfyjSk7oNXijwYi9+CkefHNgDugJjjyPRepN37jTWB+FmEI8rUp3dmWo
4IoutAZtR3C625LS5AVO41NccTRl7bIKfcgIQGVahZr+JsFfLwdIcqxkKLW2Mt0Z1jQx3NhHuKQS
sDbI5XD32gZV9gbCGPv95bxaSxAVdv4eAleBlRI5BdTEwbAwJ8m31S+CgjozBpbs6lOFoDzk3g5A
IjRZI8Mp9sY8SVmcTUwblKuekhm+o/ODtJJIVGBfRvkybWQnDHJeAAYxOD2Lgh7M9j/CKkbQ1OmK
OC1N5TpOtydid7c/9ZAHGVCiIN8JTudylhGjGn9ERrx4JhCzUOJLe63zxITy1xMtts/RFemLoxBr
nYv5XvOJyu/5uvEdGBNUhY9WRI4FgpipMyylbYBAF3N20V70+iRd+Q4+5+lCxVOmlQkZUij77akB
ABXy6j4ZZRGkBaKgR32JmNp/okgYZC+96nxKgXqEXtXi1XwuFQO1haQxACKKf97haV7Kae2scOAe
Fh6CExqPzulF0Q0bfPTAOJuQa5qW0w67nTGCGnMNDMDYWJp+m4ML/cW0NjW/Hq0jyLs1i/PlbI2B
RlNqvhHtm7Nf93SbAmMj2yJZt/PK9EmA6ptvUNT+gicCys1zgPwlBrQU0Ttrb6NWoz5g3MT7abQ1
J+m7lUINAvzuO+BD0ZYFq8ZNa1SkKsmSJNjYBuYhWKjps8QFiUdIEsO4iFIxbooy1VUZQsmEmKLX
AQ1zMiGShfkA4GG0txsMrh9kh2w5BNnhxBtYg49nVPhBUaEa/e5eSNGTnWn0ih/A4Nj3DEtEHqvz
XFVfyejf1DmWbm7tHWc/hiMqDPVpdFrhpamF7OpD1mGp1cQY0Aou+K92toeAPD/5vwv5vWXC7xqb
BpTEXNjQJOMGWgXFniKJBeshlyMVolIP26ykx++RNTVYL+P3iTP/NYj0NeRhnivuAj1NL6k+M4tP
QnJHMwyD3/Ql/VL1Q988nbUAvvl7KiUe7BUPnmM6zNNFN1WR/2Dq8Vb+CQmRcMqEeyUHoquZFvfy
NbzqWK0m827cNsLwg/yxJAcBGBdYMWlYrePboHA150SVw92dt+HVxKh3vHolm3nQzruSaFjLhRrj
EgKQ7Cj70/6UVKkL5semU8AryIWsCmHge91+vlVchPPfh7oMmIXThB1306ScRs8qIkIPniFxSC6w
2mEvdsaiE3t5hGRJb6SUYuBfY7nJ+0B+GKEdUFuEi1lQAoQxaFJdzoO4NAqKZUZsq/jbViOHFpZP
g0Yp+WPjoKX2lwMfTpsh1N5HXy31VgZFz0Ueyh+kn8F/64bkK/cAd9tACAneVPmQepcziLxLSvLw
GZVuI7XclR3qicvG5zRgDlwM4edo36/mKE538dI/sMPSon9qcHt2VAAUbk8PRh3uWm8fH2zxrFbm
EmsYx4BrQB9KV6hronzkqqvkUVZSi5I/BI35PJ5VRMZ9PMLn0QpKLb81iCpnELmbAy/cBvLzQmVR
ngDcyCnjJo1jqpIBkqYd41YVfffD9+w06qZnEalyRzCQEDw2Enze47ZJQRDN6oF7fTTpeQhbespp
CIejKcYNCGZRUUXEWiN3viM5vHCDqncmBj/9VxQeyPfjFL5HlK90Oy1vtrcjxvWoAsTxfzCEm7aA
a70qytqehAOOtTbmOMunrJ+3YgqMsq78Dwfbw0ONDrEiuSh0EftOdwyS2vqrdn+A6rpuKZbMZSfz
vP9gh3UPDi9x7rcclNyKQYhvvMCE+2sAd7gN5lOLe2B7OhfI1IqDdYv+7SwN70ZE7kKmYG++qUUy
YPbljlzinfsg8ayoe3rVhE9UJoX0rKoUTFBxY2rN1H54dCl0rki75ZKGwXoM3i/sKf068mpy9ofA
fJgGMQLKU+SrjNurTlRgQiPiaIwHf7CjK7RK3IGkMPWz2tXvXhQmCI7qXSVF9hWx9La6K7Ut9bf+
awIvWVT3e5ZoOob4A+liOvuFIhyU1IUpoK6gPeKBRTVuf+T0Qs3zdd6GPcML2GqEZWsRmaf5NYsU
mKvY+pXMYzssGTL54c+cpjgaYfcqPB/aWip2G8v1/Sntgi90pm3025Ahba85I5Q/VIvTx7qFjTKS
cZFv8d/TAcQAbym0njWDHBJP3AsSqp/fuqDySba7wsG/kBq8VUCOGV+EQ1I3JTqbGpcvKDQvBWnU
u2FEzOkFM9LF4uwL2KDkYtLqa69kKZhEoD7BdKxwBcJEyJqMNwSP03edYXqzmvGAmUeg079h0BMr
B7E2SdcBRIKd9ql3ZNzNjvYJZNDvNnfytllkLYii3Q8qUgoRL9nvtUOarCxHJ1w1s7WwMoer01Py
L6AwzNUPDjeNet2E4q0L1D23JLusiRQk4DDYqeb/wTPcsLkKfkN9r51JL0WJB06rPQIGFvSZl/vc
do9A8CbBIx15IMzRUnjdOeHFTHS7vtxBFMYyyaTDflbjYIIFQg6csG2nPa78gqBCGAKTPNQABdxI
oncAYCsUmyC3tZ9qN6RXEM3cOi7ttCnWuC87yo8katcs1uBelK5PfQ2B/LL8rFxCNAlZUDMuUqEz
yzjfCMOiyFB7kYj04QUsg/4viDxrYU+rQnT2UfL8VRIx9CNOORJP5/HdJHdNZ5tmVJ+80bUw6fiC
t/TFxwmEz3agivlEOsAYBnCwJRQtuN/PsUo4zRdRTUGjUlhpCsqf/w4FGl9qqtaVEUDGs2v63aem
4FhX88EPrZV4/zAu4CNKYNEVbUVP0HuYSLlw3S+vcWVEIfZIchbFst/RjLUH+Q51g7RxUoFSrTwD
u3URUpnaFJ8QFzUPN5cX5Vzlz6oh/9Z50yLd7mvecTKvJF1YilYddw4FNXSRkPKX6ZQls/nOtn6j
jKGqAhGRSeWD/wpgz8AaZz//k//kvh17e+6GolVg2JRgjOtkbqLEf+I6sR9BbwEBqVS/hocJjQUQ
JAqKKRXi3g+tZiMJB6nbmR6K3yleTHGccMolIaVLZH/d99xNjgMOZ29pWDTNjOgX9w9UmobbjSdG
jvPr7O8z2gaWFRlgcaUdt4Vtrw5LDly67o551/5hOm6c/UPgBurbW86XOnQLR4r450tVSEsj/w0x
PKpqHOuA+nz/uqm2SPtbNEgi7DSO45tXPfebtEV1uku6qpI5ABvey7ob45+2FJhaCca0eCMV/2tb
E1rTrxZUtUKuGxI7Q2vXCQd+dt0OfaATVUOXFahL1kBmRlSW9M1bdsyhgn9sVZWK//8OV1qli0Qh
sC0zosAWXq2515iL25OKEWgqmcd/vUm3tXNLqg+W6OpE0B2IrdnZmTI02vwR2zGKhzvhT6n+yYx2
G57VvhlCv5gZ9VwC8hY5CNA0sYgdAAzOCqrS0LzkgKbXQ1Nhx5ntXMGaHtUS5jJtES60+Tk8avRl
Wwuv52VKGasaKkSbs94/uyRzPj9HWojl0Ab0mOYqtrI6EcinRLiHF2LJo7uzETjHd91aP/JRo8MT
5RZOf45W81PQAKfi7+0MQUzJ1O+dDTTeR7EHk5+Vmfx/0WjV2OBUny/vS5zlzkaQzmQbtfePxDht
RPN/+VwW/XxDW+/6IbHHPMxwsYwyJWQZVvt2Oukj9JuVOaukuED90S/KBYdIXbiGweYbLw7k2KG6
cfE1XkyGXQoup/yViOW6vXh42tFWkJrUHSWtqaN4s3Y2CmbgWosBQ6ZyTavmLbCq4r1e5rCMZPZs
CgP1WWRPw20h2MUz1Y9Dup9HS30x/dFPg9VNGrutlb0xf9jNc6MgSW4fmiSMJFLxHGxaqe7v6h8N
xtM9748y8Hjgax2z7IdSJPf3i00p1JRD6dNBXBdI9+FeYoKu5XWIvJ2zJNE6+F5zCRpze92hka3Z
80Jz3d10iLqu5URwhbFIYuJPqh4UJxRlomjNYDLXvYAZYvqnvT5+XuV1UfgWMUqwD/Z/ZcTg1fbe
NPf9AlnKg5D1FTuOGbRRmOGQj9rX85Vu3olusEFbNN+VvfoujTWUqjRaIbcRdbDJrLlbBNzynBtd
TfpgZ6fmSOaRVVYonpEVeK5D4fbfdRwl3xO2fm45SByxoZTcYztoWyFkK4t6VoYDJ4Jv0WE4rAiN
lhCBCrx2k/ROjp0GncvWPihlhQJuL23uGP9HZilkf6Z1fOoM4vQ4gQaJY9weuKVuL3PnrVf01KbD
BO6S3x7d2kDO690UKd6h2RgxTbC/qh3hljSQxGf7YB44LEp7V7WHbGguWk1NlB4osjLTcbU6DQQ8
h/Fx2bWsgEJXWdGjJLv9CK55k4q4VdfkBH6ZqNYMBpz8At9L5f/J1May3BFHhCuQBnulafnChy8s
jYJorwQd2mLSIxJgyN3m236BYjb9BYFIGvc3Y1nlaIrDTRhFD8K9ZPVR/vVaF8xuBkw0Uta2LEn8
shPItqJNVwuHzRg+JxjjUt6iCfxXlykS+uIz7il9yBSinjIeQrVcOsXfJ48G3egLNFAEjTVlBMgR
DSVBJifBVoGR5xXhXlkK0B6mtUMueAvYRYuxBNTHZ34461OIJj3h9UU4HtXX4hKMu08TH+tfXGfT
ecztcAZFKqhAR1axvazM+OKuoPeA4PNJnGhpdlXe2MmKyd2gs0yzwDdzk8HPKOn3Q7CwLKv5C7da
1gN3oNWJ4k1whneKqjtZx61D5tiPCxq9wlK/3DWmbyuy27zA2ymVgv/2G1LUiK9NiG8auYPbd1Cq
ifnniUfag9ZIXvh/wfpNwZnC6YE0i/k2SMZ4fD0IL9nam1ZwBVy88AFe0ngk/N5MNccD00xONIKn
1i0FSzck8tzBZHI4loa8igSPMsRJFUtOU/pOJyA81cDSRzOeSQs2rxds4ZAIqD8BYhHbuqJ5VRUH
jaOLHQGZb0JX+bkQ1KQlQCwXjlpncUjPXCYULPvgUl9tWfs79KgMSdVceOF8Go2hCFtZVvGe2lB6
Ul+Z3yLmr6Rt4+NplGCi5cj8D8LTHrYS9F50YltiuqV1jmt8pOE28C4229NlBsg5/1OVZTZTI4hZ
7lizpeWV89wJOPE1RTkAXjhEc5suO1P0AuQFXA/p8PrwAHJTd8My31haD1lHlTrPZ7mKYs14mRjq
PMUyU6MDim8AJqlMBS+mMYm/INGuWqmIu9vDjDVT2FUNm0Y2IeCyWUMZzgHTvxjnory5L5QDYnRv
GcuEplrVKo69gwPRycLGiTAiq532wfndwp4On9ZccmL/pFZA2zHbx0yJNe7npHFSRX6g6GLD2v78
XWLIkoigV0U9ggzCncZo7j/JJcBc3tWeKuPG3sOT1KHEkkClbGPoFOvo4jhDG1BY4D606udd/aLT
1ZRUgXlFtjB3c1isBaQxBg0d9qwbD9hHJtGGNvWGBs54OZUM5KE44+pob6ibI2WrP/qhRJvKsfv9
ukfTYEE7xFyc3xHXaDb10OJA3Lime3h56UcKYAEMZK1QHz95LEP5rthsI6SXcmmxlkaMNmaW8OFH
V4kzQ6VCsgL+0awpNcu8YZd3h3ZuKnNdpOsqT5tVnyKIAo+dGHPedplFMmR3ktYGNsiVBjmDyxBk
eB/5B6VIHLlOo8cAaLUr4FHT+ErwAaS1rwU4YHVq2a48f8jrQTSLj50zSKAalyQfNdQTHKjgrbss
VPFKwbxdhb2r0jho07USQnYakKNjEEsDILGm8QI9G3Tc0zArsDRL11OKD7RhuvU/fzPicIMunvxD
34jfrdOhkYEsZ1h0TT0oWYOjtCqRcOBMghJ4juiqRSl94/fqQFLMtHSFQa6hfEnOdDRLVAJz0BHW
0VA88f7S7kg35dUmFPzS5d2peLL9oBOVgDOcCQcTVJXDxmjw90yeBzttGlsqyVEFr3EhpL5Ei0hy
NKJpGuWvsNjcRTXKmVmYXAhrz9cyx7NqShPTc/+Dyhjr/wMa/9bixyZ4qe2s/FjsXWz1+I/b64jE
uHSpL/YjP7KRo6hyZHwMGw2VrebirBJvzpvTztWyckT0uW+F/74qqEx66q2Op5aY6pBvoS/yUoPc
DTdfUzlr34hxxtl1jAaT8AnSVVeaTgFrOyp7afJYbW19t3ocqunrVhS00V8qdvcZYnSwi32AkVZ+
oxPcZlkoLKlBQLaq42zSlHRYMOjLaKeRVbJtco/SELZ5CJtA+wC/jX60r1BA5uSQ2h5FTPFYpZ1N
6K05k1h7tyTH89KyhsCkW9k28tTQOYt/Kwo3zrm4IwKD2ANXOcxPChDQtoFGf1CNEbRs6FOjRxjg
Bc7WxLVO7DH+jci6CxXZbJr3ApIrmbhAvZjqqcFoVe/0VmdstSpCY4DlGMtC/GBbCljdwahAJ4x6
/lotxf2oIhy2HjU5RPL91xH75hOU+02qELDs13pBLyg/R32CvrM8ZAu0TN2VmD0FjkOy1m+Dsp52
LRmu4Ze3412kre06rL0F33qHa1QRUxl6AWqLODzToui8fgizJsiTK1q8SYIgrKUiPIoRuFb2XZ7M
s3d7HJP1vhVeYCE4LnaBbiCElk7nXstmDMUwPMYwKS65uMIu3aiBSnQl7j7bh1nwf2RfSUNMlPaH
+Z1gF/SYW4HpHJpuCOj+rcNGurltSioT0RAvpWOdcdBeC3vwc0z4ow1/FiogA1EjCM2IT2U5A+8l
tCNG7mjTYPJ4SQzktuqPypC5rMtp3xMxI63nB24BUxoUB9JBwM8twGWIAxCSk7YiIrRWKgGlHzuU
nsDKyghnxYnLInFMPpBg5gqfbrsNk+2fppi1Uv+b/2MacRc5lDwwOtJ02NQ5MdbMj194thv8ggEg
UuL+OOOxPtwEauWa8JNX1TGnP+pZaUR1zU8IiaLqhqmLbX1UPU8N6251NzrelS0RMzO6fohdqWnt
us2m70aU/RmlfPkR592ABuTxUs60z1cDx9TDGkRDkbDyTTCTMmwJbYyzrySTPV8OpFXCfGYdltg+
cZByg48+RWiqDkczsAU116TbW0iakJWM0IWcXEK+BHWxDHWwar3MBGKxtfOFaudV4DBO8iHcV1lF
LRtNH4YbcZwv35Vq0OaUaY9oXzZtjaGt5yjltblwhPhOpTUwzj30XLujqU2nxC4IKq0AFqdtngDz
gBZnlD/PGRAgbct9FtCkPpIbzZ7PNlfm/oDmnEfwIATYOWyuB/tUSKMnl1d7Obisv5KP+mu98mO6
nKGnaBCxRfgxPwdNpQgvzI5r+Kq9ho+C1DNDI8GMFfJkzrm4WxI+N9wt3Ux5mJGzrmwD01hBFa9h
5cwj1d2k3Ce22bblGh1Tj23qYnAt5uf3qU4BiF3AsEb47IVQwFCwHy6WntlRCEYutae3mTEY/NQg
bXA2Di2o8Z/43Yc+jPj/+XoFhgVjelWhVsVetUbSkUwTvBSU5Pw3leQDWDP7SCnbm92vJDRNtnj9
t/mOivwluGXbm6J7qtEjrCIe7rv2ZVyBfOtThNASkwXRz6FPZYl5eBtRscWc95M/8H741D9lSZdD
bCOuBpZeKl2GRQBiGpp0+OsDS8q5KvKMb0csgAN4oWASjhWk4FJcNHX4MU4RZVdUBSxDvxHe9U3f
RQRog/ZjPWPubpIAk0FUwfjm3BTwsE1TA3dWRn1Jj5jfILKTB633MCV8wpi31zJIEr60hhWXvmmm
k36RW9QnLmsQcHioK854dTZ3GOXKtC9IDBJzIIoqfOFNZuSda7G0f6U7efJb1eb0JX10RAGC68u+
+LCVcdk9Cs+zB917nLjwIAa7ZjyvLpHlb1PIMQYEMHT66NqBWMwtavsERIqV/Sg+PqZgHT8sWkUR
fI3dDjxTx5GcicEuty/gH4S56vVWDPF5AGR2qWF5rCZJ/xpJZirj2Nd4By+pS5pK6e+Xfp3w6cQk
I81/F/MHYJaIjUGRLX4h6I2ws7kOdrT5nBjWD8vWtFbRTfZpiyKAVxDA07yywOSJ28tZwi7iLFIy
aXpHv6vBdkQk4P09HrafE/QkSYjYgCRF2niiT88I9qVo3mWbdokFdEipxxmrO4jUjrWmEjaZYL4v
TlLDAwdakjvSTwwDBhvMwHCUsWkVnQAxpi4ZOxL/OmM1NTVwzEvnzIudsne+VZ6QEW6SOaTQQ8K6
g1ELzw6Ygy5kpEXIs/BT5nQSgypVMGV73ngn9x12K2vRIXYiVmoSDvrQqBfW7euij9x1DSw0cY/3
J7c6iSIqVjmnWZejL0EMd7Z3/e7KPFBJq1rbd7PZ4D0Rjko2HHglPMTNHx/Ehai9DBulTT6rtMXY
jYWc5Rv9nnwBnE8pc37m+0tEn2VxEJJ1/Ms3A6xQn9htGsIC9y11tIqhZdFY1xs1cqbSD6/v6YsK
WhC68U8nGWBNuaMNqP3x51mDKTKPqA6wwQqPUuvxJ8fdIj9AuWpHPL6LzpCY38WiUTfZoDdJ29QR
u07WOMwUPNQeGMdXRIjLPFgHTF4x8YDkMmDBbNncJdiDGXJDgtxon8vp0DY40j8mTftwoMqbSrKg
ZbcJTSt1YtpuH47Dds2SG8gwpT2zhUA7dHgWPjeYb/LWQXbrQ1rRLs6j3JcB5569Hil59G1GyMDP
Wu7CSESqUgVZeW3dExl73x6yz79NcqSUI5Sy6mxetbwjA1v8bbT7LjvSY0VYjGeTJVCajTKsCNU9
F8CEJzjOCWMvpr2027SppQFkasDa5/XdBGKDtZkLkCTjPGv1O4/ljKnkqjrl0UDttrNCGJqX0fkR
3Q1VJvnlWQU5xlT+4B/8KiorSeOI01lUgqiOMXvNO1r01Se40NXx2oqEWEiZOSN/GPQqvEe4LCXk
tSyORYbdHFlSWQQvvCWH+ubyBb27fCfQIgr1s0af+iqQ3hpddoRmOYUPv3VraUGE6c24az2ggN6L
0MfO/xilHSrqOPosE4wHS966ciZQbMhYmO/LJUlwEh2QRwnCsLKsIySgr101deASV3p21wHKHbhe
BuQANxIJ4LpLICrJPaiUno0r4H8x26YlRCqtTPFXvXjVTX+kVi4J1w2ZdVhqf5/1eP/Rr6RXFF2d
UIcTEAA4SQtcMGP+6w1sKVzAbMz3SkH4OSHWlFGPvloV9wvl9bLi+P1y6U4JN7VgVGlVat2+6tHl
Qrl79Im/H/oQqWYBCWLFnT0lu+diee9/klFngY3tpySC6shRNcN64DJmWKt7WKD8oOzNQR4P7JVj
MCo6cK3ZEWVNqOv2lRsEIhfuYzOWnZ6K49RNwP2EqxWcALm9tgDzyxy0LBIftPQfYTQrdbobMr7/
ooWniCqfRp1yGKErpqrFEHqPLmQzT/CbN95M+qwCbt5cRQz6FWbvZPJwNHFgDhaq94JlbjzCAohB
PyRqeK8kjcLOzpNC0Gr0wMtVEUjYvd4AYyp9K6LJjhUcLa8p0i0hSUsxcWJfu4Gf/eeVnyxPkoYU
lOv8JsfBNr6tNhaTg2X4uuOEkTT0Eu/xq9G8kMnsYm1DxN/ZgFEYMXuv/SLdWXzNoJ0/FS03/lzF
yx+JyKVSxXHGgNfyaCnY5F0gsjMJwok8pJZfjVItQKHnk2SBjTr26cIkVmQNck7ujYvmjkHMH8OF
mGApW4gV55Jj08rZiDjzr3goGxNbbQl0sUSjvbrKY5cL1g9CmtvExSPwaKu8j/mO1qzdY/ZW8NFb
Lau5TN7gDWlAJegXiel5tUBI1mrRI9YN75qLYI7urT87K44Q0CUBWfvSUUHMO574b2LWRFYHHC9Z
R1MHPXph3CEbbEnr0MkjvvlW5h2v19Ue/98EGkQuXJ9lRYhx2FGxSmowK8jBd7KN1fBdrdMsxHVS
QdVmbrKg1YnEPwJQ/D+emoccPdpNb7vS1ZvsjgkIirmBJx5RBCQGrQJqhWV4fPbranNCn7d/MFDd
CUDK+CkUXvEtPD+bSoUBg1NTYoSvQgOxsNJ6lkP4xyP5dpvlgOx129C/7Lc21CxOpQjVxNrZNelO
FuWd7FwN2WbscUN4neq/OlN2SukKVTfPZNx/Gz8AsflgV5vtNKZpZj/ktRqnffL28raPLPKlTi/E
2VIBF20WLHndOj+95k/LsVObfNYuNTAeMyemjV8cHKeB8HsTRtZbZKP7/psRs6adcjnXDr81r+gL
r4cbY6cZPEVeXSHc053rlKxihhKcqkFbL07zXeixfRrGIMU55Ae82x1Qbn3R2mhoRnH/7fDevPTG
GViMu+0gwWUTJtZxT3SCGpwX3duVE/SSjKHktwY4Qji0j2t9hphrYOy/Rr2E62CwlzrNdg/pjqrx
zDVNoEtGirF5OK5B6TOUXyS+0YFJnSVnj2aa5i8U/bjDq3+IrF+Bi74y/hR2N4fxM7FN7sOrNRb/
XPg8z20tLbCgz1hnYTpCbNqNBnu3BqNEZOQ7fmnz0mrvZpPiG5vsxfSL5p6zFKpAEEYWgueBiBs5
mMAoTwsJTnte3hZ9cW3uPwrS4EDKpKGiswESKolQ3BGQfybxUdMP3xy0HpMVth26RDVlgKzgja7A
qlLrm4SpJTGFvygb2r3icExdUoUO8haTW7zd4W9VePpcj5Cjn4OgXed5sZeQfFEyzRtvVM8V4gbh
w8UBJtDDp1zyIJljW0KQhTMr6EPKIsZ7hgAcJfoA8ZzdCnvQ8aY9PhxDUHEIz5m2q70E5XMsvGJq
RkPLj1Rk27VC9IrjfWavtZ4QTjeVVwX/5XH8p4BI+O/zD1NNYWcAmUQAKiG0fztXnlqkuo2Srx7S
oYdoZ8Vmm0G8JPmHfIpAWqJZjW3lixV1citEzxxsKs4Ifhuj3uKLTK2b08tMY2umuvbmYO91lwKt
Fji0wNG4Mn+N7BksnhpVFWyD5SquXaVBJtH40NPl4gy+zOS3z9f+uIVC/GZDFStBgE1FwAQnWXTK
sRhdSJKV6kJjGYIsLC6on/V2+WzxwMzP2jDd9g9J8pEmF9MIjLLSfu8UEP7jqsqI7/hXAuwdqh4w
VahqCaU/EzYi/smY0FTl3wvQS6V59rKhNJrRWv0Gdm7GP2VJQi1zgQ1EHM0krEL0g/o5ubsc1IR0
xuvfpiS9b7RDFkqXoQmbLUE1grP+yS9A9wN0BXP1iAp71kJBzVrFPJ8icOmq5o6V28QLOU1+rl7u
SIffALLoEO6Fug5cuO0LcB/WY6wo72UidXMW88PLchCeZsutotWovvIQmi/nsuJIBfHVkAzEyzeW
gTNMSZcq8fCwjR7n47iCEeNG+tRPdFUmsWXYMKwMreEByK4kUVBRHNvO1u/uuLT01DuP0jhwFbWb
qNff+QqRZuH5wOv/2x6xctBb1Yr93+LEkwJB0+/5JznjQZPR1nblWWe2MB5TaNzR2If3ajRVPwrN
FBEgtCU8zlozjF+sR0vot3NMwnI89jIl9zc7zHwoNf8pURCWnYXg7htc2a+6A39/uymBpKBq8OBa
4eBGkCt/UtXRVpVfWDpSbF6QFOEOpBqOwD3R5lBaWx+UfkpWRSG7CqX0yRD4crRBmBWtibpV6tT2
rFPxkdoCxnynktvWqYV0LKM1cB4h/XSkIZxWFdWPbj61BG/lhvFg4rTebS1losU8WV8loTEnWA4b
BnRry9VyDkaEI0NCblbgIReKMBRQEUJBqPyCNYim3DTi4LYfsDxem8JVxXRSuy0qy1FsGWL/sqSm
UAeOsgMVipGGEA97oz5uPn67vfy93a0v3MsdN+AfCV/G3H0Pk2eApqzecZWbdpGcyyOueK1FN+8n
Us3z6kP4pbSAr15W9GE6EWBrxv5ApICUJHLAj0ryWnY6rqB35yD5ALJI+1UJ7B9sZ61RDEGcKiSg
3fw42b7ACi0Am8x2hxIlYT3/nt9lnK0TqbAzRsicRjvMK2Kfk3s5+tUeCS4IdMQWqQlYuilifKx1
nFQTK2OfzZQ2+lPdqPu2D+tt963X8+wRvNf9KFfs2oyQUrIU8jHG/5QvIq1mKSIFE2Vb6hDQtJwd
efIktbahhhCY6WaGA8u2DFx0J9hZcyMS8EbHq3yuYfMvNwFQIgoLvWUSiG/wJKWW1GKHmHrbSXQz
9fGR/ZSbLr0A/LZImgjMdhzkI/vxsMjSkvbGHsztKnCeTLjIypOaPx40bot4sq+5rPOi2GYDWmfJ
FXvs0/REVBDDIhFdLtDSS5QRRtMOnSAWMeZ/QmQz+91TjIlS5zDkXxVZh7tCj4qk76ptLA/03aqJ
QIhL2b8RqhtNRTEgs9JW/Fs/YnGOANPgR4kkPPAE79R5yobi/5Blof5eilDQGiIYRH3d6LeKjPwn
83G32Z4OCA9gDFOOqKHFB3Y2DHk8GHK89YGtf1TQCN3epnTph4qCM6JPQUjyEjRNpTI1CgNO/HOR
Lj/UnsSZV0Uzati2jn3ItJ3Lsm4/b+6in3ENDSTc4ov0LiOUAmbmZUUl2KsS2cBa8e6LXPXFt4Ds
O++07e7ZPi8ivL06i189D6b9ksGTnUXxesww7XeNhRm47tmXPMAzjeNCEPFmi/CgRGPrJHGJrfy8
ngKtG4alNN/h/L9AWLxkmL+YmKKwyZ1ykPEkyjcCBFRcDLgzCbYEWMdDPKOP0ddNEmzlggTUC64A
oLIcIbuhY8yF0ylJ4VFGL9OftFcc6GM/EojsR24UzVQGFFQ8m8UOGRPGhdi6wIhtDtyQSeAhrapz
cLeDHTpIKnzbIXAu7vbFznqhshTpiMFEa+ADHuiJssWtPk4ipn7NPrXy/+WA71GVGxjNeBmNPKfu
IO4t93FDgTLcZILPR4Ws89V9uLaa6OZyg1/lffe0Q/bsVOZ7+m1uM4+SsXXk2vI77D4wNb+ACCta
4DYZXVFqwMQo0cPWNI8KSxgYw7LuBxqMdnAaJj1y7U/AJ6KyYt6SnRmiYNbAKi/T/k5ERevPpsHF
5xoGV0DCKubOpXP7c05FL+RlY6Aa5GdK0FlxbC5Yrg0GnMKc4554WULNqj9/9ZEzxJPhNB+G3NZ3
Oy3lupgf+khX8Nc4z1lY8idmNebjLiN/Lz39U2uQ/8En33Bj0cM4BKJKDB2KxtT+A/Ue7PP0Zgh4
G+JhxeDrUlmBA2xpBE7ig9u5+XQymXpRY53k7dE96OgFtLPhazNxXVTIXXom+WwWCsNqIosUwWn0
3ptjdnGHaAAd1tB1zsSAz1IQTn09IIWj0DaJmF/ITxclil8D4qNoTZLXck9B8T5CmrX133GiTl5N
UpUtWxWgp9a3kHTQHoqlJF+nSU5cw8M4I8OoElJcl1eCGUYM75rrFRv98GOZJbI1rQr/PoBMqhRE
a905MrRBSE3zK/Mdq36BNPMeW/cXiP/PzkjCml0QRf4huqjo4P4lKQ1GCjcxa4/zIznk4ej/cKKV
c70nN9T8NkSHXwbffFBFUA8T6ONaAJ8n0G/1lx2QxXUJO+NINr3ABuZomL0J2dWHjNg/OpK1o/Qg
kjkD8tDyXEEBWFhBugxQ7PpKOd5OEy6aVtuPC2MJsxWJsBg1xP6B1BNRrWNx5vK6zutBl4kzwrs4
5GmP+aqUHQgcbY9vGYtSOWmrVg93yo76dZCQRaScgwpvfPzY/X8x7wM9T2leghy671p83pNrjDyH
gQS6FioCqDB2GJe50dnD8IBkHUwihpZLuwbMXyEJdh5fRTKWJsbiUEJt0QvQj6EF2nujfRtrXUvF
ZNmTbm6jsFhzEo82xD2zqLIyS1wcu2f1iT2anImwWbt7b2sllcUZ8ou9zXwH++4L7VPFSrs0KPet
8e7mW5i85/kTQP9nylaO3LTksf7lFO9rZ4m5dKoTKh/PRhEzvFBfVtw8cuo99OCulvyiEsBYOCmW
ylZ5IN7JU62QTUIAN2Z9XdgNzhFIuzqPRcTh5dl7jFJZ8+RXd2nr7ORuytq7Eqza5lMUchZ4t5PT
gJJzhyFriLyg7q+vMhx+gf+5a2gmjwdAPUNn/g0Um9rlhB9lkt7KYv8208KUhh/I27KAc+6XmdfL
7/bubDDCF5gpYz/ke3G639eY9WVuYbIfE3k0+Hljic0fT1mcUdS3YhVuRG/6YJhVNOQOI+xosunN
3vLjYB4CQSzwi+nL6NpU6sa+y2getWgwuto9K1fYGUwPHRd91B7reo6my/XwM536deLmCwEsI5AX
Rka0/6g0rUzw+sVhVadDQKcSQRFvh5cgv3yCU7zEcbWdj8odXPW1y10ALT+LqYTYnpY9mS7fAfXg
0kkiPWc+qTGhGdBuGyQnZ+SYN6qB13+oHpP4BDGzqdTfsBDKadBlkU9WlG6TaZrndensaDLu+dZl
sWF8+FQ2pWIq9MnJHhppFeHsvKVN+8orrgxpg24UEeiHuvYqG37hhF1zqwh5E2rDFnSa/DVyx14d
zinZs9B1SYQ4MQYtiwiuhcb8bsqtU8X63vELwsDcEwpQ5mzyESkeWlecgsiIaaEfFdOz0DQY+Csw
AxiBLdeLhh3rwUmC8zSDyWN7/U0CSzUumdOo8uIoan7KXO/z2uO7AqFWfexyxHaqzgV7HQCMYdbx
XgwIg6GfgPk2Eqgw7UiQHhMi8qSKqhrpvLTGcNS540hKeiKFCLOiyG/4Xm1Rj+c2j8AnwtMdIp2D
k2AwNd/7UKvejUs6tJb0ZzpVx3xFhefCPHUICOIQhbz9GL7Wi74vTivub8yzVyeZ8o7hzvjn2sD+
JRDkStah5ASHviK5UiKSd5Ux4QdrFIhz9s8LYQr1nTvnoxbOah+o5+KAK8r1hhChSoO+bne+ut4j
Vi9FuSmLGiO2xkMaomMY1QTRigvxkCVOSsWJMNBbWsTERIvfmgaml/xcsU9grj4Xr/hGqvX5gHzb
3DQhteMMaJJ8M6E+VzXAdHcNIa0Zakfy8GbAHMra4qwL5Iij8HnkirgXZk3ohnoFBDGzu9XyXDIE
5tS4+56PP5axFmvCyvDlDVm7rrNHhOXf2UgxwbuMD4DmHE8WGBxktz+Ajkqf4QZX9nGLlKdGoI6J
vrK1tDrvdYipfGNT444ww7M2qAeNJMx/PZsuc8w+zHkJ1IOR6xe2R8weiW6wMRZXqYsWNsbObiZ4
O0vTnFRiF9zb9nCz3njgPfAruyM7eyeQyF4R2Y0beCC3JJAkF0iuL6n8NEKHd3yIaxiipIsnS3SZ
e8trFYouWq0SJXOsL+SnXXZgzMDss31EbLmhg3Yrqe1Dbi1sc6Pccj9JBahDt8LTKOiOsolRVMEi
DFTzoO45in1O6Djxl/h4nIq7lrZ/4B0buK1+N5ldvvV28hau8W6KZYcNKXURy1NBI9mqTDhXaEJG
rhvNkKqWyBBqBv0/R09Yojk8/954JtcwnWcgiOT14ttbMUL8AN1aVeOpyFrID/H+1aJqHZoUz5dS
yKoZLsy0MCGvgd15sCveRwWKk3Q7Y0Sz3X+iDu8VPvWpr0j0uFhjzic3XZmoKktDDIgoj/w9uq2A
seP4uBZGeOf/riKGeyy2MzBzmg9Q+ekWhwx11xkSMKGxr5TMw621l6bd1OMUOHehYp7Wqaiz2IUc
8iiGciCPXzLRF1hyAeWiJx4hpY7+eqSslSEurHByQR7dubr/5QetWhdzAlo5QQCP5TQJnYJPSfJK
4PXInEjdE19foqnrdFitUH8HJI8SVZzSVpQ1X0JS4Ci3n/DjRd6DS8uPTY2CBEitQLUkhFPyF319
/JsBuEpd8gypifYA8NTT8hILmVxZHD519PdgJGidi1xoYbaolCcE5H0qmMkOLgHOqC3TTqUFWil8
fFdvXaMuAAwPmKxpVIXQhAodABvkwXz840dzKmhQJfEQ1sUWHD+QwVMyHvs6zMFJJhyjJetjQz3l
i57C6FEIaWHZpa7m3lOyrqT9yFOEkN2ICK8Zgj1fgBPW1ZojKPhxNJuomkJpE+o7OM1pGe2XUY02
hHtChPO5ABIkxRcmOF6CnWynyh0ITa9Fe7VmS+xZ9sqfIjViYwCeLOSwPBRpqLAXeIJaFPLF+Sy1
V3us4z7gCmP5MC1eZOs0aDix7qL0t10O0OqgfqcDT/ZO+AYYsqvSzHbMOCYmasXo1naWv1DQ1mC/
KZWH1mRNxXKdEe/O6uiChRFmF9DYDDeAhUqVt1oXNtOaGKC8Nr8umaqPAWCgHsZe3t7r+0sBZHJg
2jaSPAOwcNq3/cfUee23+VwTEJ/4XIxqyvgL1b0h1aI/lSU1yv0RzR7mwn4thv+ZP+J+/wt0gzzU
dyLFhQUpxbFu2TqUKpsZA6DbLscBPW8pBi7T0lGgibK88Ls4NVHCu3790Lu7jXt+Jx3WQmV41QZQ
i+O42NVKPtDxGRaa6du7l0fblR3OYitna7bOfkGaEs7K932DEm8HgKVjgKAYMtLUfKOiICXv8JdA
ny+XvJrSE4kvROdMao/T0FEmNDnugNXgQGLTSatWKovoHg4e3N11ujfCLdjv30oOBSWdtfm+YHLy
QYydoonMtTDCJ23TMotu06rUjrc+dwV/SZFXflPIwT8JWaSkxquajbD5TU9XR6TjUwtMRZh5aO1X
i011Dy0T0sbcgCnI6exWc93znsLLFL8K6pIs/5cizdhTyZNA4Y5UQDXUE37mGTc8LHae8E6V8Ukd
GLEUN7LGEpbHB7W756jgMFE9shaSIdusZ15yLnMIXQCAzcBWrSzSXFLTgLgzx77csZMCR4KCJseb
BvNKeC8N+zhu3+8aisnNy112UHCh26gJPqXEs4oRxDoxNxKOCdcqIAuKt1mEnPB3gbPbvG8Frgxv
0vtloTdODuO7m+vl2pSR9XmzcvQZT2bWAZML+2jgNKrJ599QHG8op9uJ1YJDf0edVquRTOkQ3tm5
3w8nY8EF7rDME/3wT8H+xvde9SEboyS5MZXkOrTcxujfmU/X4i4pdCnmF5WCDneRu9z+vCY5OFtZ
vRaMlGWqAXU9ZiqfALjXHCk40jZCKSJXJErfsLvpR85ATiq8HV+wnb5iblsbGF+R8RWqeT7XV78v
hYIrFJ3bbGjsPHq+sJwlHli0hYjqmyXFQa6HHiWNZUMfMo5b/x29o3JbTggC6KrzeK2+knXEIzP7
E7PwyakLU+In7Ylby9D76EcE2tr0EDhXIuMIdMmFT35KprShxZQVOQe4+C4TLiXTRXEIroAIDULW
lCDXuGw+2uFSrIXZ40PWRvEn1O2TZ4rFnm+IWpEYFjOuvKMsFMnRVXVD5JYpl1/N71IikOMuISOQ
KJXAcA11LTadF/jOLm0YvnMrAHdUfhzwmmGWg0aQ1EtkxvZNvX607ebEZSMNfp0qE1XM4xjWgtM2
lDEyha2Dw3zjDUjwD5rnGmf8Xk3Z1S95flT6yB5+D+heF52h4PyW2RB492UJVPjAQyLCO7xtIHtB
sepPf3/8tPws611vXVKJtRks3+RTm/UlAlH/K4TZ+gKVSeN2os8sR1AtHVkKbo4/jMw3Wmfz4wFw
Z3Y29v5Ey5wTcLBlU3uQRd2Cq+Cx5gRNXxvoio0doaM86LEghX/KcDIQAWDvN+NMfPcwAHK0Q1hO
jfPzzdsfkWfFxN/+ytYiyEUonEcQUkKokOBiUyVbBSKjTWUuIH0y/hrvCGuSsQ+EAnw0F8Up5gCa
VvkzWX2SHnq8H34P6jrifLXnMu4TTNVSsUGn8MSIZOH2iV5Yv+hxv/56Dt3LuRu8Fza+aLIrZfm/
31TSinu6vXl6K/g6GUwYRL63l9+cG9h6NoluGJHJXqrYGmL+OuYdaoLbQQjNgy2DvFhFRH4+x2m/
RdWKpbS6+ME1tnyUOxur8Jvt2EvNoXFmU75smpH9yfW4mNoH2SV6+VMCBe/TAJwQa+B86axs6a8V
ckOiJEJdocNEll4NbluWhKBqy9iUC+rrfbtiAtz6ETYXjljn8VY56SHpZYgKOp+85oRizvLQmIyS
qJ/tZqQUCjlp27CCFL3AKxRzr1rbrdAbJrnILvPm9SdgOiQWm415WCm2Di2D4+EJc1mgmbDcZcU2
uTl4enf4XZ1j8gh/fnvr1Ss58PpdNLkp6W+uWO5DbRlnXa+H1IG4EUBIj9OorGbeQlWf6gtha9O+
k+wnrAnD/2hLhQNIiRZANWbp4j7JeAF05Np2J1kjB7GrhEPH338A3d4a9TGgzxORa03aP0Viouha
z3hjxgcLPgZCZqstSu3XaZkgDOKfm58wUH+F1L1GjGOuSuldF3lbCoX9d4gpk3YInS9G2zg7sIW1
P64WB0FAV5KELc7g61aw7S4DZ6u9Z8OjXgQDj6mxTr8gfxoVMBBtUovdgNHIweXOrunp0uxMdOZl
Hn+imrB7Uy6jl7kzaxiwol8jT4E4+CApAoKuFbrSkCsNqpP2lKBDyrSqorRquoLxoOhhgSVd/Ulc
rXOHESoaB37IEB7+Qmh9F8KIHqtdYxvJGLveyC4sU9ynfSF/VG98D9LRgLS3NdM4J+W33ke/GWRl
49RiYjBRyVuBdrTlwOKsGzH/6lPsSSzrGKuIh3EXmQtsmrfNulkC+Avy6CDWOLynvPWKP1OIT4Xh
OlnL5iEDKmSozwtcdQrsX90EL7jrEE+6gQ0xWLHhBJlWtCoimtssrd3csaNCiGqug83YJMEHeWwM
JZS2H00HMB6XC38gVL40LhfDgLbwHF6ytsw7955ORY06yEm//RyOqHjS0NzRXAWa2pP4YMPS9VNw
agPU64P1ao8P3J4gmoLM4GctYLzWOfEetNLMmMv8Q58qGgdcJ+V0bbXJOD6Y6kuUdaS2hVZ6+60g
c9RQalsJqcTPXoInHFEce9i6mFIe1AIQubvaNfjUfzWY+nrZF7sYhalbivZehNTRyF1SyZBdmbHL
m5VomngpCVwHEOe7lbAFBZXTufbH5+HGkLG/sDBTLqrO+a5t6lVCZ1vDeu+LgdCaarh0DoZmgUwO
TIcFXqGhLBei+B6/4YA/LKGBUcdHFwcWbSzJz2eeoc6UQmM45UwGPoIkAPnbR6PaGTgXafF6qBqf
jFyZ7ZpWVeMme5IVIOPFgqikyE452fQMnauYiQju5WmVC6BjdX+O0NWwfjWP6x5Ie6vQBWG6i1v1
YYDmmMFbHsbDmvbow5vmC2QVwlCVXdwpqNAxBj1GOERVeIzOASxEaM/bpSnXmRtl86V3OA5ateNI
72htk4v4WikXrsAvHR0UhR1jS1RsftbFq4cclHdnmU4tAkli1oAUiva3cP5iidClautfrBXMHHyN
Ppv4QVDwng2prRT94dZhnfKRUI8PIuLKQCrZ5lN+24m+UCmJf0eH/deEbbtlUcD5wf8sjgGmuses
7qTitYcQpeafty0y7WVRlRfntrki0agDZhmCJTQwjRxMQ6jdMQPSx6DEmTZtZHveyHtRCxyysu8m
oB7M1znC9cfaB4ycJzEQDgOdHgHdqn2qif/7vYb3g5L14ZLotRD3WGOnwMgK/vs49v8Cc3qK5bjg
3/B3+uyO0YW2byIx/k7XVZ6N59E6hw67DiNiosJsCRpaRsSNpRsjQX+F00NHDQqkX13kbURDy6v5
N5dHFLIbYMW7m9cyc/HGTxfh1oEsD++gHZVlpr16SrTM+i/IywkvceDwwoi4DPQe/58ZAY6xnrTf
tn9xeSu2YZeYzO613kjpRFZs+IPe2Ni0q9VleaJ3p06NTO9apv+/RU64547+jQ6JWWJpz7VgrkbO
3AbLfvjeMvzYdTDb327FiNr3pR9dLsSKRE/8vf8bk+k256OXqd2OKgcRT7p47ULkrcFRD9ub1sgR
kkv2e8aNBziqtMFwAubkHXwMlh6ToVWdMLI5Nnhes3wJGgyFXUv3jZnRL9QJ5QnQzzJHx+GKMQRH
46oIYfvUHEDPVtDPxQvLkOzG5nkSmBUviUppQ/Yk4H6uWW45a7uYuLvu3Wwf3yz4X42iOORUrIOj
AgTtLA/G+aa6VCELr41MeFTQWQL0fbuYDjMmG3cfI3Lv/AGM35+H1tj1OIXAfRfj/K2PYov4pARD
2VK2pzFDZQRo3Q5ZA72xofWI5kJIrjf83Hq87ap9eDaWnmUTErwlzUAOtDntU8zmcb9mv7A9BP9Z
pmM9yxY240mfBftmDKTvdK97uVdF3rVMjvBMhEcnq30fc7MG1DE9MpBlHeFVjMk45cQstgIqY/qF
Z4TezeiBbW0+2YpbkNBNPXynsUgrhwMINYMdVlsO6lOli8Y3nPHWKZY0zQStErpcM5Qot+fZrCVH
iWdjGNm0q30/xX01TuRkR8mO5j/bTux44p3U9MONlLLwG7ZjPxH7g6HOaEkwOKIuYQOkluLJczlh
piXPyQ4t+smRHUM0FybLJYbpEScQrww0SXf/hadT3PYDX3mo1VW9ii5CnOqiSV8hO7WmUsaGOcbq
p1CH7gfVOz1bYs0+k6qyf6cks1KkYpqaXBMQVwvNdatmCUXxtgQLqBhhnAQzJide+Q5lpE79+WyB
pqp6ETAZRnB2VFpqqe3T9tngkJYOB4tMVYcwZYDlHPbR2uIx3kE6m0NP9jKRIxOzfiqPuXvckTtv
SERcYvyeOs/6B3ha42ZNzx0/+h8XGuUBooH63vrBNrQrNze1dFNzINGwCyqluslt+YC66PZ+bqgG
yvUzBDBkmd0NawtHZFjI/mZmr+FLicA7gZAQ8oKlkWO+Res3LmO3SMeB/aBT8Q1czpSp80fQDvDN
Lt8ompITaen+tfu87lBXOH3Ow3UPt9a4jEAa/ewY9VbwPxtKXcSeV5grn6CfzxXNOUXFDZQDad6i
bT5GgRyYW/R0/tmb1NQL81HSnr2xjWRNvfZ2oaDWvcyCqz2HS5moRZaVfMOMxTlQn0iSfbzwFm39
pQv98Fdh43jGy1rDmDsgspZ5DpAc21kl18TK8R4+Gpk0TKNRHDyj7pIKNAEG7cYbmUghLCCBmUH9
HXFo8xTAjVqJrw0oBEcx8cI4UuUuF0o65dUgGaPDtyHYY5eCq9u28M9IHQdppUe5wHsMzwgkEinj
sLTeN8/F3FxfOGnPEwtZe3n9ROPI3nTHqeMTsWDMdMTQdfmXHl/EfIDEYJ+9wg8/uw49vrR1Y8oN
nr4m3ziTgmGDYU+4rJ5PvocI33foP5uJPEd7ZxV6hUUmYD9RONfylmRUo3joteWiqO4laCavhoWH
UizabQgqTNr38SNAT+2USXgFzZmadgqX7gbOKRa6xPjDAw+3n7qnQLN1NCGhjgIt3U3o8nUuy85s
ddULcUboOWiNvEgZN8H53Ojzxs1eoCoRnZ5xPcrDMfuyNvNfoFtKmDvUOKmQsYlSUZ+FkuQYSGiB
v3Brfb+keAAwsvwoEMQubvdnJUWr/7ZUR1rZ3JyYGRyZFlt31IG9j+ySfxAkl3h4CohPCdjUwac4
ESt0SJsxCNwWYhZsjklHZlHoK8vWsdU5DAhs8udvg25bML5RmVDwz5SG+W9KVtFE/gVyjK61z6Lw
UodU8mKjXkRGbYYN8SYtHSQ+RuFkh2o74/ZpE8mcbhj+22Hw9kwwbcvE7nml/fHXOOGMEfCTpZ30
psLNRdRvClLfT5EuMpx2u7gvD71ayxo02dr+IbbeNwzd7zSgAfAmmSHlQ3yZsOENlRlyBBzkGNwR
uXB0WvGFS7EIjCdn2xu/KH1IBAYoxbW7Sh/91iMsLenUCCO0dycc0r9cgyfWb0S2jPFLaBE3H13c
keMlBECuNF2r38uOYRcEd8KKhQguGdmWpM/8VbzZAsDyQ6T8CRuUrxhditHysbTGOx571bXKGR45
UyTHbFyGaxbpFDkA7Rq2YxDZXMljB+VMJHF5MGL/Y/M+srQVnSQragOLp/EzzKtiKbCixay8EIwJ
tWsTr3QdI+V2cohSSkwr2Uhs64PQGu0VtDGwOOJcw93wnduTyWwjbu4f/aDNExA+tin/phyDVRWN
jO6dKdO1xi43feRK/vSsVm0LDJbDD1bIhU2j3wxS79oq5ARW8NAC1cmw2dz9GwKmwUju8Vw4qL4A
eAul+VyL4INu5UzoeoeCqug1Yq7J1nexEpYCpH94roXfRmA9ACg43JeCkhr0smHRAWdZwLGq5IzM
Xmt4bX7M0G6PpUo4sOOs6o1nvFRkmiKBce5qquKUolKZNKYeM/UmSNrhrX0bwjVJImhpJpGxdtSu
/qDXR6EZnNiNZxtElwLEt5meidtHwRuHcoI5zXDAzllJ+Fnyr006Ug+DH6auu3ng5DG0MLiko64P
OqJ/dSJmAb42doxbdChls11mdwxDwFD0L5NPAViMdG8LqdZd9cByimbIGdHkTNBCa7sunGkj6JV2
2YkfC/CcpKMVzFFofPLJDdeSNQA/e2DhlO062gP68TMjWJxFGWB/yk8VMDuURF0z56hWLu5F1h0n
cjiF5KkzTpwitDbwhKNkUjYF3g+/snvSh2LdCd47e3i/GHjnc/6DYnXYD2TKGJE7deR9BTcMKRK2
h0hPftPMav6qCmyPhqbkWVdfB04sUzCIn/CY8t+u+G0+ks+0BZ/F9XUi1LOJ64HeXO0L9pfpp9ZO
xF8Na2GChwa9BxnTOPT7oWqf46KL/J13hvd5LGHKFNcHbwo0ccFzakeStCvncqLHKQtBqBPkfPf2
gHwPfEo7d3nr6TzHKnRE7bLmUA2fs0zLVtoaa99BTjsU0pgqAwi2hi+eBxFDmMsOjJG3XNryqKcb
k0UgdrR98a4hy0O2g3mNJ7o4osXyMHftXLnMSkwwHBNVYyXMxpKfJ3fz6Opl00pzp2LeQrl27y/X
qG8XLjg6OfgxxX/nb2UUSl5HYIX47GtuScXGX6rxn+LB3c6aT1uTI8W6WubnGrhkpD01Q/KDWE6k
2DtYUBpFVyLKdnNLf6Q/zGY7+6p2P3uybY8NmewIJJ5W8Pp8QhJigwpfMzlcezheM3k8Jp83irtC
ea3qsSyebGPnOU1rv/dTUypahYWw40MgwRLHZJv/JwaGz9MxnSyJylbBWJsZ8CmLA8/ovnvLs011
f2hmCdEv116sM9z3hq1l+FZDeuOTS10D3bEJ8auREVkKn1rOq7N6VPKxx9nZAhfz47Gs6JKyCWrV
vmkiztLKRjZcHprPjk7wmM5b1HP/+tNpZ/QbpNs11cXDKtExTFrREakuIcLZ4diGr+dZp1oAjPqK
AeIeUdHIScsvPr9ce+FPIT7Bc8ATKWHNBsaRijodM2TvL8p0FQJKF8D7gFLGFD2V0GpCJlpAA8yV
8KIxofaawRTV0MpDe8IHCzkL7KwZrJ5VNv8juZbhvfTDd+vfTHqYAssFTJqn7cNVGrNuxJ9W8ku6
LzUfZOOQdYw5eUpMTTbhNFZFGGL7XGzXn6yxzGSpWbAzb4mIKF0JvOgg04j6aEeHmqV4X83CPXNq
dVEg01qQcWhpYXhvvv5SKITWupf5J9OyRJOxPO1Hr3GIbtZxRdwdUjT0MPU26keXLw/V4dVCJHF2
0cP9TjyGMBDMNUztMgJHZPDqhBbj1u9KPl2d4gCkUBZQuFL8W6rAkfpOfzHEQE1ot7cCDkKrg7sU
ESkDMkNSYwnkRZ9KypW9eo9iv4y16VJqBv5x2Vr6Lm/ETUe0LP4Ez6rubNStzD9kOCNPJS9m0PWV
1j7jLuwESffsY9BO1pfgvLY13yI1J1/JOjsFZwkbvUir+RmMOvR+U1g6lxmV+TxZDEC+QNP21rxd
utEdnppJX7xfIMLmGqtU2jSSkSc73DPUYRSDDfLEHPailvNKoKlYjigCGFPAi0JbhFTR+/lCv5Ir
m7usU5U2TW68QUHUSrBe5Af7rVTRUYPHQNjZmaHYDUmeowNi8+pBIs2wUyJHl5rsw5eHMUi6floD
h2V/EL8UPtmiaz0DxgTs5Ewi/iEPsniN5bmm6rdC0r8Qp6iPdBRrI3b8seD12R+RUaQhkOtMvR71
3lQs2xBs448kU+0Ab131TAiDAQud7mXIoK593CJUiaKQiksYyKGsZiONfTshV/nUNi2MZL6EOyaW
mKZf8xukc/dCzUEfXnmkN11PyKgYQZ6xzwD7cFyK+ku011XOC9ZGO13dkiTR5mkC+jPH5OUqA5ZX
NlXv7pMAkUmAkeZW1tGYM+j1e6SNmS8eXiSRX8IWiXwc7Q79xBD9Opk6Id9j9wcVDEJSqeEuyHdJ
Px2CSWETElD45xCpRD5yFzyV/vKDCMe0zvk3MzsG0/XpfgHC3LF5gJMUa/FhspY3lNCeDwDxm4W+
uAYmWpJEyQ32VFKtIcyx7CQd2u60qUMBP6GmOSNlJtxM4XY6/Pqh5tZjC447MsAhNswl7bT+7Qf2
jrSI1zQmW3y2S3WoNrD9zEjNVuymlp2rJhC4OIELBzjJ3itkAM4ZQPD4ev24h7w7xVtZHTcQ4sFT
LCSUdHpghVVixcJaL7vAkk4zalM+io1PI+Zrui6tEYihOk8zv23HulEAok4LTlst4x1zROIpltj2
FFhpsYVCzhM0YbkZlyxCCH0L8KpTfsUKk1QVRNy2rgocRl/fGr651wYteufvmmTTn3T37gUJpeZP
xmOKwvownBPmif40J9e8oXlgrEWJftjLc7sjbwfgsYyenJwfVyAIn6JiJHDktn9n3ngnMu6j0Rir
uJnIszdILaKGqekMEpmEMSrvzEj3nyDlrz8YcY8hZZjaM1wT8Aa5W0WuPfUrL54KZ+UbDorvq7HF
Gcz3y6CdhKM/O68lp4oewxJPo2DJ7iTduE2Xo00piHkW8ZyVYw6H9F9o41LYYMDMnfd6U7133rk/
Urz1UJ/GJ4iTe9xCuAn5ydU766WS0PG15tXCSPNd4QIWH1+YxiQlQEZ2fHzR7xWlttRS0zDXrKkb
JJiY4otrQz+hu0AGuSBt2aN99tYjl1kNNzWcIaSJtoZfIQVy17zLazp8XiUfw5kJi1KuNW6GO7XD
CZYLt3tUgVLHdE2kuzTdglkWib2r94w4xTQH/dJKVP81JIzPPuCiFeIEMKW/cECqa7anNsNKdeLT
4X3MwN6IWTHHULwJPHnKOkknWGyfKvzs/VLr4XL29HebuOWtFtJXtrXOjSqHYczX43WBAZoHCqXj
GTUerbN8FVjU3kCB2xCw1LxDuSPszad6zbYfBc6rAnWRBjqFtCKS9aMsYNbwl+VH7Fm4BrHHXNxL
JGkgcZxreWCWWzhhZ2R+3hxhp0zkI0j3oeUsE24QxUqPHm5p/y+4YhwHkPUllSOv2b3NCeuPcxGX
nsxrVd0PLFRRraGX60FhYs7Hb6A6sVbI9DQaQI8Pd9FaBQsjuvNApnWc/wb5HbYG4wYhawBlMG8G
2v2uVme8/sR7sTxxlkON9qr5y0bVBEtDxqzvRBYVI7Z0i7rMs87zn7JbbyoYZkjunTjeK9ssPW4A
u67y36tNN7tmgi0/QNA2k2T2s2gkz+jmidERxSUuXrPNjWfsUdarezuwE8pTFQyPaYDzRoalb8kq
pGhA9kEQSOAFg+Us6YUwGB/H887Pb4k58QqSdEUYiPpOTHCjhOXS7nUKhJgakceCEpeaUoPxmoQJ
m3wMpZZHcn7ed/+5fgl4sP+F62JU/N0WXlXea+YdJg3YLvveLOW/96FKSXzdNTl27UwWKrZTyvtI
AFFWZafOe9YXi/VEJkLDiGVwc05yjDg9jb4dvU+5BqxfVzXk8G+nm3k1UpjEb2hJ6PP1zfnD9k/S
1V4IE4ebjMPT7dzWfy7bPIgKn1dr3ZfYvOKx+2CCYzwGG5OW6n06oQwdaqPX3pKF3G7U3dhon0Yd
VLrYX/oHMtSV0RNjzYSgSa+n9BVUrlCtKPQuZauqV1ynedbwMNF6Srbj2aG+rVQG5+8qqvhVf+ND
L1/DjAhuVTAZ0HuIHWwnbaDWv4DegVGYy6klZu5vaGORXGwrZ7iysgyHxlXrk0Efy+thibRvPl7x
Utwp9XfY3zRM2rVhHurAWbpe+js+iAXmfz542yKmV8KMEwyHn8B48Kzp//mkm2nT51yBo5KjjdhF
xIAx8XhglaNzt0/88AF4yO+kqqOPNHZjG4H6bX+QbmnfT5BruYdvY+ICnFqwwv2EGC36bqRUS9fC
fJrBJ6dwn/Hi1cSkqZ6ZgrlYk9udQdUGVbyp+TpWp09bMqS1UTwldCgCybeBkHkHqrX04iU3kWCI
8qEXBP69RWQGzqrGmB4neOvR3sTBZ0owU/Mv/0upeeS1/o3y7rzcM89+MvGsKc6oKfkYv9qTTIVG
qmS6MFLaXFX8cykqPVdODQSOcnOVoEDn0n+qLAMMVavkVCRbGIGyBW3Ky9cHK4a78pCzM6Ko7xIr
IW2KHOpZjBKASkmRKRJ5KJwzrn1yME1Q+ThWouTt/BLhAANIBDVVt+gLF4IcHvwb1LbrXYazsJRt
5lMoTI7eX1X22Ued8vH6Hyb/RCedsjrmadVGQ0AXfyWdAWdhkNaT7OqXLMatL2vCRKUFGhvKVwLP
0y+S3ylbFbtHtxTyLD/R917PkwSVGejqR5V60Z0A8IQTuJsqEEDj/qlNGtrRg4T0UsKtR6RWuC7o
wxpSh+EqqU/ZiHGmg7YzGRzFjRVO6hZQ8+Fn3Illz0UgK3WR36yEpV66HCs01LOwfyjPbpoHuoa+
abeuR+IZLwJKRk2hKSOxqAg+cWsbsaitKc12sjTx+5hK8zTHft6SfgNfSnlLm6fVaY6HvbZ9mYHW
4+SMuGCLQ66Hb99xUnirrumsyz95ymZ/RnF2PealTwbe8rb8E1C4lGXZP1k1FHs9fDLm6WafpSJU
/tWz0X1F2g6VyuwsXUsgsm8qZPOg7R1NhPKNQc4Y1752XQrwAgYOV79D3l8FD33WdXNrLRNt43Jx
IAECThr1dHsAlK0iinnWYwSwWDfK/K9Dw29vWGpGy8TTTO2YNlLKv/uJoXOrWN+CVu3FSErBAMgk
9660EzLI+1Qw4+6x/3e+RzzriNmCcg6aAEo3u9rkHAaCDHfpn2z8tluEtO84nhvLpqtdreaKdkym
3Ar8ciYq+7qWK7k4SOKoZHDKWrj3uMNp4npLA1xKJgYR/SccdOkkUzo9ome60MkWYu9rLFxF9A7+
+F3t7KS3eHFYljoWKG8aCUUxRueUKwpIf7QF0NsGBp38R7GgXkuad+S+RVGAZEHKfX6/1EoX87bN
Ei15nXATPFjo+vb9RcbudrWoJ3InrhbB14RpUNiRBWob3Mqp0e8enX4poDJSGSgTlxA3bp66Om4Z
N12qmzEVY9HB/yTMHQmeu5u6pp4sdkiDo9lvDbsJPF6I9g1hoy+JNdKwYRGgTAn9/ycP6B/Iec+c
0sics30qTFXEydIT8KSixWVSO5rfTZ8QggaYDZQAd918blAOmEl0L5s7PyxKiev3+N10KFQiahnO
ZC8d5gVFfoQ/bnQz2Sq2ySQGsDkEiBFtxzltV42XFId3VoJBrgYRalIUwBGiPcxWZ9TDIokIOvDN
U/kxcDW+SprgVGlO4NnyrdcluEhnsg3Chup9UooxStb/EQGNeaiqqSePygartWnEnmz772iScnYE
+V/XjhNnyyNtctZ7ktMg7Kb70UG8x2oJBJcDNiCZ4GrNxeS9m7sIaDAmlQd0ubjmOXybs+5Kmn9U
YY8SwpMS37B/Q+QlzvtNCvGoAejxABUF9rQ/sPFuAWz+DRPXCNe9Hy1Ccj2ef3IWQcWHHklDrjEa
7XcpVT5owDnGK2LCgkDAx2/ZsQdVYCV5Waq2codnUTzBr2/B6RaI9nA6dOuKCBo+H0oq88MJf1+x
hEGMVuu3JXHWpclYK1hD5Nkx2GmEVIXYzI3I7uoFCnmiiAl0YrWfQfuJXBT/FYCSQfSXNjZDHdEm
qicKsiAOV46nS1KSFZcn8ij5tJ+8ZOU8jEkmlvQy7EplCApCR2FQ51xw7xcA4hVnsMcVzwVnnoLD
v8aFMrKZpp56q1K89bO2nBt2c+8geMAhpkOY3n2gaxtPUlK+IhqOqoluimogGPH7iqeXQlqnP+Xa
zj8xZN+fmRwbLYFLJrfKTNPnoSM9fDBv5dQNrVbTb+7+CFKRB5K/wH5EhM0rmtPqmoM+tRHbf7Yd
uSJ8wxpduv6Zm23gyyugJQSOmezF9bS74EIWSVjSM09KY86jfykJ969+kkGyzdx2vdEQZrtY50+D
7z4jbwACgMGHdmkXMZwHhR/e1yIARKhSdMdz6akD2DaImIJKmuPS4vUNeSyZ2Yq7Ojj/yZFxKdD6
GF7FAjIvPogjNkVh2Iv+TJxUZieYP/FD5pbQiRdziin1w8YSCG0X0lHmZe2SAB8XbG6E0TA7++KF
vC7mQu52KxqLLmlPop57QA6mi8Banze/7UvwVSznl1Um2MWHhLxBUYHvbzv4pHEDVZOKzKb8v8Jj
M3784kCs7fz0NEFHJhj1HMTgnbByCf95PQ586pkzD9Z+aguSspf9Zlf/637hhmyKbIU66ufqucPK
GB2R1B560dZev+6ESJe1lWHFpwUOSrseyKkunNwTZ6P5NGuFqrHZKV6BHjsDWeQLrh13ydg6TozF
cAEKGrgyIvB6MH+JipMWkd8GIo+RY4sO1ZrO+XIlxDxs9TAIpY6YhM+FG5KTqZpxY+06U9D77si4
m0USVCGKCj2LjglbGw39ysIN5nHdMRE/49WB59emfCAoMrNdAvdT8Ez4zbNoplTpd9H/s2Q841JR
RNOzp68EsOcaeFhZuXm+n/7/4yRkiaavVFc9+dIAwmuUgh4SDQVJ0/eevvBoUgBe4TaFtaxm3ISB
A+x5yLVjyCs+vpixcghbry6+qYM/wegvrFFr7UAaOs1lNv3qzkwkBo2VUhrIR/KZYPiAQyqPwJtQ
llspse4THXno84Pj9N0QqfAZq9KRbjUT6ixNCra0bccrqx2suKwnyy/dqjLDBNCjbo80y0kWB+0d
jre5zmdoFI7tne4tvLCigPsNAIljF+ounRcY5mnvULQXdn/Xp5wK5/Oug+oVUyGmIopvQ2C2Kyrl
m8tCOfV9OHXFPRjsrD9TvYpK35SazGGYDVgAHarOHo9LFd16r28mHrrKdIeYUQ7fpWvfBv8Y9yUY
8j3FHr9N99kxyYPlg8jiBzxAHXNXfbq5V7OtnmySj7PVk3rj1c7dd8zYIq+WCAI3q1sk8CAP3xKf
e0fPagZiwlsXpKRLgMAB+TFN4h1/mOWeO1cvaBsAycAt1knaq4dqrR4GCHt4BpTjtO4Nqm+hI2pq
buNuAxPi1Z+zOVfezjpPnaeUJPFDNI1ts+yN2/nQqubWjGJGwUQ/rpGlGZ8+K0WEpZ2aUfbWTZqF
AvKJtdd04m8Iv5KNUE/9PThVnM1wuaT9ZMO5+PqkrXs4YGGuw5xW5AoViilm9hrOQ0+A7TDIkLQt
R/5Rabv07alHgyC94RTnqTGArN+hrm2IqJWcZAcqOv/71i+sK/p1dsgcpI4/8UA5WEjFnvJBq3YP
rHZt1f0Wc+XGbUwEjKUykMn+0NogntG22ksmJ2W551E96u8X1PU/Op95cO7JC89AwOUOux6fNEJl
drRw9wJVuz96sa05iCD9F0yzVV1FjjEz+MgjtR0/WIpg+VPgWVuxUMtrtwyiZih0NDBWuaWrFJPh
EUnpnAX+Vp4mSS70WWkQs0f1giI2t66JtFEfM7UxSdRKLcliwfjNtbD97fRDwpwoPvinb/0tVy2c
MFjiGIEYqiKkxOnOkAjZxQBrWXrGRZ8VUwYTEnOagufc9UcUyxq5ICkUBbCJdhVTzJeFfryZIpw2
xs7gsSmPIgL0yy3A9CI3Ne/UtWnyo2A3Dr40R3uuNEeNwq6DSDhCvWZpB5XHWH1ub6hwt7qfVKRv
rWAnwvVBfjNj3563AyefzuDxUjVZ0/DlsskPSgAzph1Hdb7WbcPLoHp50MXBxhQzHNCmmyDB3DGG
duPDISoE5vUXNOLE1NYLhB9XRI71EEjL8jORI6iovKaLHHRmLj0bGpNpG86yFPYkaQuAwb068dOY
qq6TwYKJlalszNRLQq337L69iShTc2ubQtOV0XYYGReXg/vABJe/FqpAxNn4asYRk4c8rfFHK36f
ns2iq7jkqI47s6tpdy/6JHdVjVfLYooUUHhOHHek5coS1rw0nd+XJgyVVyh5DflOT18jzoYsm2CH
3U7n0HCKBte8nMGKyQIEjJHlHBAlxSjzCawgQybDv7/Vv2IxXkyM6wv0wD8LfzrpNv2GfL95m75V
ev4y2RVR3HmN0lL7SOjA1sDEgFnH/g4U9WhSKaxP4gNzdotxAC/3pxXl+80D68EAIq+Xhwg7B+UM
si7Ko7M/AcTltyUi39IrlQ8002dwKsiFuWiXGhCRXBmK+DDkqiSrMvzwI6lxq/CPa9mDyYwExMIl
M10ip5N1gBXhOWKRLDLbaDjg+CAfYqHjB60jFZHDEmRBiDV9ZtTS/FSYg5RRcAK2+5gwhO9j7xv4
gLr4OB5dUWcJQBlHWh2mgBYfAN8CLdGUwYw+XszsiAvhWpkH5dWohMxmcID+gMKloZS3ClHOA3G9
+ARmJofUsG3Nqgf4uv3QXJ17pkRoBp64i8k6K4Q5qKskefnnniK1DpGNAD1qkHBbOB3AG8q+/7UC
dkV0oTEl1Id7NUzwz1ZXMG3acYY3IX90GBXhXnoJgRnb4t4Y/+AMnRssocAHjZ9vLVEy3PV9d8Ks
jOTnMWb5I4iIGgwImZ/4e7713k2twh2eD0tR2d4NE1TFs6XPHlPhB6hWvKlTFHhrWIWYCm9bhB81
dv8m7GyB62lmNw7NLC/o9MDrRUcSO7oa4uwtDjJQ5Eo1iqJdUDgRpQkI2CG94k5JaV9fhV4n0c1l
rZTlWBcc+AEioXX/GeMJteLbAU/Rj3iHSzJjTa5VoPxDhbTQFmfNFT3Ms40ws2KdZEYAz7LKkdO7
g18UA17Zy+vUikcV1cTk/S1tyrc5mjE81t/bKbzVGjFmQL6y4C9qfO2N9zqgbRB16l21o544PDk5
rltstS4E6btI7loRcLZBYgKFumOlMzZElZqYQyryVR9skB9xG0t8zeovQVrJIb/zsWgYqFDyU5hs
BETxrcJewgSZECWkYLahFr8Sq0YznsdzwxuecPsaeE/myASqxEGTX5gHOOFLPYMhc/g8LxaEXeBk
jQMRJvsO91W5JggC4j00DzFxTWXoW7uccjse9Y9ZlOfproISL6n5XDZ2VnZ69082NN6o6PPk35ru
UWaM78Brr85zwI18HG98AzNf7S9Ubhi4rbIVhJ2XjdKN+mMbdFEvhvI2vFpKLTm04tdPVAeEPYln
zEStjNi/U1uvUED3FBXqIWv60hABdUEHSkpL/bh2Tz5G/lZx0X3HHsXQOMqj6qTottkWLoCIaLjw
BsLctqpuROGvFBwXvX/ddm0YIAim5MUMW5S9EajsgTB9dNBeDFSpyZUEmdFl0v/naoYe+mVRS2Xu
6nM8FwTmAWxq1Am3ZdbzM8SZvJxprk/XUR5GFeX/BnbJBo0VxzzUeMuT9PqZEM2OpxNSxM50pSg2
NCM1S3WU7MgGBlIk7bPJEEPVJct1B0EGA6fKkB7las0J2Y+DaXZ1HN6vQqLBSLrNjKXozJ4SHCUL
A39a11W4QgPkLGp97QrmkK7+LRh5MS1S5o9pJaDdD1AZaNPcYPDOnQaeCcL1pZQ6Cc8tFu5JLFlQ
D0piy9jSdixf42HycjrzeZmOIJ7+yZkfJdbr4jt8tT5MVIhkuQURV2qxbPAMJCvRv4OYac9SGcBB
bCfMXevBEizOLMdUu4peQYWOgOyn/RUH9ZSdzOvkTH3Uj3/AqSx63thNPuKVdtiHnET75qNIIQPu
lGdGi4fCh1P9aLMn3yoraufWaC339bvgNxfiST7lozM7KA+wMlm0vyxbnXc+Gu7D1Jm9zixG9NrZ
4BLZSA+m4P+suGPR8vQxZLOWs8JetF4RJIxtH9XbliqPgOeen0z0dwCfAw6ZWoz6D7FOUZOsbT5t
1oMHsv/F1Pt0B61QshXV9sr7vKYGskDViMmhrDVsGWMNCwTJ0v0E28DYth9+16X5SXSaNdtQnF/4
SZoQgRg7mfjYuc//j/CZs2UHGrTgz9KJ7VJoCvQLkuVLN+FXpl/2iRmMdiJHjIeeOiGUif+d7DH6
4mHxHlhE5KJXa07glPetjqjUfUxQz+cVwTI3Z+G9oH4X22SnNjRosXVg+M+b3zohnarZLK1qa0dP
gsUGQlS997kHaQscvTJgjAlrhNM92AA6c61QD3gqwfTang0RBEQ1aDiMJbxalWOT25uKzN4oF6hG
i17Ju5CrP543/qKsEQV/a1PYaKK6REOafua3uajZJDyQvkoyzGj5jtAWOpVdndjAKGBGClxMR0ML
WgT9oNKAMSfZym5tjvAYE0eU1WfpuQBTpufNHfT0erxydhWeZ/xaPQx1diFiYvUxlSAe4FLsrxnm
cz+KemcSrqGcOCEjL8akD4fXEyObLyd6F7SYGUlS58IvrvehCHMnLK5rYGDQVUF5zAeESoh2pdKr
7cF+jqnPZdWn2qkLeyomNKwFeO9e1gilJSuTFm/0OxXeZlVEl+APA1rFc/zSJIlO9hwrkrAVhTJ/
KhXnDp1C9fh07kFkrVKTM0rrLgVNJZ2Vr0eq3R3FakOL436IuxIWJRCBboNuW4Nsrp8lr0DxjvIn
jNzdWZDE/0E1OCOaR7tfRUmd6e0SKmqdoO9tmyrC+Jdx0UNT8mZBjQX7XAdMzcLMa5R23ksy4nW9
rMTbGmHk6NAPsPsc317PBgnccLl4ivW11zRm/KYJCgAZaejWv+eIdPOrUQ0X/awWk+OFGofNmbai
AC0kKiBQel4cURNRTNThRjuoEwcZJ/sV5yOD0xYoXmjPWMHG59lrXmZmJsf/9DiX58ULCi1KVX6w
ojf5rlvIQxiRygpzt0hq+E8OTKsy/JO/leqdnuR8H04Op/otMLV6RoykNciF/zaU183/Fd78zJzL
F8o16c+0Mo4QUbM/5HueOh2cZqVq8nrZRrxz4K92Q9r9UN9ZnPiiC1+Sw33bBG6E0igGcp9Cmi1C
oNCNAHHhgQlAI9g4GPm4lnOUGfrts/7gSpvuHwhaQv16m7PdxUby1Gh1Eqrcopho99VCDUAToDW4
rlDTU2RMiU62RI2gDfI6cpJeUUnwKVsRK3hXaG0tHpLPtoz0U2MdlunDG23EV4Saal2ybG/N8Wf9
tXvswk7qmTE5S2tIZAGB8pEKhdpP/o+cwC+j4EYWRqNfmMBU+jGqgCvT+NU1T2bfoPRsTvSn1Udd
EZRjLYQ3N+h4i2IRpx5KHwawzsRiplhItnNkktpxRv0NArvMp8Sh1Qv4H0Qor7XTrtWSmty++u/k
d0NF/5IDnH+LlWRhdyUPVq3W0TgtAadNQgL6ZKQ9yPlFslJJ2vxZvDBLdgWC77ODM2U3ZmOaqU2C
SiCMRvOJYxYcmD9V5BuErX28DNYw7JqBUfXAqNASQNkmK4E6JKIwP78TuieQWur6VRbma3aTO+c6
seXVIIi04aheDznIsD4CKn4tluIGZ9ziXGoDmV24sNwLjfmaX9yEmkZdMDjJxFXbt29suRHEH6nY
Y4IeDUl1l5tXR89rWrchxfKEt/rsLog/XG02FqlkwEASCBUGjXdEcmliJm9TpVpbJUP+HND+Hefx
DtBkCcmGi+UqAPD462mR/iDCBZZeEDQ0LfUQ2hgS5DgdtoAeoezpLVuPgM+w1GmN7iKbcAMK+ApL
PbD0TJG0Ou73y10B0ZpmpVzZmnxypkCS+3g3k53wGQjkmLumgQ6FFszrnawHEF37kNCYexdtwHSI
S68ACTGmUiDo376ldnMbBtEVtp6v8LGgATJaF5OiDT3z2gF9i3OLIxdFLH5mR0O0g4XNIe0BOI6b
S58WlLdav+twgH7ZQ/rt0PPwMmxM+EC0EogTxlgAMvXVnamNKie1TK246+wN5arNHn70Gm/DrMfZ
lXk6eTXFZ4pEiqPTDfiengMsmcWcVipGkPxAf3qB3UTnrSgV3r4n2D6Nk4iHmJ9snauzb75UU1JF
a/hh2f7CB4aQSgkpG7DqLmYbkLD4brnQ8X+Y5DgRM0mcZ1+fs5rR1F8r4E7SeEDvX2z9wUWFVpQ4
FwAmBRF/h85njhb/jfywnV+DxmLPOg95Hwt/rrNs0bExXuLNAV2+qp2bHL+I+dc0ROvTkMwMsgnj
2Echu1QN9GWj8BHcVWYym1QHnuI+iLDIR7BejDfFH8mhATqpb1oV0O/TSQ85GQqIafp1pEcBfBOz
Qq0GimzxvzsxPikQFqNypX56BjS5l6InkD1kADs0C8Tb+91ry1e60cqCa4zsHUmy+6VhkFbE/HNj
MLwOFh+jNJVelp0CM+TxJTURDSXBiWkxkhLTpa8u8kSJOAqe5kT6SLQF64sLB6nUyGePGj3vz3wx
T/csLiumXEjsNDWAsIxnl4wGZAkhOtC1gwG2lPgS6qh/vOfppeZw9HS0uJrR1q31Zgee18ekomxo
jczXHIMKohWdpJ6HIGxbpkIDropMwfvQMQYTxQfpwCgN259/DVSaK4VIMhd3wTZsPmizT1LfWiWg
L/Ju4WjYAF+nMZdv9ucnN6+yKw0k5e2WlYncqjlfMsS5B82YYZRS043XVUTmLXYPor18Fz9vGgxc
1iQ/gd1XmxMmEHZOWXMP4s9DXnTw1VHLcdT1jH4b5nc9yhGmePnZjghiqnvKmHsbf9RX9uBKJwYv
QPNCUlr72bzSq+zjkn5zS2m9BxdCLVCrnI9vRowum0Y4PsPQE/xNShliqpd0lBl/PGR4M/FSpp7Q
GCe56cEE6pgDWef8ouw6w+5qtGA01zF0pQ2UbFEo6es7Ah+hTZtNHpXh3dQpaeI1N6Hz2B6PoiSz
SVvfY0x6q4BbXAMgmoIr+akY4MnXRMKGbM5U4kh7LEJ+lx1S5Kt/ie49TmvcF3oniRGEP77WQyiQ
AezWCUS+JiP18JmTjXjXHlSfoZCJXfZ8zVCOlrmEMTnCreL0rriGEu3UC611vU/UhZtz4mxdDuh8
q21pK6EdfO5EN4Gc+2MWxF03r0eBgshCxDL1LbJKKf2ovb5bGIFPqIn8gvxVbLTKg4npBiBcUP72
GInpWSHBv/nffh7eDRbeAM9NSrt42vCnQJJo4SQmb5K+q3FMUMYIs00hpoE4hNJqbKhTMM1RNydi
a95ABb6WRfDgcSylr2VkbwAVnGp0EYojJmyYMlWujx5vwU1mR2VDMavw/FwQJ61JLBVLd+CqEJsI
iNCPik2HUMPtibxwU6i3qJ2bNijfM5b0903xNenozgC3bpph9fBXmT7WMSzMsQGQ517Y8FJ/8E9w
tCoztM2DWA9Bq/bB4g6a8jSdRxRvqEx5C5CXR8Jm73YoInWRgzgj0HbxPCJa+UCL/p3/c9ydodbo
BrGGbGC+Ce6mLx86svXuaAQWIQgy/yL+yTuW/RgbfFlBdXAtaSB3zArlHOtKWKI89sCfFDSp0XEM
KWZewnmiwcMkS60QdYMyAx19PxSFEmAvqU2NGoSqr/OLPXdhWwT3lGPp1njIXjcBjv1YGEnsPDJJ
xusAxEgytLPitR8SrlzQ4Ruuck75F5PyXG8C/VvCqi04J3ANfTIei4FoIMllSofynT1s3HLipUu1
ec9GykWpTQeevVgePshuuQMc1IKf/6s0PIG/Hf4wLWk28jtt91HZnRy9lWmWkwGpsBW9teA9SZSL
/qRBgUy79i774e65KT+3Ydk2cDlIeQLYDQHxY2TpR6IYEapexuk8iAWJCBf0tmGyzB2A2rCFe1x5
9mE5jil7AuVf8PQBxKtPY04iL9+ehOwRoROa34hmQsImw/sUQ4wUp6RNUKwEwu4PHl//LlTV5QXn
5iHBI+u4QTfD79lU+dcKbABRfUnaJFYfwCtptLXo5z3PKuXZ/yTLNl4M+iU5zLF5pv+iJ3sKuICc
8tcGbx3DI+JDhN4kS5YeU11/a2Z+KOnGPM61FWVIFgyomP+YhJUKlEw9ws+eLKFIlpwqRoF+7C+f
UB1MnfHsqp8cwFVWVxJeTJUiN3XfdYnfMfcYhv3d26hZT0B5K9LNW6zLRqB7eXv5phnUJoBmPi3t
U+BoIFQpxy88Dq+U6vrYrZ9UJFXb0FLpWTwcPpERiY8NjJoNtm5XWet7H1pA7hhHgyK16Pg3G98d
5welaIercpO+zoTK41upz+oZj1B48QZ0hUUIlUJwva1ghDEeAo+KpikRuDOCWxzGyZ0EcA79SKdP
CysTxbhCfTzQvg3wBRpV4v8KyzFLr24jjBMvszpZ2Ay10KnWiFCay5HVIUTe0+FJKVvnICtPHu+v
9oSkaBhXcrfnIWuejVCE4H8LhwEBRv7GrurbxHWE4+5e4o5psP6dN99B3ShzHkkO7bo4V3M550dP
zTMy8FI/ghzYpB98t2bO7qagftn9Su7oDpw9MJWd3pxMx2lI0eSa1m3iNAP5m0aFd3fMzXRYzo93
keOERwcI/XfYDrB1ZVJP4jsRCD/XYuLSWsFenvgPK/I0DWkcMfH/QsygV28nQuRhmD3U+qfT96BH
2onoxZItjWfOhGnJIF5YkV0ZSqr6K2ibkj6XMCP8sh+tyTfPvXr9Q33iYOvODwV60dKq9oojk4uR
ryVNXroUTQ5CojslWRsaNx9T7c7kcvJOO4fekHCc/kXhXW7U2aEi2tiV1xQnrWgy9sym/2RN4cLv
VhIJD3uQTqqT6KBFyOEUfQFEtVj2WLE++uyTPevLu8/Vi8CJGa+OSOfXVablVE15cN3vcdc94BPt
4UYGcqvj3pUeegc33k/pyJKiX2mMa62L8TbRTdbirlZWJRvci/8d0+wvesZzlnGjILDsJtcyOkqr
KcKDbkxiaCKwlsCXXdRl/xH+xtYEJuD8iW4kuM0zDyl8qR6KNZrvxBivbzXrBXDiqtSBFeA/aBWV
AX1YPYIKMHFrxZ0IGm5RLQUMMSECZBKrPQd7sMSeGQdSoG2N+PeFWWtf45EPMwWK1woHM0FpDY6p
Afsh/XF+OTVT7VGPLi3xfJ5IYhr0++LCHPmzooSK66MiUCidogr8QUtFM36o7bMzscz2gksrAd4i
Zqnd8XbDzGKC+J0IZeN+o7FJ6uEmTzKsQ7wLutH2YIrdn418WBJosvXuD+jdbf28obx1+7PdHGTu
jg+EgRkPDRf432UtCQFap7ztSHeaTyfGhZO11SYzkFtsphsgdL4QtCV4suHWvAfr+HQX9eqeWnQ/
b40AsboDQKqnkcGKfwDGHNlmO3b6fqgTp4XFCKYJpfFL8JjpMynyvmGlNEaYTggnp5i9RmEsWw67
exDQe/oUu01DIEAk2yCnz/HRKjD9g0qsPsdYq/eawtXsyCyM+n1jF1sVRxFy4ch/LLKYVkQoK3MH
QKmi/RO1gLhlu9g9NKZmjILWUtcS/jcZ1a3QWzkLwVR7kXSjRJllCqLSW9jtHPEhXzYnjAQAHIi0
Go+s62BZ7sMvOzrHPzABxwPwGcLhkUwd07FePdTkqhPt8zNGIR2B0BTq/Gwe0qxhMgw5yAKxI2oh
T/sKqlbUq6KAHI1sgXbEeP20+12cvBNb+wLx6DGtK4bE7F9ohQqxgTmGVcx+a7d+wP4geGuP+Nox
OpHqCsbeNtzKdt8hcEIxZOI9GIDPatV627dqQcrXl0iGDfOuGC4ZWFYEcDKtGnccghRQzy/5XAzU
1AiSpiuJk0PODeEKfrprVyxjf4P5mqzLeLJp/cH3ardzIDyzSVGcsUX/vlymfsvoxuC0QLAKbr6j
/kMO5SkQLYONweoXArXnsaN3KTWSBCimG93zoi9u263N4sMQNZHvSo47vixd1gBdZpbY9GFRy0jI
25jhSwAjrFrrR1auSWJ1Oe6c2aESEVwFgaC8AHf0TuNBrYIPwXhq49kptdcje0DvJqxEdO3ygZlr
g2wrob48eu9qJKFaIoKQm8RPuBnNYrR76xUDrg0JbEwryTWjlXwXjM2v2iVYsZBGOkIa16gxL6Tt
A+zfdSOTXwh//GASU9eIGlYKScwDasa/oIXLeEgRusQ9AYUU1MVN6Uy8gsT/2z91RzYtmVtIaRyc
MfKWmw2ZCUyGzFqs2Rjqc8JPzhQU4D5MgbXUxnB/5Cd+WK5XpoPwULgU50eEpNtCB8FriXJoWQme
jBBSBZHvzl/pBtW4TLF6Pwg9WaDA7j+RApfuZNvP/lRNK42TomMKTfg4/NY3fE9IjmnOzI8uONzv
K1YR6V0TaDqxG0eBfAtnx/CO6cqFQfCINWh1fGXqTsTCkH73ONYaGp/I0Dz+FIN0kWcpIIkvkYOO
/JKm/mxE8cOPahMMLthNQOK2YRmGIZDfAp3i40wOytqj/wqFK0Q5HG3LF/RR67dB5gwL09Ag3zpE
LX/iqhjPOAoTQArfjBhfjGbr2TZqL7/WRc7awP0SgLmU4ScIzxqdGiJTXdEjsV3w79s8M0NVYkid
3KeyRbQcBs5kw4ObrPAoQuKLkc1ej1IyDH2RlH9746O6lyyfTN6srzkXb9vWHI43F0kaHJ6nz2cD
Iy0xMJ58FJ39sBVdJCen3S4FrV1CfO18xriDJ2eShe1vyzIaxw3N1VFtP9mBGS46TS0Oy8kK4SAZ
m4Ucg7wkMbDAkn1FjLvDL3K9vjOgJpEDGPyzx6cysf1oNyyg/niQ1/dSshmiLIkE4bEHKskm+/JD
NIaIsw9Q23gNqmd/1wgOkPWuALZZa1fVsWT3sI+5LYq1FLiAMMu4/LfUjc+GH0RfTnzMjr4ICmZu
PTtE3Eq67F3r4lazGoq1jvYAvRCOYDGmwxRrZ2T8GE/qWyD54gLp/nxhQjbaik4c6bXPiAecz3Yq
Za8MzmFIPAe5lm67U+V1SMAD4kn/CX6fgybMG3Vl0WBm7KNmvjMRTYWUWljquJc+8aqg/i+VN3GZ
+IQCtkX9y1tIuY8FHzI6Q2w2rC9NcitL0VOUuE2PkVicWesZ21SugQGVweNW9cv5gx8sKBezRoO6
flxNYMv0UN83wCZxqpX/GiZ+TlYfDsGbYpsch/AQhNpCJYnNZKVIr4lO60LfN+173doVnUndDOPg
OEMiSFOyl2ksF7kAz8omrZDaJ/+pYFZkVHO/2uuMddjB9qQRBkEDtBW1RQzDcUPWhKCMKp2cQJcZ
mY7iUzthrGRAcfutYoOQOMA6lIvbtbH1pz/6yKKsmaz/j5DedNOmcsZCRQEcjgq0I5EdYcRolcKb
ZEGt7B9LvHcuHVswi1EeqNfxjh5dDum03sP24skqQp2O4xdfqtVyOBvyRjYPpt/10EKGdXB75y7R
kiCDJ2SWfJNIKUWlvbN6FLu6QWq72zoFpzbAlZ7mlt5U+lhgPExyKn0KdVjT/uI2hzYYP6dViZp4
o8szEmY3TJoqjj0r5vY/VxricxPsgTGp/nWIQDxM7LRC25SqUMwh5xn0UESZXcW3OAgr3xvTQX+c
5fJttju6txEapFkkzeOTgF2wbL6HoRTnpiSa+IFbjGuSrn3uQndWrX+xZF/hhDefILNlvWPP3e1N
X0ZKZKXLlDwoQWmt1WUS3dnlapGFW6/tz1VHWVnRosjZHGi2bYfCe2jE9CpVCuqtNyqaRqnFn2GB
zyc8JFv7Dk6MpGAQW5W/MH3b1V28+VxbK+CXmD5HzgA7A2bZuuOHEIePmUVLCAR9SpeXoxUYwZyk
BWKjE5KC2QV2eaOjJbdLAJPjcBdnp94eP3Fxy7dAap2gOyQblmT/h4FE/9NFEaamBe1Q0ur2gF7S
OIeo769AJPRNPbFzt2ACkKmtA0L8BtsCqt5xA3gKYggF3TwK5i2/Px3/qT+w4s0SG9leJyJSIDnV
8xNMWjns0k6OEXzSSdql3hCuOQd3rCgbCKv70BrN1044VyboYtdW28dtAldk08XKNLSeL44XzAs2
7zp+KvZ2VrGE987MjuM47xzt7YZOr9xYzmSqKJ8/5giNh2Cg+M+VudRE49/4WPxbP4gBhEsNjNzo
Upa4h5U9VIPbfJNM6FYlkpV+3K4UMcqjOuExbrAHc4+BLK7nky9INFQ4AY+f5K30JCpEe37MYsDP
p7UMML+usoOFZYBME5b7+lY8Ii2iXTlTBK7n34BJbPKyZ1P4DFe5uT0W/aRxv4Wy4vUniEtqRDGc
uRs4bewPBNQIg313C4+R9R6P0uwG7Yvqc41nSqAL8YV4JorgZNGof9mJLBrDVuB4XFzl0phwtN3Q
tUWHCVWp7k76EM1ARTL4ib61hrT41x36Y4uRgkTt6dXvhwD15sxeE+ZLnz3ZPQyZuVHWtHS99UwM
CoQbe5vuLzPd6dRteL9nypQY8LSkFd8Smj4TKT/xjjgzg5VdqH+EFg6+YwCEuXT7Lvwto6cAKaO8
8+54Hrx01rBpS1h5QJ7jhMuyL+ltsyuQ2O4KTS3ZxeOaA6zMAz9t5oc19piYlIVInU5PC7Yp9Mh5
LvhZsaUwJkv1PlvEfK8spbocU+VCt6a89SzNC7qcHCa3fWp3txDd3stGheXYa8w32WU5RhaeJvj4
VrvguXW2hoKz8XGeLhtP/kBJZHMta3lTuR8/lx4pCorGNkuaaRA81IZ1jJua8ulVjafRyZAjXVMU
QvSRboe5qjNJOegBngPofBAogazzL62VdIxdaFhP3qMi44a40J8WLHEiqZWuBz0E1nu8ACaTJrxI
Dehn424fJ2H/4zD6ER1lyc7twCUVapH5Sic9MztbeaoTrjXt5fVinRW7FVmrZ3IdW09QBJaoJCnO
S4URjDuVblflBKgP6xaCpiHR6IayEtoAXijlr9bvxxPlYagkTdfh5psBI9E1fsDSGI0Jn0uo0rrG
8KAli9mUKGDv/OENz4D/riSetLAgFR9rLY6eIhTRSXE38B42ljJkeV3198IPvHPBNfv2G1XXD8/2
F9VAcLl+u8tG+B5NwEvCBTaDZ2mG9xfrng9INClENwEKg/Mg0O/RuS7Gd7WdL459TiCnTMZj1mJN
Ctdq8uIRu8GOlcc597Kx23tsmftKkydM3BVq4YPcZcQL8U3tZzHeoIID5DMyR1GNhcTNa1R4ZriB
6qx9WcxAiAPwotnb6mOuaM/EU5EOnYY+QhUnecnRvOG5Nleo8rMhD/VNG2JB3Dnnp/lkdXdanewn
0fTEgTlbeiWA8C7n+wvYjCmqT8fAR6oausk3UfI+Dd7/0/RmFeDcJAnCW1Xl/p6W0Hhaw6zSM0Ud
3mtTz0Las/m9bdbjKfRXM5vjxaYcT1dZfzRBYW9rZOUBYwoRfyJdfalLOXNWriQ6dz54yme99Fkd
mUNvsNTh7pec+mPW6Kjr2D7pCx+3/R72d6cVlqA2LvbH3GtQU/DWWkXgIeq2b7oT+NWWNZYdha3Z
M/92wOkVUKDlWEnJj4qPwqsobsBZvkQksRmNVUy64Vwf1I8f0JfgS3HsiLNQHsNJUHvI8xkn1McU
ZtNHZvI7qbXa1jm1U1o1Dq7in5GZy5rW5TjRYRZco7pIvlES02/3Xo/am9blmTJJJ8YGv8jHub6n
aQIGHOLNRm5VfcXqVBusr+l4U3IGr9MHMmqV7Xuo0UuA/EzVOVjBa0XMNlzyyhcx9p/HaiJEbcVY
2eYkWIXOj60JPb3Jq69aQUMa1Zn80RzCGCQ0MkMcGddLueiLuMwqyjFQodYOLI8H7hw10OV9VB1a
5mjqeGW/fuqGTo6vCTNkS8upSLaqA66iQR8x6Qax8RRfVgeJKnJefl55Odn6jgR6l2puUySx4dnK
1PRIySWLnVqtC6/gI9TGutg3lnYUS0ezV/+w9K/8mFo+8Hn6KHRkIQRAb0GMU6pWQ5c6noOcrugl
8nhMv0o9XCnl/6Cmxk4EdcZ5898qXQRJMMv294GgBGlgCTbs8gIUC+Z7Q7QygFpgCK/sFrg6rdop
ULvMN0wSyEEqeLYJq35Roz1n8XKNZWZ1K3CaL9j2hS29ZJ2Nxb+22oB7tLkzoTBp5RPnf3yFc9xj
CP1hwk8KRSM/inBiPje30jXHqo8ONBbQt8c9Y8NNCqe+q/nSPspdNcvdj1YpAgBDwR7Wv3tzaFv9
fnhRWynTCG/ow0MQzuso7ZJN54vHvkVnhZ+tXppPVnXwFs8Y9uP3DvKOnw01P1kKvSHxLNXzMtlq
iK+b+CM5HnFUcDmLQfOYn+Kymnu77s9MzdPU0Uyvg6IDUkYm2lY/4WBQsYEDWFDwy/hMGr2XRPUd
lilc6W+qaFRjmqRUMJFzVNFeFgLMCmjT6Y5Cy593joWVysy6HnUakhaOQaoE4jJIye/9wQbtRir/
M8XmW5wiHAbutE56aauCbG++233D3vQIbp6bVNGaKBypwGCv63fQdusofovDoopUAVkGu79p07vg
uod0WlnKZHWD1RniKLRtETCxE3jqb+bgCFqQvFjH1mzJUu4CF7uo4dzUrXg3HFdbwlPZGPF537Rj
sZv1iFmGNbvM0QWGvzjbffSbu+/ObOzhPGRgKNNjgXaK1sRmnNg/WEJIzqPRh//YgxadN9u369Oq
GuGf6279fW993kiT06ydrswJjPtvlFG4dck5JMDwEO7jgQZpR4Vrnc/iF0c2tDLTm2lKW/cJmW9a
Gedr8CeQFzkEOyLqoMN4rue/cFLekbqBVo+P8l9pQsU110Pgb0uG3nQe/IVxNtXfC0qU/EO8qYPd
HPImpSRLjNbwdZ7zy6Ug8Sva3ECDPr+7Wy7gbqtUXZW2kUtM8PwCqc0vj4n3kXmYmiPuvZfnLpJM
ZtSUH7IX+iq645jOHzA4IdvTFBbgfuzzLqOLkfAx8cHVr7LL0Yhjv6jLlYcPuk2B50NTeaLcMIwm
gkw71kC62G2EjMRPV+8KGTTMgfOgjRESIhTP7ZA9WZfUETF5aL6+w72gce8dXLdISIZoKrz3wsyk
Xs9TAaCz09miAze2A60y4j9QmRbc0H2efUbBtqqg1SGmtThTIdWVEPdjUtyTQGXkAm6Dch5Kza/H
HKOoHJc5T3T2B3fjLxD5c3Cyeu9MWMOtvmXac7/TiOtyMrB8Axy8GXLOO7w+UBJSl0ETpzGYIftD
CgyTS1QL+5aL9Oo/GFjwTrW1QfWxywoe3df6YJKSxniOU7UYjHNtHNMt7krrWi6ePvw4hogbJcYm
KPWANO/fN51ozQsu60r6CxfpLcJGDy/937EVmQqvVkMkKz1fVfN5m68Ji6FPBoCJ2ybMKZU/k22a
rDZCzdFlK/q6qB4MhJpgRNBMUDF7IeM32kZ3+DDKxBqyskymupo3XnzR/MQ5KNhroCnLSl2hITjI
H10I0nORDT9Q9hxMAI/Q3C+V+7EFtHfqVqoFnxaPRrtTTaMQbqFjUId90tq4Douq+zXpRC0Z8lWW
BajDWv2gL5zpRLebGqiX/xf8V/kfXS84s2Xirnyvwwor/BdtLFhA78L6PBH1jCcqGl9jdDIhIi4x
e9LTQYUoqwUZvTeHE2h3WVNZHlvrnfQZIF6pIQB4JlqxiSwKyiuAPchz/bh120seS3y8o4ihfbIT
Gwoi30eX40dQ5+Z5RAednn36TahD5lK7G54keDHoV4+etXP+cYzx1ZrkAMFPg7hLQWdkvHW8+q3R
clEWR+W8hUgZ8a9YpArl12k6LCPf+jyAqak6FxOPzc94ZeFHKxi+cIgWSnjjvbYiPhE5jY2/FEOg
EvervGYFhDBKUMwZ6jX6iYvltuRFFdfHLpasHUn1uLKBsfjofrJS/OQk3fjQHxzJRS9tKsWZBKx8
pQyGq9gloIJRA4I1Fh2NlmHMKO26f6WEVsd4o4WKZDoUtBoPQwbXYSJlAG+TnPrF8yhwb3on1pVW
CA03qI94if+f0OU2BboxBo3bYBaTJOtlAqTx4pt4mbUJpcm6hMFO8GFT+KDgAz0cYtLTahXxpgFt
tRyg4GIdv+PGiSJiF/zIL+q89Tw8Ifxc8/cqnK2wgrz2bmtC60k1ZabRAPAW2XxVPQ6oXNWnmUnW
5ZcmsO9h6cQdJjhnQxRaBOHy6n9hmW/fGSlepaw9/Mjz+0ZaR1rfMVjedRNMuvS2cNfFtlyHjtOc
c35Lh477qSBrVufJzYZdaQaJVtoubSlKl4xwozO6AY0rNjNtFbqs+Moz8cZe/xGJ+pFu2bBAofWa
TH7bZn9YACLcmYtJ+mGR/ycF5X1h7ushyk/cOG/NwRA6eH55FngcjLganwWpfOhQ2RL+R5e7PElL
mwM025tc3nByQqsMiPxeYSK744+2cyl6MxNSf2O2tnnrmX2/Og36qYCJdYwhvicNcueTUjn7hxp3
XJ+MuzGAFnPXe+KLMcu9261NZdv9JYViXnQSF0RlUq8JahbU7m+o9kCDilc6om0QBC/LPfcBaPFK
0PWq9CGlrF43qxU7ERk3LmEzdY7u5SYdGaU8DdGbOcHezeCY0524nmqJws56QzZ9ZgUCsX/XD1EA
tsOREBkkQwg2oa6jgW0Er4AJzCvhhRLzWjZW9dFi4I9924rztrtaYL+vUhtwlAkIwkgxSxecc9JZ
jF58Nt0GSmCaZEK9Crp9Dvf527xbndUiFrpBBIcwOoGlPA7ysh59WZJY+59M6nq7JtPbXTFzEYKU
WnetFXFfDlfYUBPm2WHNvXgqYUw6SQKY8o7xYRiYj0sUWg1pqcDqRrWBZjUEVhuqsSggCc4/p61b
cQBWXvM0eku5O8fRxNshxLXwUMl4ndSo4hgvaC7xTluLg8YIj+3MMDMmMpXEZZXG/Vhdmir0d5dw
UJGlzNwyDY26CGii0ZmxTLyheVHHliBa5ESDwHNkRTcMvT8xWerfCvItGQ9YcNxwKM91X+PmIufS
3DZdbzt6SjAEPS6+td4cEsYZwkV0/UZvq45pUPRd92bGyLS2v6s6Z9BnLjSxOpYrOUsYUZCCxQcT
xvjP1J18Xk+IoA+rUNtCBQFtGEMW4VtCUjhBkH9LnKfHs4yxu5RMu2D//uCuYQ+1fY+WFnn/n2z/
cmHQRMzKhHo8PPnUC2DkOkfUCbwQX1VLAG2G6JMzqinkqhc9Gsj17ErWpUtAHstWBvTzIx5m5Ibt
6FLjfk7Wtan5bkPoPhmLTLAEBfOoAv0MlQAb1WfGEQBsIP+yXqm6FqptR5RwT5LPy/QYCffTyr/8
43MQXHmEEp9ueqoyE1sTQGkNdl8hWDx5VAIKk6P32npjh7cEXnEi71J00qxTlLvw3+ypgjUZrDVy
vb5vM8O28gM1yGu11Oj8LmpE9z5OkJ4a3iXyZjMOh2n1hkzvbQWwf+80IDV07ooIOyMSXwsKwWaz
A8o05pPA0LSsRYM0UFEj+gAh2b9mxfDnBpmO1VmiNkyh97uv2tmRa1GXRgwNOfrgfGXlnGbD7xtg
tllcaQRkmw+zerqEFD42vzGv+xA5ba6igpTfzwWjP2yJvUdurjF3cmCzTB4xqZYaNqWVfj84JYDN
tYKFucMu/DuVzPuZUNEiMVAowZVe3gYnqM0Sd3BwgMW5qeFLedfNtB2Igo6XA4DzXhVfe2sQLZk0
bGg7zouPO2PXVg2Kx6GwhMafKLdBrjVBntrI+qIyem5h2Q9BJz2R+F6kseL+3qvoUF6wZ4xogjbp
05NlES5klfVhw1B+f4yTwlOK4K+miglHHscisX36BufpJIG/aWYdMGSYknX3db42I/mFKMZSXHeh
I9S8ebdY1+ry2OqqlDwdR+R9Lz64ID5hQxu/eDn9cUcrnm4+sxFJPuK/LONlW+gaf54iz6q4ziBr
yoJNPTb5WzsZBnmQ8kE0AOwQih4poy6GTQR6oxKBJinlNvEceJjVrJLVkSCtM1mn9SVbB0At6dSD
8b2aJ9Dp2tkc9LniJFGRenul/NCtdsY/HUBOB/j5U8ti0vEAF5ms3biCbU2pCx/337M0BGfCYNLq
pL7vDaMQNHva5xZOGK/kK2YT79BsDIlYWfnrJSXYTExR5ZERCdsTfxFElLEjkyHVA37kOsNSRW9J
hXobVOXIo/AixWafT3laH5/Wcq45YmLW7ZZ7Y6H6kuPFITJlDw0fgAtrgVqwcbWtiEZYZ1+gYBwS
Sb6MWzqDNxnvf+6TM6xI2Q5sZZqTglnAJDD8nrg0myp3sRtXGAg9JFBEJEny7DvmRK3Euk3MGP4s
Sr31RACvzenb+yOBilq//h2dhmO1VV8wSpEeOqcJSZ4G+vkEX2eQViy7Tkodn4yqIbwh7n8cqUAd
4HOlUKqyBGdsRX0HyxEsKqJXbMBU04rMV15xYekZX8qs9ExfvaQOnIAhhXMg9yefaARfcBr90/DB
SxTGk6tLE1bbpxYe9FgqTVQO6ll73H7oxueOeyvr4v0e8IzDIyQRJn94k63rwLOzlfJqnDYLTMDK
s3HeAMTt+xGL1zHjloxJWJ4y6BO3xCpglLUFjws73+CjKIvgVDNbtbL3+3cLYa/bYfGO0DdZMhz9
5vsU6ZEK2sxZgkzAYCUdwTSGAA+f300tDJddkfGAwn3bmxjD1bvz/uo7J43T94vLP7CvK7b6byYH
VFtneqbcYmoc3Pldw9Ko45YDzhO9EHtFyfnqxiHcEbnBaqnOqOvr4FUWw9t+voOWH0UodxheEtTe
omnnXFn/WdfNVEDQdUP+Ph5YmiMkv1AQLAfBzSgZoml5KJ1zaCwl8F9OKx00zKgTRo/zLV3scy4W
MuNZnwPz2qxgXQ7kf9rDJLcqxNIrCvtGPCCD1pjyhFmxQNgD5oXRSStM2RSgHOaGj+TuZyydMlTH
KT8QFv0UUDtPGsaK7DnUOsBgDLZOOYu50otI3T4nNFgtgONG7h/L/rWVPKs2hdCSDi7LiWPLM5rz
AgEeL9/fTMAZ7iV00jOyhfAavpb4lxkhCXyob/1hp8Gg0qj5XEXr6sJdd/jP/7li3Hvl5pRt0Yy2
0VJSDQ4k7xO9JifZD3begtwXFIgDjrrmDeMg4P7A9uJZPpZduD6cUntG0VMM7zz+uboZKQdCZJE7
NnIKx6zDJa2Ky1d+GsMyYyMP+PLe7SZSm0lmPf/edJRJbCpafYlLBBrXqRJlWOK6UqwuQNGYrQzx
eCW2T31a7Lhvz6KSd287Nllozd2USjYF5pduXY5kBza1uaRMY+ucjnQ61EWF+dn/jsDI5L770+Cv
EuxtNSJxKC4HJ4D+X+zNKtolt7Or6I7DtHN+ufXVzZfO2DDc+Gsv3tWBDQQXfWdK/Wn4LSI8DhHE
vvxnrW63zllAtCZ7FRv6LwnBGyvWvJhzIuW+/WTJrBDKMbc/oAcd86QDzFTM649riFKKq+bjAjnV
egEJzVIJnEdiO1J6a45O8irPk+4U1hKfP5ixZPxBdnYmN1mUMOCSsL+QZH7M5ENWzF5i0qUmhf6f
2RNCmD4ojfcrFudMgeM2YUfVCcToj3+CyWgq7Pno0b9MI2JFBFE0QQKZ1lFBaUaEEfOPrE7P3Pim
aatBBD/WrydIQgEY9qCMHbcQ55rt80syfTpj893GsBc8RpNSUSWc8Ozb9Lxy+CeRO09QLRVZz//v
vF9ZJPT3eNg0ugefGCLVe/gJq3geX+O6uirAXAejYSl22W+V1AZD8F4bkPQb5jEQU3doQP8sSIFJ
xH3RtBXmRpQWuukSLVSd6EoV57Z1eFWcop+WrU5KeZYp5zlRq6x89jr755MckYZcwDVUMv9zuMR5
Dw+JCuXFoX1OgqGkNYOaX1WxZV+Nq6NH/JrbETCGGXyIPbzPwKv3c99IBj6gnjF3oDvSzd2u8EG9
PHoeIiTjr8j4nEO2ayEJJoyIPIwwUolUZwCqISTW5QlotACbDSrw0DixmxSePOF7EK11dfElLqDx
FqMRdjt3MQKspyMG+/rUpx9sg6ln/u/4px3V/+sPtOIm1/Px9QoPPKHj7bujhAF7JW3py1vURais
958K7fpxGTIhHeO9Q43iWnxeRDsnvNwEgPMfnJkLNHkbU8riIb1VADHYzcNY2tI38e0/rSDmb7zu
dC9sTNXZ5DPUjDR/SDIexTGlq6qxsZ0JBti5mTWDrB9vUdnxGGCTeyRiHMJZV8iIVhuoISXPkKjG
YYOqt9VlHggHYQtylahN6nThkAuRpT0H6ET++M+gOqKlAZLlZrfUUhuHlv7D9+ZBurfMgvnzCZUL
oonclo+lJdmb+4M06uxHjbL4azStD0OnXP7/f+AscSfF6jM+mjO0VjKFfTKVZJAOAsEkHnE5gwyq
IHSEoMapBkML07I4u9A6EVZKT18LA3ZNZ4cOFPFSpXqT/45iDbcY92st8uG8iErHzn/XKXssGV8c
pZivv/9473ZITAPotaKfETSTy4lsbgI6flq3a2Lst8GLWp4JbrCqP3e23SMJAxtvOC3cnW3ZW8Xr
u9fGacvglGMJSa8QTUGVM3kchVQzzND2SF5UDNDC5oUikPLIL5D678NVX2YrEKXcXT68k5n+15KU
XfN/EFiSPM1w62/i4PJD0te8H3JgLT1ieKEtj8lLzd5eCde/VJKTU8WvhLWIKVK6ZFl24zXUau+M
muNSLa7o8ta9MD2tlCm9JcC8CRnGf5jdVMPFSxlO1NSjmlcggYuXxdI3UwQtQwbf8gsj3K5ZLrSQ
qRwmwOM2IXFhpmKzPRLqwjzVuaJanl9047UdpUNb/xKSzW9chLId2nakri9KeQtN3evzuKAtLO8G
WINatnak5avLhSO3i1VoK6hrYjPHDKmoJgnvvmHPt1lWaF87DzuFFVZJRXx23Rpb+MJz5k3OSimt
Qwq6qk1bzDNh65WErgeN0TKuuGb1xU4+xrHPrdoqrX3Wd/ZCVlLXwXU2zJiYut7bK5qUlzgJJVBP
L/uO4fPtMK7TkBOypHeics5WNqKbMjdk9i7q879HO7ybuRKJiNf+K8OcY37NZXD7AkxYkkM8oqwh
z98x62wPmV+O6GqVKNTJJkxucX3XeRRoEEOBtYEPHOGm2C0NDR+1s7hMbe5akItkvAKmhl4F/vYc
eXzRE284GfIK72XYq0/8GOD2HmLdrPbHhYeGhgNQAcPAgFOZzA/wPWLGnpXH5usZmkKd381zSX5V
IDdaxrDsJriSHn9VoM0RW6h4ZOId8EOr4fqQ8sy46DJ1BwahGnCcL/G0Wzi/fOJWezjBo+1Ka5FW
DUQYh5ucROQlglEe2sgtXoQfYFjnAhX8ITza5YBkbwI8D/tkLuU4SPRgciOEAdevanwQ9vKH93Do
GVHbC4b3/9Ag9wzstKlnWo/hUEuWt+vFC5+BeR65swclw9HVJG0AEHFHv78Xf8R2BjHL3X+2HGxd
3yLpIzUc6YPiozNMQ3SmP2PYrUTiybvZIrF2h2lVbiYTkPIxuzSGKPYGKoSDrBuzHNNZHHDWc0eH
lPp29NKysSvTfDD3V+XXyZ2Lnmi5m1J73FlAUQicAdhDSdqy2F15uruSvACGracz5q7aCKzsra8M
5uGMtmk90jt45SQP5bzarnZdLwvpPBhzqiuvnj4y1qEdgMzBVq8SgF68LX//P5559DKVx6bep3K+
cHwijXxMbsY5MR1peZAhIW2wYdp5lWRs50pbtApFepxJsrmVwyqFJi3/4JnUL0T2/2tZw1HcLseX
M76MkvTwe0l23ur1x0hXNbLg32Ou+ZsEWDE1x6Us9rZhAeJ62Xo0HM+KPqVZJDL/1JPqEDWt7JeN
WNkSE8FGbYwT0sPKij6HlrruSDUSHfblIjKiJAYaoCM3qJUuaSAvWXAXPV7htx4+gTuVJGK3+Gl7
DmJ7tTWA4ieFMB/eX1Jx5TCoJizFSMGUi/mcH6LA3zXtfAmuKz9TuGz9ACuyZBZM9wcUuAqBhW0F
TR4adhEjxhg6khNhXP6BOz4laoiw4/z5vrRgUcmngGDLEvtPTKz4rxsCaAyqYorDcwh9uovBM0//
iD1ttikq5cGO/DX5zZA/3ZXI/pGkbUDh7pHwVW4gjDMk82vJ73URHDLprGQWq8oCXtZVUu5QhHTq
cN2gPKeUM71XyxacQ+rJ6/9MyIuKcwnbKH2wTwD0u6PWUDur0dedexyWusQ1ITuHlupTEfwBe7p+
SaGHkzdj8IyzWrCvnyUMeCx3wRgRKYxzU9//R1caDgv/gTimOUQCFSkH6BPhgO9yGn5qGecXmepO
QLWQv5ixX0VIBNSDU3Rc8xmQ2oIjdN6vFG2Jpv9wbadO9pvSIXYUxfAAiuDk96erhEQ5phmqEE+G
fAxHMZhH2IdGfAJ2/iRPcxusCLlJfmP1UiI2CgkKRv/b6x1SLOCkOQHDocNSpoA6UHQ2+WzKMREK
EGSU3CFQ4FuLEKDveQdEczmA+1E26pG4SPoTaudvxwYn67vTNa5mP5pxa2WNJJ8O1PX8rajaqqDR
nBP6lufxPxnLs1Z71uxMCEVEQeJEd/1cokItJgLsqC1vZHt9mRol69sk00Y6ZTVL27jtKWmhPT5H
acn0muB67HfEc/g8mcKOZLG1vQKaGDm/tvd6PBKe6UMkKFoNADoyzC2lyLJIxcpQX1iyurmd5Bl0
v1ladhZCLfOBADdsIUGET7nin1ULZpcr4RiwfkKaWrp4mbf1i4KwBeyx2crc7ZSOenPuB+EWael1
WzHi8q2OYKK4zu6wXNOgkdBd88D06ypSQRUpZ4eMXBYrzKXrdrfNqodiGqJ6fOSeUpm2H1UfidEv
5LMgLTIVS/LQ0pAXjf4yXjyOySBuxOdRpdTvKHzU9LdXwMk3C+DtWQROlpdfebCNt2kAQCY/412E
ghMxU9sfhtbO9gJWxZoQgBr6GISm8ILAAmmEfwh0+YLHcAEZfEUbCeQMsFGGvxLJ+IWcQWPDWIYF
6v97wP6sNxx6k1xTvWofjLYK6VBNZyRDf17uJTn3DYns4dGCBFaCF/Fe/6JbjU8xOFUmmxAqsUjX
akZ6Tgj05x6qOv6xASNsVbcSAqa5BghTho/pzVI4TYMZ1CN6nj9F5jUgtCha9EgjDqzQe+0VsLUb
5aNhF4pF1VMRli0B9kIL3dN4ChH08kmxC3HnNn7UIQ6/GI6c2DxaHIxXdzpbsEOIiz1kFH1huoqj
ZxfmZp84zwddSgDBz0/87AXRSZr6J1darsXRpEvN42IB5m1wajjStwvdy+SiqRDrB3iM9uqZfs3I
ZyF+i7Sb9KHOozf99xzCYQk6AkKiRPpZStOQGFr//JHphWb5Ky9uqnv9Acoz6p7AL9mf91Q8HKPH
wBOpx6fBwkgMHm/0yZQA65bpPASlnz5RQpqZpWTWLdEwNWokOxBeJcJSLXF5nS2JCMBSwRKjTxj/
wt2pd7Z2605sa4DW4kpTLkscnBQpNbbVXjCvJVN5KTkwuXBbVQj9FEYVqA/HetFED0qE5WU6txTH
r0BnOZgWjxKerAKT8kQN0mpAHCUe10KDSkO8vOdHSz+9YaoAPFy4ArHLRy/SSNsJL2R1g6alTBgu
LstTeByZdQ7Sn57vmdzxVL87LZpLqoANf08yj5FXS+lqkJ5GGowq/dE8k2xN4NLt7w9rMcVFBtKN
9P7hRYNEappQgZSD8l9/WzAXlXQ+vTbiDS2lIF0GNmY9CWzwQZgTOCpiBz4WPTvtQd5NVoOiHPKl
3IXHGzxq9n5YZiKpf0iwj1i5xUEWgV8ZK7N0hzhTQUr68a7BWRjGSjRRB5zXfrud9PVZH/v/u4xQ
DXpIZ9zJuwlpmsR6V6e3+GQlwaWT8QaRK2QR3RhTr6RT9hoVsOeKctwPioG71uYqSSg3+GhRgfI9
6g7mi7OWnYo1dT0QQyvyUb0A3bwuHqKbFaB8z6n2DPHPEQFy2K2fINlCEaSEZKqNkSQEST7Gctuu
1vM7wIDYeGfE3CAjj0VLzlVR6FshHNsxn8vkyCPYalRqPIkYZkg/SSJqwduqlNHKi2nBlpYTYXeA
47qu5m2fMM3byEtGagfdc0yYi87Vty50Xzz0+kg8dE+ZRe87xyE+Pb1VFNFw799hfEnGsLsmQG3g
Df3f3JxJauHJDh0Fx+nywaEzUXzFZNW7D0dn9axTs0nkP/e60eFmfAR1h9qp8AsM+B/L54wBVo7F
RmP0v23hT9M1JROfnaJ/BvbvhizGiC3c7tjDyPhy5+5ModJH1A7zEWexKbTGXGqf4FG/GjxxV48F
mnMcdpOZI+KGfLLssM3XjAJyHeikQ44v3Zhdb1qwRW+vdscJgF6exrfdFTYjXCzrGvVu4V3RjMd/
ubonFsmKq22Qp3o02PwfXbLMTCl+qVJuvS8c1S86dke+wz45maPci4IEXORuzbEpngz5pl8TDsCC
cZCBZKwzcNSzQ2SnU9ImETxAMPyyVAMLXW+nF4Q5g+n06vJ/SJs49TMkExlmSGiVu8+cpeycYbkI
I5xNaAZBp+Nn3cL6XrqEHYAAuC4Yu+48e41mzOlB/ukom9z8C3AW5lQE/ysIBReD3aYC2E73KyN8
AFLeq9dOGhk4cEUNN/WhgbgSl6G3aH8TSbBgV3bPnBUaLQsolXxTfbPhABQBbtIaOHElwCGXq2e/
bLq4I+cXPnmRC2d+gxqTdwiATREsmfhrEI32EB7sszZtPwOkfo0PMSXZmHftLCztYp9MQlv9TXOk
2opfy5D/FdGYaOzJymFQFtk11mTT/4XfAnQWZ5Q5k7XxIrocJcLES7Fcn+2Wt9cpSlfKHYHopG1C
sPXuhz/B5GdPWNpLDYA7uOtVZx+v19rKLBBZV2SA+AAy5/jUSvwcqU9gotlQ5tR3NIcAGD0PNSRx
WxZhwRHNOStGIQBa8HCRt2zOyNviWPtgGdhqFWjsq1r16457dhuVXHMCZuala9d+gO5d+t49sQJ3
Dp4+NLuj9U7DjzmoNAklyk4zXfJwbVPtLcUptsD063C+1OmNQmYSRm8h96wSSpVKSG/PIArhBD8R
zTiEfPYyFDtO7ApmJ3bYsv0tTV6o0jkxPfBIvRtDwzNfGO7s8OIP5XNeYBLTYZyzZp4o99+MsXiy
6OjV8UHhDkrtiJ2iqw24ZObPpZ4xoqbMwaDm7URc3FxcdcI25iD6dSgWylPEBND4MzKXvp1WWSj7
RQhAF0JXu0tXNirE4/8zqYxsEH+t/E40jbVfP4QS1Tf6vxQAFIRs84hMLop1yxoLc4Ck9qa3L+AD
57AS6II0kzuw9OfgV/QedvOiUF7nyxqkiiaCwfaijAeWF4YmNIfUWPUcUwm5JRbXOBsqQO3AujES
W39E5tL/ObBo0dwQ95VQLNiwmubSJuvY1/ekYV54vux1wiBRvkxX0rFmYYo/QnJOe6UIuqTxseyW
6/48xrBmcJQGeCtKZw8UZeObKtWDGzWyKs5Nips2NdzPu8DpfUzhJpHMqkFkbOTiVl1QvP6/PhGd
lAmON5+RRWxLn8eeyG9ObYro9w6WBekNhONmJgJHDsHk/W5GSgn6iY9K0lEyWfcjcsUM1xCCMxAv
i5RWJ3FX37WLN0wYz3UeV4VZazJoqtyVN1LFajDESwPnq03F6TYsRtLrRp8h29ErS5Tdk75yezQ2
DC6+Acw2mpBPIJKZAEdxxVs5ZIt8dQTGCEVqV69oQ/wLwFd06n/sWf/kteXOneDU17t8KSMRWQGS
BQyZR5IiFrYJhIOElctEYWCl9xHnU6R+ddPP0Q5o2Cv3Mucw+8NvJzmDlZAnuGFi1hfKEFJDi0D6
oGpJOgmoNSQynm3Yz3elIzwMmiNVGTIY3SZDPMi5MG9YO7q7+kdOVcBWGT/2SlEFad34Sfv/yz74
ppH5iFLbZjO+TjpkpsdkNTZeLyZFvPpYnEuNnbnHoJaPygfSC76LygXVcJgIjVa6CzjbOSMp7g7h
OWNb6ixZJF9UK7+eiuAC0R50nolJx2t1Thl1U3VcFL9aKcA1wPc7SaoWIICNQplPz5Gbx1kcHNti
ZmyNqEgGj2LkncxVvRvMOEyew7dTph62iZ6FRa2dDlvzmtw5y0kFKRmAOwKNNXAb76+3Hd0Z9CLX
oq4gd/bO9+NhI8b782pKoR+nzmLSMO40+UTRhz6KWDSPjb27WZHcZVcZxoDxi7stBJf8/AipdunU
XY8OgE6Cmk8RRohC8sgFoy+aDSL7PGNuGkzcOeYohYLib6tq3tkUsRwJ/1ruMbV1de42vr0vYahV
+MTJGjbw/7XtadZnBWAfJ9xPUfDsnny2LA6jAcbl0t8gZMo1hsa1wovBjSwxUsj0Td1DAYxh8nFU
HZ2kiolgcN/vfDNypAf/PCKVcdetdskYEYOxl8zk2ZlXMsql2y4qjjzwC2FkiBPks0N8WDg++wdI
jSn9ZmEtujciFxwbDhbF9aEniJJhHURaKbnaas9JSVuD0RiloyaaRxAR59gPaIfdWFmxw7W0ccgr
xJYM6ECo4nuZT5KPMR9LCiaRB8A5fWoiJWtlHXWRvis5Sx1IO4qXq57bvKQMT78geZaFxBy1bx+2
ZSZ3xiGy2ctWU3NWer1ToAZ4ldajPlq/2mfUMN0MClHek+HM+9qb1QregaBDEnP6fINr0Ggm9zWi
y6cxFBqEGjYlAM5gJ58TmnncIVKkv+2Jp2vgDgXoaJAvS2v5m6PcRDpvm8wlW6fDkmD/v67Jqmu0
bHUoJhE+Fz4JYUQlPcUl/Gj3C6enQRnEkMUCHa4vm5oqjaHYHdiO6pzn/EYmy9AO4LzyrGX6ob9e
HiTA04+3dCFRqWLOogd9llOzOCng+mVic7FLhVX1xjOP0mjVsBPdbiisHEKSyPGLVqHMi1uqUBRc
cA76kmHrD1pSdqZePci6tqSKahJwehQAMq9QC7mJWC+gS2F/r2LeXz+JnGHvLzGR/scuc7lU3Nvd
cQn8raOmgbZfUZUYJMxEAjWA9fDlJdjz8ubxsmMw71t7lzFjmWjQ/c1c7RPnN+1z2j9gs0NNFibP
BZpRBd9nlhT8vSpcuiFis8nBuf1fxYaE5j1rh11ZbopWSVJWpUA1+XjmmZMHQdQHEoJetEZA5QB9
WfSbHrogJYiFqOoWYj0xoRjUOFjcBCiu6WYhGVYA/dK7w7TmG0ynURM7ytOV2x1l3FsIHGTd6j8/
R4k2gw03d0AJgUEOPJkrouVxKPPpkmkwCOGZuF/DyLVae0XQw19WByrh6/0UnuqXyMGs6HFSxs11
B4awvjZwmMPaWih0NYfctXx3jPFJz8DiJbmbB0OYwT8OwudTz/HQg/AZZXyRIxZtAJIeZMvBKPNF
XdDLpTFrmB6Feis67HXBBCEH9IgM1HrTbEsRsrg2lYD4O/MYvf0agjMzQLbiMHS5k95/4pbra6ib
vILmoTuKysp8J0wF59ZXJLWrwCAGT+SYSPALhV9khN1o33YD+3C5wS3ZxvcW09NujPUlX5nO5C/l
LkXARfrS+AnERm+mo4cq5VwDzrvxlWA36YkfatZbdtffO+D+NmjP4VMAdo7v1U2lOlUGLT7kFt7Z
Xx68EOZQ9De35V2kItZSfq7/AfjwL67XyiPkQXOypd7w5qg4YkjTfuDLbmG7ukN2vHgK1ulN/3jU
piK0bew7/6QZY7JIYkcOvad5QPUnghVElu2WNXNcHjn8p++6H1cL1e1cxltmnfml/+DBN83AXlYj
71JLe4FIgi0nml/LG2hSprKBjPOVPwcXNIs+qLwyGDobxKk0Qi+706y3PeJxcBHlK8e3S4JvIoRA
8YQApUTZFSJ+EFC1em/4fQrX/QUHWNqsfKTMepXaJzXF2lskCmlRErb8f+lhNnuKiJyvRsGxteBE
MmExoYtuJOvEMRCtid5x12wDDpR73htFjzF25O8sPHVUwjgj71Kqsd7tOM09MWyp/YGZa1Tbdcnn
fb/glE1gMghCGwp2RONBW/1K3FEfi73qKDmcf3Nh6ko8xZ0J0EN0CAvj0kBYj5QnfzbX3I4rWTec
RQ7MjYP35UZFrsEaFg9CS6bzWGfwu8dXb2TtXmlQ+7UL05iyUpqQzVwzQBXzgprYTMx+gjly9Rfb
VxIgqG5aZ+KkEMzgyMvV6+vd8+CgtdjcNQmhRtkNUhofDEyPET9AWBVVUIzxSRYscr5c8MfuA1QM
7K3F79PxiVTIiuaLA/9usMfi+LD84IC9NP4KTugIwetG5g6Q4emO6fM+apIqasrY4RoAY2oBcGpS
EUqW+0CCy8wmIHV0sW7moOHz64zhF5RwiguOAo9SW0e0D+C635icd/cncbffEaWt3uC5A0h7PI4x
JCruYyGhK4WTIDioN3oNxMcBqkwHKVBPoa1ESMpuSTqUcJS1sYwMvXR/Wg5CzZgnzPC1y6xTVy7i
t3/w2VAT2g5Nz4k2Sg8hhmLwwzmeQF9e85NGQ+ahcfebGlJUbvLgrZUGBbBJMGlU5m4j+xo3KA5n
nREmSYzF/sRdKpq+e+MIzSEfpDxzRcPT/CtbCJt5hKYQ6d7eb2I1WwBne1HUGvawfWR9eMnHQ5AU
PB5Q4L5MeDOyYewXFCC2w0ncEr0Unxmv3Ki2BIu7v7tGNnQbCQMga+K5ZMEu98DJhZxRNFFcedkx
rNelS6bp7cj1rNZXmqNQ+u571Vce/Mn7Y3xbKwPBOaR6zeayC7lbXeXhJqH3tajqgmwefpdRMVS+
9gpM+1Syf/ZTdEIKA/ghu93voZy2sqivwNGA7f8OaNPiWstpugk0bYd6lynrXtAHK2J3vs62cIK/
s7TnTSrh+XoKxOZpG3aPS1FY/kO1jrH44H3djimH93SM0nYRcn5AQfib5KpA6JKHM0H/rvuu7s+I
T6KrXi/mw7Qu+ld+gRK5Rv3aNomrPXBoN2oozkt6eECuvept0T6zfqQYg0ayhyBlvhYWcIJhQT3l
PD/zaohyDMb25ZO+avn3K0DSE77AKMl+hNllo8ZShtGQiZIM0E7tKirJkdWS8mWem8pctQVrMgL2
AcJ430ogk+zWM5aw4C4lFw4+zUKWYsUHK5mVQKbMF0TqESvaMlV0p9LZ0N8y1rYXSHiY5PUJFJnu
muY8KEd1XVq3E5YtJoj0q0NcWLUx+V2yIRnm1XkhhqOOB28oBesIlmxDUZygRs9lCRAFkiojK8wl
abSpHqnP/wgWY5MiSMk65xKQcdjLYbEqM/GexoZecw2jL2AFwBLkqjy3z2a6VRxrI26fJ5phlmnX
+XVZpY//k8X7R8ASEzixKU/3AT4cUaWI/EPBU76lknOJdoeu1JeppTP36GzEkOFp7Wgnt7wILOnR
qxiZRVZOlKiIDbjo/kULPLbHspbH7mYJ5UyFBYGV2zPezVHhsUtxQBd624X2SY61RchYhFYKZVlj
7M3Ps5CCuIF75nyDBXPxpYWreArs7MWXadO+7WM2r/GtLyRx5zj72+N4f1vgYgAekaHFd3FmvFZg
C3NgPzpPikuH5f6qsslmYTyHgJy4uhHawGOAWZc9orm1KJ/wmWTvg6lmDls9hYfhgxMUH1XVUut3
m5FuvrjD/b5dlIJq0Zgs6KLNE4/UptLBS8wxfr2k9g0gx5mJPD0dD625Qj9VxFSM7C82mZ9AdAv5
G69JnvjoC1jYVWqMe3JhfB3qmofBPcexSLi5X3fb+kpdCu9/fh3J7KQmFDNR3QfFi+F8JyKNEV8z
yyqPadzZzrycCQNFNgaWeZpJPkArwgNJeq9LmcCl/IiIK02CcI0lcgUlGfBIEX9OB2KTjOTAoAnX
72hKdMG3cDHNiR7teeLpl76sJxmt/yuhlJUVQYO0Qq8gIePo4DqQWr2zOpIrAgrTeXczV6V0h/P/
8jCdUvYcOlUcM1nILLS8tSRIaDMG3EfVq8ABUDDR8AE4GiZxqDW2RXkHtl3jtohG5QZkQPfRdwPW
3I06mxvLjQHa71DNXiL//Yh40zetZIMbE1sNMyKTGNWJhZ1e9R8mVcfNlMxeM98RUM0DIg4oQh5t
r3LuBrHphR/fvqNeJ0qcKB3icIjvMP+VbfG59xooJXtHs2hQGhHpStOj8Nx0BhmitV4Il9tAp71D
FrsiCaKXBp7E5N675ePcZ62V0hN5Xd7mQMEv1qiLsGp4kzklX6gLp6rZm4f+Pim4MQ9Kzxa0Ls3P
rCnKqdYinJ1QK+RDRLD4beY0fygCYKkeKYCGxFb79PQ1/5WdY5/gqgOpjhNoIzQXCIF3i/OObTGA
28efRDCQutl2GBds1C/0C/6wJ2OxZemVjwq3SsGnqcknS6iay5rF+7itl7zVC6vfiTfj2aXhrAny
+GpmztRjLf5AqLUMUe6k4y1VO/E9zSO0cH/TdmtXwPlfDN1rwYpu/5sghwzEynERuCIU7p0EEAmJ
/NkWK11J2VGVMJemrmQMD6rhAvkMCC4iT4voWMjlR9Dou5JLzCIrEpTOojQS3EGc9uc+9XovOPDl
8a9ii+2TtfsJJS8rN7MlRy8UNZ8u5vl/8DGT0wyww2NmSOqCRj1okV0Y3UZ8TumKmpSZwFooIevX
Sj6/HHkwICExQCN5V80vNzLYwMA+00LUfC8eFbQDBlWfUnYOz0WVggvpQeM7MMIlKqqXmMU5catM
m9tYqc3i4KsD/doEuhZAsT3UO63czTCyKgZGY+YyFWfHRpL80xu6fqItKCHVeLEJcfKuvl2yRlGG
3cjoh+rwWVX1eF1mO1BLfWWx+uzUazDrnYhViXqm31Hajq12Q1xRqWLPcuDw8Prx2aBqwoXBvuGt
gSpNIgag0Kbpsdx/axTTR3gswiHZhzM2yp9QbMegdEp04cItQ0FYh+rBxEXyNsUVCLCiswvhovIh
/vE4hb77wOUpdqh9f2SuFtOPm0SBZojmsqe0oW6uhMzEAdFpV4/y4NFRBtx1InA8mbJlYIYQ8SJr
gWZEDYlfax8Q7umjWSWOWoF/2cPYOwRR7lRwK/1HKIjrN2AoGRrVVPs1Pc45KK4NgRZo2BJPXRho
6l1BSibP/OqHPg0fcXX3LDy0fYvp062JUIBmKY8t8Fjor4HRG53JQIWX6RgEd11ttYgM/vD/EDsO
msEiG4DcFoNRxuEvnIA/GuAug1De3FsK0VV+C/J7dMSuiyc6oBEMx9gIlJmn4jJSwmOxpPwf8Xec
wWZXeSfCxmcvpKVlRIm9DBr0covZIIbViy/N+/SHuFYJFICf5NcEOG6iEgSFPo/5uVUZd8sltxct
JxatmGlno5nl46MHXKvlDdpKZwADizUB46+SSjIFC4OJI60sUGpzRv4mb3JUrArR9Imm2S1mrMJE
E8qMwPwUTQM0l1I+ZjQGC7+PEvdCpCbUqh1+efQ8Yza4/EOk7qDHwxduA2J4rhQLn32dr5QeGd+S
BadFhTEbctnI6i3NGIHQPtVo4vM7XxLKGYJISGwkaiZJtk1dhkeAsdyYwa31sAy/IxFZkR9p9U48
60VAr8VTzj9IjWXCcYHctJKnp6g2hxrh1jz6/lY5Ea9F+Y7N8J7GSrvRUU5vsVZpvTZgYAaWEonK
N3gaYFWXTZwIrsci2Hw7L8kHRTE+865ZrvNloK1zDaiQlsMiQnAvnmTL3GHEGN6zZFrh54vqPvAr
vINQgX7X6/NI+lhObLtA6FLv1ZETdPhS8lri/o6lvMosEE9RGld9yiSvmB0/v3owIb+1FZ74Xke5
Clf77wYuz+XqyImbV4sBpFPb+Te7haF+WhXCWdTzU+pylW/r1tndzsW/JC9H69klNvXT/HmSxWe9
eEjHfIsU/8/2UzIrp112+1rvLmPrTvGvnyrSlxx3jxvDBHnHPjy5GQzWERWmgrCrUHXGqbPWMcOQ
yIGpWxXh8z3Z+IVOVpZ6G5siieJVgcOkxwMC0OloiTIEVsbxjjLY+BlCkOik1wGexdwN1uS0yURC
rrn9AmN5+ncjUuA1r6pRMxfyomIPXfQ9r+uGusQbOB6romyibszFFhuPJFz35JterULZDjDUu6MW
caAqsQLKJCxvxXmyVW0ADb1lrWVOUmHzQCe4EQNDDDhztE4qemvoXBrw6VKmbFCWItZN6G9wPVTu
PeDnB6ge6k0aJoHbA0nvwv3L0dt6nCLVrIb//JxgSHQ+yCuwR8Ang2kIYVcBGSDwEADMhg9+JdeM
Zi80eP7Laa8YW9B/avHJZWC2eMHsyzbRsuIkkCCoH3//CENcaPU+KCKN8TALMUSYm2v/qLN/lWpm
B5mpydoxIiS57wWMF6/U/8wsed2rqTHRdstrjH1dKCKM1Pnk57ZYyUdcqHFmtMi3eLQu5Iykz1+p
BLLe8ooreHHF4w74DxsUQ8+mXbhmYvvWO0Srv/euPjZQig0cbxD0lgmgfl23HBuRutsLIvRJiXre
bz5FkmpiIImecR24i46vN+CGOwOX8EiPsasr7nsahKRE5muT991LGfQpXb8Tr8ZOu4ctX1jAbmY+
YES3N0ZgnY/eBz2UIWVF9yj/1Ozl8PY5IO/H3PUyYpRfMcd03Z3Dn5C6M/EfK+U8/riHgd+51rYx
jx+377ZtWGMCNBuzY5t79r3cQi2E8IZur1xDA2r2Y7X+bHMZsStBpHo1Q5ukgxTRQIMmy2FWOvhz
lVuyt1d0EDT8K2jeLzKzVzoLA7M6YyFSKR6nNRRhakNobqFFmDy3mphghq80P2P2AoskwRyYuXn2
h6B+e4RrKX1sx06hiIcDWp7EgjWK3cCw8sqRKzBl+i6/nII3sfkUfhRyrixSRM8rU7NKTRgzYgrS
ucYjocScsOil/nt6NpwtoarxakPT1lPihI2zqUw4AUjW6rby+qJDFW89/un3ojFLRzYHH8/0GL7d
FGyWYKJPIx/x6onbtgrlCclapoLXC/sxqNY5mOyymWsdKdu7R8pps9Kj1ZAz1YO8kBOl3pVQlzrR
FJAIcAgPDuqiiXhFh2hW7HkDNcT+W28u1kJJwU5Fx5rxpI1b16BYfeKOvbEpWKHtaUB8B0xxtZaA
OU/EGc9p8yH4XxF1Ayp02Fi23At4uSdSjvpa689ohkE3+zGeJhOizPJg57/o7dty1XJLNzTxgaN/
ZHG1QSNo5RCaYcM0smM/AM5B1HdnYw6nVKWDixIQZm3DsoZeEPGjYk+o8TYHNBxY4Obv3UN6qk2F
5lTjahuxRGvgRxK8UpeukSZso6ZjHfz+kOVaF/nVktFrYU/hCX1G6ey2wDAT0EugX1NZEssXVkjK
lZhIYPo6HBJdGIVxZJSZ+ass+DwaFQFWEgMyw636ZPZqRfon8PwOcE4rIlClgHlVCI87jJSmg6LL
KqjVlY5DBdebb3EMlHX8V7bPVqxYKVRkbDeI7JzURIeJV4N9i9gKkbD0HkUIF2fdfd9VdcQVu7Sd
R9YNvAQ/FPq4Vwd/Xi624mfLU5gfm+c5+eZ1EJ47yQDA7pqxNeXnjgWbshiCbzLjd052oPd6O2zS
IjpA++QI12GXdhqqmpTTwiH5whT3ZVi1ZgxEHiihtQgNOXuH0zvWZJp5DyAP5hUKXOkxSHMG+BrW
2T8OauK7kqo2cn6lFYy0p+ZPAaarWoxdgCs/HqbKFBpL7HtFdS4vLsMCY6yFNfOjhxg+fDgcj7Xk
N7YZEhu9aGiaTeqMWNAwuJF4pCuYR8T1hueYM23oC/vZTw3gveChivhT8VPmBeIcWIvdB9Nw+pY5
AReKnWHD+dVMT9DNkG/i60z5nFhZjQYCniHodT8u02UtYh7/5KTeyqP4gN8W8lYIwvrcnn7qlkZq
gEBZ+DJ6gM7IXKTvYmZqBYxhGhN4al0E/1BHRxOjq3k8YLVeqfCutj5vSA0WZYmKwrcHNa3miDM6
3z29XX6xbxEGmpik9zwNw9nA8R9AIijY//b1x+a0LlY/2Z/bpaMlCcOPm+S2aAMyS0Bum4rrliDl
t8JjhQzqGMNsoUdpJRi6SJXtxAZrahob5N11Rrqi7rVYlqd4r412yqss3+YqOaKCX2IkgS7+Wxqv
lG+HcvdoMZx5W9gx71NqLwVeUipBCD0p56RTo2JH0TBvwJt4zKrb1PJKLym+67luBRX8TqIBgDz9
2+DZByxka5zfdrOtDVYfrfctvB0hfQVEljDVl5bT5+p/A99XfXRbfuk9ginra4yFWWkM1mJ3FHYO
YE75JJ/KvCjq2sCyrxR22osP25A80oIyckibrJUWTCD0nwGsymCOJZ5EOcKuw+1i57QC9T78D6i2
P1j/637dS0qkOYDQtC21wACPMnCHpBk9BEsIEFoPuOyJIDAefcy6lp4r42xtEXWja2AWlLZLRcBn
mbO+ogHqS2kXv6DedOclSYG9SEKjYxK0GBg5ZOsCWhEpW9757qtsmdjPog0sLrepTZiMMFtdnmvf
PpihpQmdpJ3ilB/K4YJ/4MXD+j58NdGshwwyBdJs2d3W92maF4eQc68G/FYiSrohUXqz05hl2LUU
0evgun4xWvljIcVRrj1x0IAmKbnF5v2E4Xwdt2a2SO3iMB5cPWzE1WuaXJy3p4gs2HUbQejnS2oZ
9gX98Mo13TdRcgH6dj+K/FHVhZ9hpdK9uE9lTxXhqjvFYENsOWbC2QDyGVVt8ErEn+QUAPyzgpSZ
u2agapweZpVoqJcfGE2fT5ErSCwBgjEWl/WtFIr1mt/0cbx6P8m+ejmRbCk5aYj0wsUG5ZDyUS5p
7cGzz8B2pm9MrhX0fJ9qFAFRa6U9MXsqTtwcLdHAfB9MKgw1YAvTmIBi+nY6W5sxyJprCdeK2IXy
FgvlnlekGDbonV8gMQf8EbaNFcZt4BXekXzD0RNfaEgoFJQ1qnGl+pcDAXFkRp8MM0YzR9Ul7m2A
oY5H9p86Pxx4R6WH1UTp2QrTj9/rXgHGWHe6vdwL644cFPXMIPDKSaDWQ2BmTSYtqJl2XytR0kyc
c2oSbheW7LzOi63ENJ6CPwSszTlW96+gGe6kLKdWkOGumvvPpD9hk1tsaS4XtdfvcSkah9/llaiP
ES9LTfCEyp01bvW8wOnWgHEyxzkqeVeboZllUmWGMCZ/H40xvQNXwAMwGtSGpvhht++nwG3LG3U1
JVnzUNIwwNXs+NgJTtogv645D4Yww4+StpFwZGcdUNuoVw2qoJjkIKkdpMUm2qsllbriw+O+tmYO
iZSoxMjiZ2are3xiClarM3dUbcvUlRn0nIywK1zR3ikdLAgRLZke3gmeVY75HsUp0bw4R4tcSYvQ
jWVof+k0u60huMG2E/Lhmqin4fDHmeOdN9uxGXd2wHk/dxE0WvHxC9R5/p5hszeUjK6rUM5d/Za1
JR1hXI7GULsPyLJ3cYOC5w5JyalrSwcccZ+qlwtVtFKme6TWCoMTo14fnP5sfVWnN7+AIwYNL8iT
i1A1Mr0Y6u6lIJ1QlcfeLspTCHYhRP2r2sTKjHCG1oGk3j0pO4zWy0bLXFJWIOL7ltC1E2hC8zM6
fHxpJq89FN9HNJwKNbsPtP+IHRnTzfDCNV/hTtkqU+23JlimhiUp+raGsymF5JNUzn1JmqgFJjVD
ljgUPlB7JfklgYQy9fCMhb6a8DxqA8xDb/V7IV4aHfe4kur+F2wMb41n8tZLRix6lsppKyMqR2Rl
MKsw1vQ3anWI73il/QDC+5RywCyGkZOkJGUzhPXrFhVudCKHjVAue5o8TUM/GX/7sFczk7Z2rlIa
FotZUcS+h95M+7pbCklNDMI55fChI0kKmPNURvmHttoyf+VXiBnyy7ksF69SBZQ9QIjyrg8NyBUz
2DkTXhy6zEjSH2QOSJeCosEX2Q3hr4MMAw6LdBp8V0PIg+dssygc6UMZ067gb2q/vm9jAxXy/5PC
caFVmafQq7LwwcenSspIbTZP/3H0C4PtdbWjPfptFKYb1ssajIFiVw2BY/vo6w6T0J/fWtgB4Y5r
i4PwldPQSdasY08TVy6f++HFUJVDFm0Y05US0wcitm0gAMi8Hie4ZG3/Mocs6TNPq0V31/pRJxMd
B3JWOb3Tx5xyrk0V7CgWvuqlOGEjP62k6Xpgwuvbwrc0wEM9QTgYX15/GvQYR/wGxJ5QQ2XWGbER
cEaGs6xQvXWRYYMxJcsk3OV85WfZPDU/qhERG709Bub9gkbaKSPn4KV9fyKppXTU08355GATUpzu
tXOjJynyPOCVS/Kl0m81ck+Zl8Gdg0Ud1l6H+SGncPu/GUsqAFLJHpyaAHr/73tLDSMXWPHg/oNm
DkLIXnQ2rEkD/sjpl5dSF28NYE1m+XDn2gXyzVk38rHiHA46zrbhOhbRtxsNLkC4JVztXOljkFGQ
JppjN8MvR8xGhALO7FuC/BS52pNo2fJcvRn105vQeCeBXZa42E0HXjdGeNAEmYkZWEsDNtg/T+7j
Ebz5sUtOp+Cgjx2KDlXllMyohYqrXQ4CU9wKUsECH9jX0qQYvuC8DWQ9IGcDa2BHpxi7E4NimWwy
+N2FvTcH0wArPJiohd4JqY+TIUC1rOWUqYqXUmbfosOaap+TcjgdfvGFrX8OfdKZ3raA8vkOYPo6
qVLs9C+V88tf36p03Xw16FUTlpbTWvmVedel8qX0GI/C4xYjk6q10zwiDwPOlVaItcSFuNm3sDym
idTwMyN00a0cbdg9kDX4WV5y6LpQJSazhh0vqa6EA+3D7Gr1p0xSTpZ3+vXF583KWxZAWaUsjjAA
rF6RzOacos9bFm5WPj1ZYsFdPoTlyGvJGcqzC0WoUleiYbdHB5wBcXP1vT1lMRfX/jcjGydhHLPd
NuRvVXsxDAOqtL1PdfENRyXhr+0OArJQ5EQ3JcDaR/nAM20/TtTWdyjfyDj7/gj//oNAqVG0//p4
Asa1DMSwwb5wpDs4lq/1acoz8i3HRR05LpZmP2hHiFjXe/JyF19mojRGHIbM++sF0Vte6wMsAv2s
+WzhB3xCuA8WPJLDrtAenTMXhW2CaeFUm3h58as8ysphGXRsJJcFxksFTFYqVVTvCrL2D7sT3BBs
byS3lvYLDwd12l+7yy+sb4Dq/dtln1rcLDpcvd4eKX+rVD9q1po0RtCDahC0gSdqPCLz4I3WhmfZ
8mqqGWrZqJFI08Dm2vGgA9J6KtVqeajG8e7yKdlCQNQHLRHqTDLk76rGxyBAFukl0n1aBZrTd/hr
xk5doga9glFgVho8WnqIzZ3jPFASVrtQoZMW8lB4l3Dhs+2Z7+1ko/ak094OnuI1EtSDKbTbzPr2
g2cTsM8DPU+iyTQ4iXRXfDHMLezmZ9f0yRKl33KkXuCtj/RoA2jChh7po8/LH4e0tr9mQ+yH+Ljv
JoT3uapxz2CJjTJ5qQiSyZsSY10qKyY4wZ87jXH/ApHa/vQOPGTntr1ZgOJjW2z5zNlc0ZXeGhoc
DCWrsv8z4hTqkWp6DhF2aRUGxAfNokkcxCqZBhJC6DL9cETC6nF/ldPwfERRJFLYBxdDHULM28KC
rWlvwJpeG52thrGSgl6hTUqAbexne5/lw30Ov4UIH08pMimbtUXIXLsS0QTNkCA4eVHgky5QVqX7
ukM2RZvR7h5bsZNqsCFpQpm9Tav7ZajLc9S5l1WZgikPfZQHpr2iITGoGeR3KHRimpMJ59HPkaSc
QBVePyL2iRuColF1OnetrmwDO1s20TzFdi3XNwZTGQoAaDjPE3HkZyze4FUv0peegu/85fITyCVV
o5wpvN/dJk9cgjikwxNot6UxCRR5K+Pcv6WQqWqL49gbbf8AB3WVKfRXi54OgaRC3GxyZH9uncT0
xwPbX+mFm/gulPwjFwBhPOdAoafyHW4KZT/aX5e8FP82c83wsNUbZ3pD8TVGs570hDg+Cdrk0frY
O1QCXLMPVcYE2g1MuTR2WDFXsLeymuPVyqh4pfnzsTC6VVu8etx7w0vp6VcIVuZpVFPTJlVHjaL2
G2neAC9BuxqSjg6Dpds91AvW5y6kcAKM6zcEly1tAOtTt6BXzji7UOJVINNQGs7krlB6VozRYSI8
k3hXMV2MzNGJAVPibocjgdoI+wmhL5jGhabasFHLbOWtjLbSm1JLduGs1zIVKiL6d1ClSQlFLHpQ
ke2PgnBUZfvaoRhQF2HBhiskLJORcTHxc04UZ8AQcpgG+xZVmpr1E09OeApoVN9GUdICmRqB0vL5
d8VKePFoJQGDKubOO9o7XjR4xXy5haomCWBJKtwzoAuBYb1UnT1RzAkzO9zhaugNjjIRg0wKlTDI
XJbrDRc1ZQpLWJ3KpE657drRbu4kisXK7NBTDVQiBL8pNLLF/Zd23cdX8mTBoSdKzL9iDg2a9yjI
PTlZ0m/pUPRYadK1/e8gMtZh1dW7I+8+LqMl0ha7J3bDTh6sjeDpuYb2xdmI3FNDdCpKxXGtCE/A
sUae1yFXShIQ66omr3XEplLy+VMKgPu/+1SPBG9PNQskJ2HN4cDZtjSOhuJdEqI9kIpAfncM6m/8
YkSxvyf0QNXKNDPZeIjksTifvaVDgC913kaJthg/x31g001OBRdyzVs4V2htCL+YxZT0sOqrV34l
qdusM8AY1YmaRabN7fjOSXPVIKNaPCu0IBkzoB6XBzPBTLnAU+W1DacYT/IhABhDFDjTzJQJalYX
vL0XedmaeyxExbVhsFm+HdgaG2+9CulsK9ghcL6ljelwoIjZCt5rekB2bUuf7gE9XFWlbc2m2rj/
qhoHy0XO9Lq856n93m2WuUXJ6kzUorWsk3g+zjImpoI9Jx2Zxx5MtJ4fZ58QAMlks5b89FfkASD3
NZkWAe7DzTUTVcW8mpKqHPGCWHLoiCyfeWdpaPg+nXdSYnh20ynzJpP9dgy81mK6k4O0CulBiJ/y
UYqo/wPNkB96HrXelhVqRy9tLRgvtLwooqAsHc0MUWlaAyBYUUvyVuI0z9BiMQvlSvsUrIUSazkT
u7FyR6TIJg+WKloUmm+7uYwcdugxkX/xmv/GmBrUkmPW6BLxYdcWGFqg2YEd88Nl0FSzaXspznrP
f9yQI/vDhbKbTMFBq6W6nNSnmcEKgd7YOMyuaOD9cOCgpJOjk7dEj2xvWISU8HFFYstCLuqPlQ0Y
JhvV7kjTkUouFrr7Qnt9NB0qvMUjJFVqWeHs1f3GydsC2f/Hod+F8o5SJZS9Sr/lrM3OAzQozCGQ
syLBtTqYHCEDAhevdDkjWTz3/yzkXQUKdHB8XDF0bzIliXo8CoIHIrTWVpyxrR/h9IRMoKlZ1z+G
Fwoa5ewzod4asvTOpkugdZLDBNvXjsJ/Y52UBuQXw2lM4FPvqB/k7LGoX2mC72cCXImRYroTEoVm
v+9c/JEWcjNYWwgC0gviMVwLkhzlmWq7duD7qKwU0cEj0zkz0+249SH4+TN9XT7e2a8uKHP3hXSW
RK7/CqmPVEmJVYUGxtiiWxtuCagYVYsFbO9HqwLHf4B0r8ePdXLJpWjlj6EZGgsxqtjyWLG7d8dP
YtpMtviiNj2vfSdSXpS6lbZr76SyvqpgMcNBlb+uRmCPpfMcV+6oKeZFUz2nlefa07rp0Uz8seHB
1csrXaxuTA1/2FV8gVP31JDfeayuxYuR59655g/AKlxxXZU9eTRAdJKSfrtLfRuQq4XHYYOy8mmx
YTfrwgUI5mUFDJWPhhfoMcdyRQb3xYrHpVGWLfdz8Y4+0gK+RHklImSoe+5w8hFZXWISi420bQ3p
+c++IMD1avrbBZAHMaQKpwKebtjyhgdhmpE7OgicOjny18cP2EOoZXhR6NX0ZxhfZGGsynb6TDs+
eK+OxeZImpheyfTYoN2LOnuAMN6mNqzRtNpOY2U1YWmXPNnIFRrFFFk5GJgNBeCF9gZTAdGBDdXw
Aa6VGoy1XylvELJkNy0xC+n93PNoYAVrWlEPBXQifxwOhzRbNnps93fi54+iaGU/+w27KtFFQmBB
19FHXIkUZmQzpA10ruQVvXovmFtCMWr6/86FBOOcMLSbtQH9IzPWnvr0v6tpuQmHzb2uvCyGDf7s
COhURtal4VxWNAHP5oGQ5NVcKDxXvnCeWtyc/sO9dqYIgPHMjDPemZw6vRqIlgT91uUUp71Kd/mf
bFGludrieUwZ97kvZvqCfNyiKFZoSivp/lH+Kiom1/yffJlf4LiHF4crhoOak6B9yP6yAmhuQXHd
x0BxfUeB9xvbp0tD67V08cPo8OjIkop04WsBVFbG33cIGqc9wf0KkCau7W4POgkbAh2ip2kAWh6x
iK9OiO2lWquW/NaDTc7aXpGl48MgdNrhcawZNKlOyKmFqq9rvSUQ5NTS22IcWbVUUUGe4RiJmsNW
c7CINMg76blPcLTK3fxNurOBCcmCN0f07hOxqlXmz6l72adVLJ8wRKLjRg+Hr97KkMvt79TTkDrL
6FrRb+b7OEVZoC64/HFU3v1prwq1l8/T72kUpxUqA658tv4/CDSZIWQs/FBGjLGxXfYQKxt8GZ/P
6Ipx31i2GXDLJSZAFnaLn0EcTPPrchvwUBq9TW4H2ItaDiSTMTY6vnEzrMhVFCfkZ13htfUqFKFh
Rqwnq6UGO68B9mLRUOS3axF6GfiCqYBaFh4PtHitb4ltPhiTkAR4AMf6puwI6oGiggfkixeXavNI
OIXEwism1CaJK3rfJ7s2STezSS2LY4/gmQS1xLFE/g1/3Hq2gSMV0wRT1u2LPp2FaDQFSTrk3Jj+
UnxMESSfrOKQ7UDWUb8n/JQvMIa6DLzIasZ8NaTDzHrYOIrfPLAfLAqxSfpOrpBQNMmTiMe4vdCy
slGTQKhdlq5h4cHDlipKayxicS5Gs1jhgMbCQ2e+1Y+s/jLICa6NG2b4Qmewk4FQVtRwtfR1GveS
niuUzExQrabPGbNHB44s55Qk98yQEhI9TlkU5PeCLELSXnd8FnQ5TslCWQvwIWznbLTpHYgJCTvq
p+lS5A7GCiGiifEC7lPr9900wfYJIN6Aa+bzjAC/FZdUepuglPyubdHdQhMC1O4GjUaTMC9CVbqk
j7gzb7718Dz9qjlJD0WMyao79g8UzsUedHDvlXcm3elftBG0KIEkEuwiuBmvn9m35n95u8KwUZOK
UsdWZAamlgHm85vvFo79B9f4dVPB5mdM7eSnIh2kjH6mx7h9clwQAV/RtlU3rrWByb/ObiigXuRU
9lk3Y592tgznwc6hszP1CscLQkCqjmzjH9gwL/BuzAQE3FM5TZsAWRBa/qrynJPCWIwoBclTRuAl
eqmC829a6X4JHqPr4aB0GlK0GHXry+JhrXZid6u3MosZUhA6Eq2y0oQ1jHsl0zFWnipEwl30KlN7
r1usskn3Od3nuBYr1Iad/u4AwktLYrTDQa0rb2SEC2/4Tkr5/JqnVZ6mM4O5/Hoh5HQLlxzdQCQF
lj5a+MhKTSR8T46/qNrUzQjcfQf+2dV5QuuK7qt3j9nf+893Yk/5tg+sZOoaBZirbzKm5HyWc8Uk
4vgJo7rtNorO5+0qosI7z7vgbRDuWxPGrnKFsd5YTr1fFi6C/tErMHGZgww+txj0EczOZlyAkdWZ
7cvY0HzoxwVl6mbWUmqq1jTjvZ2Z+KyjNYVHSy9Jwm8uudRUd5rq579259upotcUvmGy8whe+7LU
7hlVCR2V3uyyntsLcVx8I0ISn+mTryHfn4Fdd1d4U1VBxkZ9+FXy8bFnbr6hEe30LeJCyGuoWhnw
Q1eSzXH1FPZgj329b/YOAfXEywMdQfIeeTrBHRTRV3CxTzwia4m4pv8Q0SAedNCe5OdEFM4EhEC3
rndmtbWN5DgmCYOksA84WyFkGhBBkD5PLkKnvji1Ue3/GcjP97EKnvtjOeDvyqmsxINa6ekl/BCN
aH0/85yj3fQC15KshuaAd9RpPM7rMisABnf0XRvxQ8PBw+skLJpIIiML+BUDz1qEtWCf5/l0ldQU
pOU2mrjbxmWa5txhrZZyyRDfgb/w4/VAktzLkswCWB91fHzhrruN8cn8CqEcjzx/A3HYGJrwVGHp
eUj+jLi8FOfh3RwQpgtyUUQqhNztn3htjOoveod8UAT3flNsqyo05CS1aPewT5N9EJ2pVLtBJ3gP
/3JlDtwzP0EpQWURR2U6+j6IHWslzL9LOve7+bJosOzEUWSuCW5Rro8IflfwvANAhOtB7xNxqt0G
OqHlDXsJO+ttLjLx+Z96aTtA+Ds/ig1LR8bWadfmTrHEvxZU5IbiPmiifR7BMx3cgxG13YpJ7pP/
NT0ZaS+pDO+w2gJ58E6EuhVuBO2OyygwcHrCbUl15vbx+bUIdTzhmmmhFFbMNS/0khmMtUA1TS9S
RJc8gMy1FsMQymUWKV3MY0cogVDXAKKuV6Qblyk3/Mt6roswzQFYrgo7wEVIa8KssyRd4B5TEHGQ
YtMRa+W2eZS2srVdyr9u+2Uq6/S920JPgEDsFUAqmPUSrUPewq4XzTNjurQoC5ms4WbwqVjB/NjL
Z81rmdkaczk7un5SPJjLoPkES2KpN6Tl3d2zbCtv+88qRPE7IJjtCWRqr+6xPtLqgVTnx3N1eqCA
UHh8RVZmqI9Iz5h8BDCTGH9nakBJazRrArxEBq16BKpLavuT1+E3Q+m4BboN4SC2aS+qCGIXUNHX
NWKokdUpnoGRrORjEpaVeCI6qicYEYuoJlv06mzwmxagjEnOYhxnucQZTUHtHEwGJ3Keb5wFHASS
1cs0BHFjGgKkPBIKS/6c35hzke4AT0V9uwLw53quLHR0brObZ8Hv+9f9bxj/t3fdWwJC128/gx86
3SIBNkNYyanZNMmq5tXXeITeeHdD0CL4rZyZB5Ma13GrETOZwx78io+SY4d9rRkPnfyGjqPEnH8y
mLtGYz0gZZiaLeCvHV1/UdJXBomyB2qlNExTDR86U0m9b4vWezSub/q1XFxmT/Ucc5JZh91+IwE8
6tFy1F5XOarfB1d/kZk0Nr15DX8PzvkHOQ+uPV3dO8M0csGpD/d5Joq0G1ZmizzW2sCGddpxCaKe
4yGVqYbejiIg6/G62vUvREFtXrgAm38WSWhIsv6hG0y2cPhmzwoqGmmIr+PSPlYI2QCUd3RgWuwp
XxX0fFwwX48P+v6extG+Nzo+em45aDm6tDeETd3s+r/4S6uGYbpnwVAVuStvjKcwOJ2RmeoSjKoS
QzEutxpngfRXyeJL0AddUsvxsD4E0C9UFWv9pqSqrarg9DvL4i4moQgFAGmhPosOBtP2nWT7sYTL
jq7OrWPXW9UO8WQ2kYN9L5OtCvEgkIQRBCIVtruO1pCfy59PISFgG9C4wE4lYlYShOYpHUyApRXD
OmcJC7SEW/8olsb0vysBf087skjOJEls7WZz8ITQ2tGbwq2CzYv4aUPQBN6yHz5xQEkP7Xpn4Pk3
jKmGTvgjo9HBMUzjcdEvdZlJyxIaakYjd583e3lsKVjePMFqxSOUp6Kuo7GOUapY+7cdOYhthqtp
3Fgim0Zi+k6dbs4UaSSQssJvtQPNFFRerdkrYrPy+2BJE5YAVFqCKZ5EydrwZB0iVFVVvp6Oovt4
ObJNPB8KATsHl4YsIKO12xcY1wL6O2ux5dFW85dkUORS+uxM0hOoiRVakCLM4SR6hIravHBBEEoX
GblQY40OlvEXpvRTULW2hzoa1QJwhOtCOHbuX9OW2te1+T5b0BvU7Tm4k9JsVvVIyGAmz52MSKje
D/Em0vjTgPlWyV2Cun8q9kr9hIGJdeFy0O2mbQpEFdalRRLBEuuowgQ3z4ex6dpwnLg/pvImojr7
vUxa3M6hVabGU6ij8d0w/aTxveQoLNng1c4TbkUPbV+Z0C8gKAY09AtEElb/gAeETFOOy+8PgqXb
quwJE1IgpKU2r6xMcy+HziEx2+qYycQEt00g0I5GT/y3p4rLL67S3V9zUuM4YbQgbGWqXVJrA1lN
vTqEX53E6hNuI4WupU9Wpl5Uu3Ji50t2rVRSNL6MkIIBSnNF0hJ4t+s4SzIk6eRDrOAZc95l3d/C
yUVCNVm9f1kYzi2yOxz+kT+KqPJe3vHvKWXV2pjSa+sO/DaFlr/+fkyi2eZwNLevkvGPTWJ3RAn6
sKb+yer9Erkg0s+M/qnwQ0xkHIF2uYydIf8BPcErk5zW0KI2QrXHOgFrIwoxEj5RakSbjwDyYZYd
Xy33EKgfk1ALfSOjBEaG88XKtzn41m7AG5NekkquEUdrSku7kD2+gQr0a1IJq9zJ2YXEdZAwE2yq
Pb3bgPYoYmsbAbrzaX4mSNRB77HIycJnhP9/zuhuoBybLlYrewNGJwcJue7+QfiWuNBUFPbm35Il
Ul0hlp6qfuk+lztBHChxLKVeTEzei5hSl1muas/5sAwaBxlVrfI8IYIWWfDbFtBATwUH0/dODr76
v4RrOgJVdK3WoG2/1riTXAt+K8H+W0QL+E5ubT9xsBz3aj1pHlMSPVGbHwLmcFUYaouxNLf/Creq
OmA49z8Vome5zgCweR0zboNkgDAQV+uIYQZEo01asJx2cUmxOjyTCQmpg6yzQps9lVmv/qOd/i2m
OJZcFgMRAxGc415vXl1Kz8rkm1mGodghQW/4gA6cdM+/duGT43I9ij+dxccWwehURq+6MaFfZBid
OmZDQF4u4lBn6E1COGseAVTjOHnrhFezi6Va+nnmCBu1KQUli01dVa3RdMvVHKrtJ4bn4wsocqYJ
C/BHbsb056jc1XwdEwEPz/Rg4auTc9OYq+zk19vMCMzEvdQpIZ7VwSrym/cs6TROdGjP4a1iQoB5
YhzP8B13PNGsWfgX/9juQgRI8mgQMI1vmF0ISxtc6o7tojYLiWouNlkiqOMYuhL7GM48rCaCbaWd
DGa/bHGaynrls27z5+R7ZkAt0QZjb+hGsVZadLYLLbykcUiSaSVoNFjhvoTqCmfEeXHQuiqDOcMS
XXaEV2DVnkIqUjw210M6RwC6CqZG/RkOQgzW8ooBqJ8NWyKlZa70qtSYF0E1wNRK/3ETMsimhFM9
dFiqNz1vznA5bwlvg7jYD9Ir2uEGqnd3rc6cV6P4uoS7/DW6VS81q9NB/fQ4XyqRdsdWfIItLSYt
XMdsS2VKLIvMJqCvtPd2uaQV3RFnzUEh922uQz1wpWaIHCQ0ygxboWYhscs4AOId0+uYRHKnjMvs
oawKaXwNPlzaFq2LHWQy6GAyGYJDyMljUMfisx/esek+mGB6O0ebmwYs6w0fZG/BM1MY7mk65tGJ
QXkc+HON7sInXDPFIzSengtAVTsCb+XVxKtPTGVTsXYwTo6fr4ZAzurzhCjSsoRLYQ4+XEhejWeq
Z5NGudvRkB1uacmxD/C3X7/quqREfAYe6LHC2hsKxu3TM4N/3tOYuK0K7zB3576OCK9bj1j/Tzso
ZUBUcCUsqL44lZneSGLfoz9s2jd9rbicEeAeZuwwG8gdtjEadkqdAW0jifWw852LI96AxVpEMfyY
cbTAg+V5QbWSzdPbMWheMr828ptiSjEkQsHOwbXKQnT+mVUKk4UZkqN8MiRL2Qf3GtT8YAYMBxz8
2JPwqooarxd1YR+ZroIhRtxp+THweUrku0Aqix4gReFXd0FRI1uU17dztGnu34wOtW6ZkFGozsar
4VFMz+/03GXvCpb/BDXMDvjR+6nXO7YuMCKFKi183idpXQ6+OTFRhwDWFqnuVz8vBXM2ZJkcdROp
mSkUKi9fevPRPHd8XcO4QSbIhApjksnx983qcimGNVHZ/YkRwBn4RwKiwa0kPvi6o7cv2juT9UKG
8yqLKjTYfUWcVS2zimUiPgZahuc9OUhagZQhQSV6kcieyjazxKMZjE6Abc5YD5hQU4NnphdJSte7
Dz9CQvc35L7655abnXvjQP7skRMpxUAyMswfcgudHs/Mx5m/tKqv4wqCPcbtf/qEqcLcbya9WIRy
NDFpari/kpBqvj8zFrMobTn9fVtl2cHp1fC5/sXehiCKxW4opXY7sEqdY9hkI5usqJcnkysNhdS3
s+TmBqXQ/nNcAo8Wh4kdR6UnUpZRyc+I60m3mVKE4GkaKW13FT4BEfCs+8PYIR403XKFOu6R9V5h
3zhlx4I3leFxAn/6J+ga3QfHrIARI6S7coXECbv2ShmaIME4Khuo4m6u+IYonZQGzfXPsNCR7ntg
ONEOZod6HCA1IWB3ift7G3lI5m+sZ93wQnhVdm++hLFA+F8eLfIkVER7+knVWb202R2BBErXraSW
X+KDLIuUqFiA1vzmZuQXZech9ErOPMnnKJnsEeboTeXJpxkEshHqVCwmITKCqLDMueCM2pxir8U8
afFzl3mWKzCxNSbVcoO862sxG0kTQTP/76CKPD6idtQ8faWyI/mYeZ0w/X+YEhICHrOX2IR38Qw+
gFe9HCDaMpf54XcAmru6ewQ9cWbumWzA/uqcyz9ArGyFoAIZEZrdaURpLkqwecK5bK0UDtc0ofZm
1U7DV6F+4ljMZJeyTElTQtYJ+4c2J8bOjc6/B3CBPrOPa4E/c/bTx1FC458/IlhxG6tOJPTbjmxb
GLWXUg6/xa46JLHpbvbI4iguBnEEipQShiwJOzmmRJ2y3JdI88p0fe8jMeB5/rTyFeeW0seePSss
DO1rklL1rpUmekFZyCzEbAMkXTYU7JbGrpg1oSAgqIqZbJOoNEnJhBRt+b9FL4byq9XFvxFawbve
Eh0iaUil4WslGegjiR71hh7ZdM+4tDiSE+3EYlHjJ0XfCf+NZUcAyEAk08gAhRVjZgLrGekCE9Bk
QQ3i21t9ihy1p3US3JahuSf4K4r94s2whg8jTjkb9PkvDRUigKKOvCics9rBNoB/HgmGsVlxDHgc
40w8mwKJsrn+WNXoxwLTTPOFWdirwz6Vm880KByZ7i0hHVaDtOWvnCgjkWPa4l9F8pKRDswfVUZP
VQvoPI+Kp/2+Ttktq66fWhQ3R5KWjoZIykbtkioFTscMp4u0HQ2OV2QShsTZeiyFijIlEISU4iEo
NIeLSsUY2w/+e8pVMKdQnYw8TwM3nYYplkqstVK4V0JcZwlqI1NWfyAxNS7qUM1fBGrdziO+x64y
XFv71dqcusKMO0S1DX/cpG3CYHwrDx3yTftkx2Z1iTPHxhPN9Kyn1NFX0Sa9b8lY7eepR4oBVIpe
Lw3GDA36YFK1o4gq0QgvLU/8EOeJHIgxNoqYwhzAQ9eZzPkoFDp29lb05oB2WagPJ3SHv59w9NcO
24h+xPDJk6WwD2kNCALMDbL7VkY+DYlYHkjQt9MkJVQMibTHbJZ5w5nXY86JNlPBzfjbxZ6guwgd
UL7dM4o+qZ6z7WrdBHg+lgu0Cn+XRME7TVpB98p5rM42N+g6ta6Hyy4JkHCbVl4YJg4ELV8AIEt2
TqoTh4R9JjpSydBREpQpkilGk9V1zkOklvN8z/6ou+7TB7R8miUbIULLrCDDP6rTFww68+B+DEGW
+rvZNK/ftbzetPC9+mwF/PfcFXOdZMwfEAMUPZUr7bG8QYs0Lq6CSZilOvpKUnQStRpFm3QNk5x+
G0O4oUcgcwoaDkBpWWUYZFuwfXsMscILA8BvlE4blBw+JPMhqij3V5rS5Nte8K/3q9o+UkJWNVM1
y+B9J87SFccuv0ohV7RdaiVMoAxE/QVAU0fXKKgq4f3i+h2h4aAk1x8ZIO/TqX6Fc6EEeQ8iCjcH
rG+yFhSnNNu/53RGMj+HzpklfunOcK4mSrkiK6BnZvzMG2z/ezsfRIMoDKshPM5E0Pq1GNJB+kdA
Pym3nFAJNPFXI4XWr3puj1zHrhEn4ViEmbnoaz0tCiIWnDskZCIlscrPCsDveDF05AYNkutcIjSU
dx6mrea/GsrvfAyDLRHJnfimcxKIGypR/i5IdEbAjUh/jJSM83ngp/cyf22QDszUp/ti1/qaTrKr
P/+RYqZboad98/HGTEm14zT4cTaJCo0jFRXPbuWuZjf+MQ2Y5ua+YpNc6cWlHLDEdapj3po/J3A0
2SPGlDU/7uEVs6NL9+OI9JDZ+Z8yHtw0zi9LFPxmCEechBW0etMfZhvQIH0rKtgwI00vTFBkzQz7
f0DyZiPdhVi95kJH3mxDGaA0gsRhkHddse4ASYMAc/8pxGwjzjbowU46woICPgOc/vntvQJjwfGV
dJZE1Jg26KSRdGEzm82l9cL7SPajU/hJiDAAkWZspTpBOxoJMPQI7GpYAqQ46VYbdOBPO73eRL+i
lyNGWPRU5jKEVS6f49KSxiGu5sG0tKpuAoh24X0qNT0qGTBOBWmj/x1uSuxoDiAcmniEPDmyvITW
UQ8TIc0rCNJsqrX/M1qdsIW744/yI8q0O+mk94aHxhrKAY/KIiB3KldjVOoi/43eGfHQ4zAUnfa3
RSxtRG5llAG7VTOuuLm98GeU8AkAUyGyHD8yVtBjS69CqjD3htOSgPF2bWnrszebs3MUK4EEDiOk
jdzT9mG3cyWN3wGCpq/62vxuFc3eBMdN/fXffySsihNGowawwl1bpt+F4ORbpvvGhHMgJFwU0mRU
mb1lwMyf2VnlABTzXpaPMUtjFUWNLNKFxNciwaV5Nh4M+LeuavGTZLUJgy8NcyeaDPG5luL6DwfW
8zA/hSZ1FMb7jL/DKrf9y1YW0RXIEyGeWezs6TqcXopa2ncTAuk2ExcSeFtC924sWG1y12/M7bKT
Zt8N42YadeYHgCMUG5aJhuP4QGe7dwI0vrfl3OJuycwGJ3tD/E//6mLgP6yKHjE2IBmtLPz2xznj
8PDxrwJLITs2WfOfM/A1QPl1IxJbRvc7oppLeot4UEStVr8R4HjyIoKAFdKgTc+ysBSQwJTKQvF2
1yL8HyCtlDNm/jUjCJwLZT+IeVd3kSTq/CMHY0cWzC9IAUQVruL1d/dqFLvKTeq4IfQZi5Vsst5k
v8tEReKFM2g252Fo51IKqm4oO02QA/LPuwpw+aHYbUiP4cnLwHott6G23CTo/s3ajwI3PXp41VXD
wO0HBiJ1wr6a7C6snJemUOJyw1FbReVu7PISyfbYAw6bl946uAB0xbSZZ26XvEoAsUew3G+H7Jql
voET0/+LolfuYwB+39istR8lUfzMlsw7SHmK5YQTlgDYORzq2kcoA+Yy4C5p3e5QOpTqrJwQK9CI
bYCRDwEhnCh6yky5djXW7S6JHQinIOM+zMxplJ3yOrET5C1IzRfYn+gOz1qvBinhtrGabC2CIfWM
c3O3Xa+k4khcJdTxVURbDECRzpu93xTuLNlk2+N6wsE63v6lNFoSkZMRVUEQSKSbFUmYqDoFau4H
3MZFORgS180VcbLoFtzsdKGeQpjhfnP0jzdV2FflL1vUG/xRW7YZAQUPijOk8Wm/GrLDQergneH6
MVd/Ct4MohNB/Km9TZfLo+tFi4xK/29qLwAXTbz01VVkyrrOZVNsvJnyeEkkdmVT1TCjOmUHf/ca
fy0Jxl1tj+FwefSOiRNlrvw++kv8IN+5fOZw6ysBcRT4ATuF4tLLjyYABFc7fe2IExmvHVws25LR
CbqtTF6oDd8/qnuESrs9+N3oActQOsZtS5MLd1iSDsBB5j7ccD70M2AdxDiqnHcPAkk0F3y5wGCu
ByClrnKgGd4Rc1OKCZJSh0LbrNKWZ/qIznw5U/0yLV+1S4d2Y6Ld3IPLIeo5vNOoHKQxBvGbZDmd
h6IwUiWylJfTDInBM+NiCuVKxhgo18ThXNPZPBzNXoTloacClCHQh/SmuKN6M8p9QWntUweVJd+B
PqfxaB2wRBvHaNHaXKMdw6Ay1B6HvyWWewdIOJEGJMoLGzKXbSNIi12CX5blGGMlX5LcIw34YV2e
UPln+iGPtYx03KHx0q968zb/9Q8f9gh6ga/kGb8UpSh9HQihlhagiWsT+yS/DF2HfMofFUUIqP28
Hep6oRsjdwP/Dpx9mrpcKWPzSWu0oQHGyYU7P0mpsWNC+H42CdpofXf/RBNsiEHWaISvtCmpRX7h
zBrfIKLQK8Qc+nPL7gt+XJUQmgU53DdnjZaaQ4ZJ1k4h/nlBDfSJfV1GLAJcjH1HIs+eDX3WIEeK
77jR8p7rFEHGuGwAa2U8/Keplk+Utefeu77yYc/ruedVwfD+lAOtvZcd++Zco3Qd5ATvGtgjDcBi
gdt2VGBFSmONVHg0CmwZnCl7T/K9meV2PlK/j+m59sThFodR9vj/3t9oziYj6+KVLTtFkXjPWsP+
kQczTz2rNTpt1GcVcUxCnCFx/n0RsfR48C+Uc+gE2j54VB1aY/hUq3DBuIm96oOo2gv9EoiVMgBm
w5Pkpyu2P1jzCNbN+Ph0pLXTnkejvy4vsDvD43i6NxX/yUWH1rYcjruZEeL5WrwCqDTy4wqXvOnn
H6rXBzDo9hTMdUQlPjaIbhgBxf3nLArz+NXp8qM/guG0OQFpHwmLuZYM41PrIyrrNSN/fijC9ucx
IImlr2MsfZ2lauPLa9rM3erfpV7LHw/Xzv/M1uyDCfUjvoW6DF+tZoIzwLSG/njtgf7oXo+MdazW
5H2KFysoOnukoPwfpkBebPOSVLjDA1oBx6hN4+8ZeP79a+w8PkbF8XwBu9EK4eJ/+OTBUdDe2bsh
xjjc68lzXxTZ7XC1Z/t/HZHucAnB/UKcK8ofmen0V+McHFdt911n9PGEnzWZ8d+QlPFFfV0ciVuk
xkfYrj7K2sJ6ehGDees/aPXcB7PrY93TmVwpRPshh4GGR1aY0XiI0ebsejXVH9SNdu1xU1UGHxb7
hzcq2M90Dt+B1eaHKNLKIebBMkluaEwWFvi8j+/eC2bZKv7aYnmEMPwXdLjIB41uZPF1MMMPhp3T
JJtcpZ5feqmlIq+jfJmZIH0+kbPP2G/4qd1bBbqb0mSc5WzQcmEvGDxwbT4Yc5xNBujNMupCRBuY
bN0JieHyCdElU59bWWK4ql4k4b4xMokEY1r7uF0HHwnaSxGxoQG8MSsx31N6pIo4vmxuKx7vJNpO
ehdcQkoBG8OQKOQwHeiGqC+WeXhO3MUxAzxVsxzzPXxTjtOqGCLN+t9E4cxmvOTJk9bQpY2LhjC9
oJoKClOZYG4JihWv70iOAmBlPdsrPbQr7+PjHePnS4OW7vxNQmCm9wJJidUBJSWBLtjR2dbjLCsL
xMjKc5KJlTUzFvBOc7zGiCBwipBrRnvyVfrcgKXsMpN1wNyDhIn+WeMRsT2Uwblfou2wnXNGh2lh
xByc9p3FsjPSHg1IQoiAacY3f1OPv35vVkKhLQrkPqbmk+0KqWb1E4h5le46RtGAG6/akoNArvSc
9ZCJs8IEtFt5zm2DWw0gSVCSeq90cXWFuux2x61PpIl9g6RhQlliFfhYvWypAhEuH/CRrKSGpTd9
V4ULOyGaUbbuLAxLOpm75ahrAS+TU0H0NPNulcfeb10NY8Md0yXtYMtiffxpXP55Phh7dvhqKJdQ
wiK3oNX3YPvIL+ty8TdhJJ6n5YYnGhGvvtCm4tvMuyeSbEqhpo49oipVx3IYeITBGsB9HiwrL6WU
GqrGIB+5+GPDPAe0HcaE4+kducmOH6wOH36t7BPT6sqDWu5uVYs+RBSlPQ3UFYHB/V9O4Y4KzVRp
N/3P4m5+4zWnpa5ynU0Em7eskMoggP3NIl9Ie5/lWwwn3VL6jO1r+Kfjx+IOcrgDyNIrVa4h1Sow
EIldldpS8HyePe2wI1wVu744QZ/Iq01mcPIW1jxT7wex1T+DSpckwjB6ntTeKdC4KqA3jeJ57PH7
KGlfo3Dg18jeyh/3cndqRe/6KNsRkcQLh1CnVQ26C9TmExkHSf8hI/YgktqBfbHDREbxILac+Up9
QIVfB99td1QI8OKlEhv0oamhVIRmor9Ecm5VinYtcn8nOJcCa9YMoyrv6fMy3ZofRPZV37oIyG43
NgRgaMLRlKs6id4TMvZ770MpYL4XXVn/2lFecGjL0N/UKuLEfaXOqKKwAm1HPiqUWhjqiVyBfsTL
zHIHaEu8zMcvNLO04/8RmRZ5bc/vWw81Ct+Fudl1FEtqKASDBdfxpLc4ZlIo4GgW3b86Q1GI5zXy
v9oq+qwgpMpq2V7Jmy+H9KPoKk/D/MF+psLKNNyPXWBByQg3XD4AfFmU9ucpgEOSA5hW6nWuvw3G
fDMRobGxJa3ZSLBdUWq2/70D7She5kKNn1HTGaCOsDYRGJKCU2Ks7OKvHkdES0wuRQafppFj43mi
ela65/IirWwjnfrOoG2BtSoPzoJu92RSB+yxZQEMXv6X0EbPl73cjUKtVzZoIMEie7IGM6cWlX24
wzRg88Bk+hTBhqyUUPGhtRBJIlbjskxcn5rZr1fEBVbe2bI6+VuVeXi0SNo5H1q0OLPdg5lwVf4T
iYGnJDkyFCbAxjKyVJZhZo00Wx1mz2+hrWGGLbdih9W1yR8rY9BCoZXOkrgYLQxaxikwgUjdtbU0
M+riZslwsU/sWE5NH+jFVr1xjRrN+sbEpHKxP0EIqZqsYsUSIKddlb8LInDdEKEkt+3bgTF5rqdW
KzKSd4uCmw8C6n+D9T77yZhnmu8y88WcPWv4TfsouMC0e76ibmr+4X6G41nn903zq8rhUfvOCsyi
KyoZCq+12xZPhgwgtmi4l14yTML7cs/jMrHUtk+fUlVKNWTkmPjMj9eXjkFy86tiSg2sj7vbpdIn
2SZahmklPY719ubfnz0c5Fq6rSR6QCrVI+VAxEWLXp0WLm5W+yq/5MPrZOZ+0PwCyGFAMhz13apc
qQ27B3d2ikTYee2xEdgMpzlETJ6wtg+/EYPwQwaOuADWftIbLB0pr/HVdb3ksJdihbFl22N4ppRM
ygxGoGiI4aItOmmgN+JKhUWqra3+gh9fl40KsLtQwMndzlRoUgQ12n3Itt3bbKpz3cba+savT603
9A0PPRQzWivhaBOU6i+tqtIcMvwg3kAsPcVA+3PD3Wuk9QaUGrboJLaN/9ttDzABMjQZndGSLJl/
F0ueHZXV8tXchTf8zIk6NBa5OCdj0wwXpSNCzg1kkIabzsLtmmkbUkM6ej6mB9IWSmiZqqkaE/5H
yvO5uMhbOupuZrmrp73HSca3IhYah+UArHEWwTM7l8Q1DNW9q3Dg5AxQRMZyAv+mw0InvmdYT/NA
vY2Bbxapg51YVZrbLG8sm+pyZJEj6rEn0ajC72v/GqBa5N7mkDO9TB1af5nRH8CvcfA1m2/Q1l0j
7JtTsNoMSAFrOM41STrvSyaUeJXhbAc7eG/3sgopTrIjRpdRr1L0+5UUKtkfNUCgEuYbhcVOqH/Q
Zs5R5ac62aOhvqN4SWq/duqEThSjhepSITHTRW7g2Z6f9PmJZu2lRDH4ZtPdOEQEwdmwoxt0FirI
H4/ZyaX0Of+3OLdKRmt34jAmAxjt6f9l0F+80mRn6Znn97fb5WKpH+IUk6fA1aFdjNO8Lih6jDCe
8YINPTm1cVCaY/0xn07s+H4DQIr69PqW+tYqzawRI+dV8oseZ7TeKgx8ONUPjv17zURGoCcDtK3T
QWFLnE/zo6hP0Yft5nA+xX+WAVTTBo4iTr29JT2gE6cPYqWJ/MzX6L8cPKEeYCt01uUE/JMXYrSz
6pORNqJEWJWt3iDI7TCLZJzX30bCQEcEHiCwVzrVIJnq8UWLH2+U/lbaHYQ4YGf2WIVp0i7Q9Qoc
QublUzGNfXd84Mf7cwt3Xd0mwRn9xajv/qMnZ85sDXOguNRoo/SutTzOyma7DimKxALZQURWrM9Q
BO5XqvrfPhzDs10wkugJ2u3kAhrCRxDP9KLlcyIqwoCVuJsyU8qPLMSHjm3yUr7s3siv7upzeVpr
F8LwiQbB9N5u8JhOwFZEKrAqlk8LjcdbvpIq25xT1dP40NtPqCeW39H0QiZBCzO+uoZZ4vLhBP36
DO0E+vgQ6ysLm8MeA+/B7qgSRbWXfujvd8QSR/+d63+WCuwII16DgvF6VAzAmRX/MPD4is7XiYIJ
+JSgq5aXJVhphUlpbU88LyuKE3R6gRG3B4JA1EaizwbrOPPfjnapQTyAg25tAYIE277sUctUo5hr
Pfnd0EbuMj4YxfVs66BWiV1F8wuH5kdNm81kupHdTxRlx+WdSjQon2mjP6/qzSfVT+7wUa5q4pMs
qM81LxpqSVHPsXbvm6mKgXa4KixEINPaRmQoEtYCnu9kWqKoLKp158EwYh2t/StVyRi+uoTFM5zk
wchWnBd8O8jybOUffoEHyV+3LbVlZ6KYI3M8vJWfclndgU4/vJfidvf84u7tJzvRVCnxWebAuv6M
dLsZRXo50LrrbobHvtLcAX+aLWXuh/Hoy0wxG9nxsUI1RpCoMnuX4L97oIbFUqh6j34kTfzc/5M9
gbuBcA4mh0ygkuXElZCNdBZRyt9yYOJS8W0Lk9LPiWD8VjtNMaaoNoux9v4NJ+zzsM8XPKbDIH3l
O6smW5G60+JTJklLAWKgRq5Yiut3KJBAxAVWW/v9Fz03ZF0Y83WEh9QuozFkxMr8MwI6T0t3YvwY
c1Ldyrw2M7/NbxM/V2Qc1Qm0QE9kniYyQ54CDi4MyI9LTzCfLPuFXnxE1FCZyh4bIvKGeM6i7S6K
lML30YVUi6OsKvn5cKtGU9LRkLmbikYjPWvLk6laUikvopnyRj3EYxMCzHLccrplzTCiZCgot+V6
/+3LC3lHT5LD8zSa5ZTxIp2k5+p3kvEpIsScUMrrR2oaWtr+t47BsZBv2xOD1DdyFpMLZy5of9G0
0O6diR1M8NFJax8unCd15/8e9732pQvgibwWchxwB0aNVWUWzDNKr/ruueJ/sz5jpXFKO7rCTPdl
wGR1sJf/mscukmse2dbzAFDV9z8J07MLF/pv4DQssDEqFFskF7LOaUKfJTyuovG7KlRnPDg1pfTW
gu+FAxI8e4SRAZix8Uzb8xBrouv2UszrG7HuInfqTQw5wF/bL+g8lmnPz1Pj6LDXNR22R/2zPcIf
fuOReavAl+MB4hW7t7NkojYMoJUhpqEnaktr/QSjMYyfOYTzjXMmxCjaLLwHao3vZ5v4ZzlVSba4
sT55MvLfei6F/ka3s5RuDA5yiZ7pvuSVb3/k5Avckslxd4qy9ykM/RbX+m90z1d2o0eZFnYaaoFk
iCYZTEDWyHPvQkXjrffcyq8rGvaWbQr4tZqHIuUldwSm0QM9v3c5eHM35U7a7oij/XK1c7T9crds
bXlJaWyuoSu0IIdPbexgmYsW4rLL+EWtBLBHnpczd1JzKLXmMrrmDtzsV3r62f1OaeCnBlcdMt+F
vviyu7+0oVXd9WTENBs65orI13D+37TvsGMeO1TQ2fnVPchr2wzHXT5/14vQvdMxe4dAxElKvvr1
ry8msye1NJjQ4vL9n2KFHZyOhWV53ITrGcyDEjWsFgmx4glD9p4/hlSSmMgNLxD4gu7APks6NYgz
JndDV9qqbQH2kZJ79iiu1CQV8jRLYtONYKWUcoC4E8M8TlKTprhSZC2y3FXVRAnbpFPtKKzx31ai
qANB8zdIMwzFA32qtAflX4rObrIqMQlAGy2Klvv9bocNjXZATNmPoMup2FaC1jEdAmLo1Z0wP8ss
9MLs+8tabWWYMQxonvS7RWwCw9NYEJasrP2UeaU5x0vJtbhY6+BLSWPvKf10ceLXyl2Nlo9j5fmP
MkzU9JffaRzUtb4TMNJ0sBKpMrk0KU0yl0uReHYkhyuFXHZX+4fT3VDtxRb2Ha4aCM+9L5V1e/v2
evg+MPE7A8VDMOz3r4h9N3FYMJJjYlK5zc+mKucMvjj2Qlu7toHvkd6WR9jUoROdQQXN233/JAW7
dHcY+Km+5ENRREpJlTC4pt8mBg1d6mfooKGDNnaVjQ2ZOjzU3S7l0uZHiHh+S8sL8o8lnqVybgxy
8uxcb8M4M6CwpK5Fz5Q8V5JHk8zjnkQ/LJLAGMEXpE+BvSM8/BVpEYXFBDxnZFfjG7eUJ8lnAvnR
OtMTQsw0p6I+FhZFo7o1dLL0VH+5mGh2ITEQ6AJ4v4XaZo2E2WNmNDWR1nsfPxzwH/cxg2lUQy1z
CiUU0E1gmRshaiOz5vmOW5MQflA8swIr7CjpLEaWFIiBywXPCw6u6aeL39u8O/7962CMe8G6usn1
VKeFLH0vTzR1aiG65q1OWy+qbR0YIaYGtiiFG5O2KNgoXDAQZ2DqMOUwvQj7vcOXoMh/mKgJNNHe
vOMG2OK0ge4KMqeGBd2lQE1YH3YN1z1tO71+kh4JxhgLG8tyiyu44OlGwCgEyhpQGpkV3wcb0IbS
oZnPfgWFhX0H84FOtLhT4NTJuhsrDwg33VmvB6zVcaJ/CE/srgeo2EwZcMjQSHr3uDmecUnF57pH
8KGUjUhct9V4dT3OL4I5DYF5LDhyhnNHhx3blLq+7CfonzOa6PSi1mD5jbyE8gWZqUUvZTN856M+
Us57Ry3KHcHo3wD01QAIyqUvj6fC0y++W7HvQvUuXo+DLP/9C144aHSGfvc3ROM/+xprkohmbPaW
K0lr0GlKO62KDjczewlwKj/yKkybdgFR7TEhzZvmjhdDEOChHw7ISSSCOim3UB1FxP8+0adgRxB+
7omnYDwHaO7N2AgYvhB5XWPCIWxyxAQmubRwL12OfrvXIv5j5LOZnbrTkfuZFVl7C3DD8WjD4APJ
RUXcwT51N0lI0c9Jf5MMUQ/92Oj1EpBbopcaRhyo1/m4812v7tQKVfwAKDErqRnrco91ZOwsW7zy
de3yhr6W4AQpojcNPhQTWccp6kyjceLpVl6XSQjwXPc46/1JZwZc2P0l6Q3EXYDidmfYDKKI5WBP
LgeQsoTNoXvnkEhNW4pDTRYR/EG/fAKJNed2bLUI+YWm47KKy5dt9OQ/+C9aVZhU8eytzbI2oxnM
kUc6nKzvR+1kbuaBJxknaSjeWf93R4zlAkNdX6x6hyeTGGx9tklR26InPKKvwPdnVkMxvasmRYQF
+Agm4NEeuYi7Isqel66o8QG5GfnyVh7r1oLhkWncJxh5W1T+EXsJW4DlK4pWjobo+b8h5V4qbHbO
Wi75ik6ysBlGMiqnCjrMr5XsikfjWDZUlh1/6mp6jfF29PK54cUbqP3K8JV+8zoxwX5vPhri1RfF
XJ4vPB/4oslSyzD69eOjI4+pgmOl683ecSgV1l5YHnuupypMdEAMjHkNshk5QO/Sgwq+aQQ6zRdB
RTymzzq5Mz41LZPLifAsoU4UUwBztGlrseWiFXey9pmFAOYwYRUz39PgAg+LXeL4+U7Q7LjbS0e4
FdjdQaMckeDYYKUaqs1wIr2MmSxCSNqluCt8ud+uOGoR3xEJVpyyv9uZ8Bj/WEWhd+HiER9P/rpa
alBW7HVbf4XnMC8TTAwIdq825iDtPFtPP6fblaiCjBaEtOfvdGnsxTQUtvKg4p3P5J0ESWvwEnIs
0TWxzXol1TI60PJSpY2cB9s6w2TFBdBFG1e2Gr/SmiR7JIREVh2JXz+VnN0eNrM8LpEh2p2VioAX
wEcCniiWxJnLPf2JM8BKRkpQL8Jpm3PhDHt/M/X7sc+GC0HVsWtaM7LAvIq/KyLtsQH2ywLkRDvv
w+bhqe2FlIwfJWDR1klzOYy5RBzHDzgSuoET1SytXBmI4ZK72RzmxwEyXMa4m1dZafn14kqdnaCR
zlmNOjJcik0mI8CIfxLID9zaWAMdBTloBdfyrjLC0D5y0BGJ/BleLoLdwHP+VMDBxSul6/loWoRE
WuW77BAIAuxuSCuBksSxHSIUABrhN1WpwQ1OG0SjHugBAVOx/FDGKCRhkqUjPPB9rylDgm22lP3o
gQRC1TjQRfZaahjhXYsoFZ6XJmWmJiEBlwSBil1Ne+aDvZyzxjehd7GUZDTnTMB4noxpJhNzo7GS
TKzKssDPQSlEauivA+rp6ySzyV5nKwZOUONoiDyYN0Zq1YUUqSRWyomt4xi9gq1O7rFhz8/wBkfh
9GNvSjLmxsnX4Ua58yg+Oj+J1o1ielpRk2uLb/Uc40qQlhG5X0WgsdQy9+OXGXD4rLbW9P9FTEFu
Rf1u077Ba2SSjJ22j1rqH8tH+ue98Oni2YVQenQc48kQ98VwpJaSu2naA7SkJLdkFxAlgISljSrb
NE3sobleNol2JCZWd0KDAnT6wbSlBQyNwRRbimy1j8IvqgaddqM7seZrGBJXJvHwIqZkEi9Q0Bh2
ESV/FRTaUg/kzaHCSKwZzvzH5A+uOPqSzN9qC35t+h3ZwgbkNjG2mGowCdx7RvV2/XSDqhuFdRVs
ewpTVW+Aw9cWl2bych8Zcs2WCbiIflG0Lfj0yhpoMcHKhwr+5sm2pOiliRfrrNhwKRIAYyamksk1
Dvvm5DVFg3FP8DNN8U9K3xYKZg4v9+wkwsPxdQu6rtys1/UEmNbLDVrxTP+uVtrcF6a3aGENatZL
gxUYj/XpmC/AVYEgmrOzd7SxUXJf/Nucj+XJtQf8iEKmIXDDegdCrfRUOxFh+gfKmX7EmFSmLVJC
bMK4wA5wa8su5QfkwBNxolPSLaaLHiJFBpX69VjBkspkGyDsUnBXJoT5RovOMSzX56KybPcfHD5l
zOewqj0laQk9FtJ31HOmsWHjRb7k+1HEBlwpPaBT9+f/qabVT0ksTM/iAj28lUVBGsxgwQaVX5YN
ml6HchxtD1yapyKv3IYgLNQibCzsekaiAdp2r3e6FlqO1aS4XIlCGNxYaByEsA4suraqIrL7fo/1
QUxKVN76ftHDJ/ZR1GAeJ6fuh53ty5JpAR2/iC957m3MVBdiDDStBU2GEvSAeXNgHw547soXDLvk
8E19DdasbFKxtqp0hPxe1cAWUWinY838lTJ4dnA6/y8uQVCUUyaUruPM1eESGNkfh7uKGyEuihdZ
Hmx88E2yqFmssru3VMrcOgsHm/9fqHqhJHJzxJgQYXho1g4Ywr0Wk9sD6pUX9IeYxykyn8bcuGN5
4NXm4Whrg0r0xzU3K/rUbgocINgwyLx/IZUJ/GWJZ2CwXaQT+lc7p8fR/JdfLSm1/jbFOibnOno8
+LkTlyXlMeiuBtqIXbbXgpwWwZO9okNzO1Db+sacpPLSq0ODPImUHEZ7ASgmBILDdEud0OvogNiA
JaPMQc8fIpwXUY5ZLuZAyp7/srOgb+eGxKdF3B5NHjcObU7NK7eHXAzLwf8DjHwIOOedcaYWEAIi
tutu9eJ3mUxsUZm0yElrKc9bKv7RVpwcam9R6G2eHGLiQBINGPB2r6cM9s2Pj+ekYWT9zHR+zcNO
2yZLPXv99vmarGsvLG+9Pvf/U+O8R4+WWlGXfpWnqql6xbfKk7tyKO1FaEvijFuuejRhYico28Nr
qG28yIwke/3lNajIV9swcR1iFo8mevnzFnkTlDQGCuQI1J8oJwvDobZsu/SsdUaApgnvYgj8dAXJ
mRpXx/aPv6zDx0aDkt1tlivAq9WYi9Kz2b4oRaC4sBGIiHYKJwbpT7Nc7W0lmYxf9UDiS21RlTC2
0V2rxy2xe2K+wGIVhmvUR4xFVAfcYWBflN7v3ODL2DljhYFwdSGnQMXaGFNH4w5Jc8swee6/S6NW
XAFugeXMmRxTqMfzJ4xsCXcImTzRD+Hofn0+2r17iMCAsSpESnbn7YDAhukA7hFWo5irGCJdzrtB
yM+vApiT8dKc0FMjrD33xf6hNPkxXpmZNwoj2AaW3BMuXqKhcGUVHnQvGh+p5VJyTKFIsUwBzyOw
mTL5X7IagVTkii6dnWh87+32SrIkLBXiNYxdWEhH5G/E8TXWBcB3+Y8YDhUNAWBj7OIdHPxisV5E
vqMt1epdO44f0I5tVMOdd9sKotX8I1Ifp7QoNptpqWUCU1SIzzgp0cfW52zwDbMjEP8i1Lgawxbm
b1DAeAE0q3B8hPXWAJNBtEKEi8icOHITC9bWM6fL7rPiguOgzYjVjr33dpcz4iRrEE81d0FTtsSh
2n/p+Z0yB9xVm7Y4cr9/Ld0OFhtfglTmtiGrW+PGlYbUzxRGT9QZwbI5D3kOj8QuN0zU8ZpYk1+F
T1IXD0UlmT0Bpn7ugTvfY3X9IsEYYgvVS/x5XFbWbaOyiSrl3bKaaol6tNsYKeXE25BygkYfSzL0
7UZorkN00/+H2PxTo2v08ig7D2iSvN/vdCcH+MYQUtQ4s/h2rQHo7bsbm0S814ohwR1Zlcvsy61V
nY+JTz1QRKB07j5JDnjFzWnAYZIvQ/lbr1YskrFMkDm9VdlqJe0QAgwTQJGqXyIIt9DA3ChRIsRz
lHg1kijsDl2B3uVw7RMC3vyYffXnOjQszcuGX4jC1iK9mn8KtlzGAlz+U1SWB1njHw6vB/hM1iW5
fu75cniaDDGHmYjZdbH587BgNe9MK0P+e5r94EcpKgq9bUKrgpHS13zMnKCArem2iFbpeOO1uZ2/
CO9XsGqQJVmkJFO4TDGAfVnryWKVxu0NUnXC7/fKa2Z4FQoB90m1oelPhVlBUnVHpgruJy0I8916
8Vu5/gQlc7HuXSvLsjkpKoWzVjgyXpr+O1WoVnEae8E2NNE2cGJ2DldEicP0ZecGeJzwYWRaOAqp
MODke13yPL03UkHvj673veeBwewmpWwb6u/YVTZhLtgQP0Gvz1HVna8c6TxAl8U3mnCC+utkqZJc
01CAL2nRF6oiuuDBFXj3qYoJ2qXTbPVQOGwrawEqCZpm5crLfwD4emrTZz6qlxWteQ/TptO/5FVH
nkLLYty4BCXy88x90Zl54wdrNJN7a6Gy8iklUy6qet8PhQ3chANEIKMCMal8wG1SePkeBKvq0IO+
cRYcKDCfi++GQO5Z2WDyFQSyhzmzA/t4Yfjq18NxpVgHeAkRkP/THDKGbxv84nqnm5lctWwTdJYg
GNYmVdtFPXckmBT8/YwufPzS5jkIRE45+kzOcvrk7a4OTRVi8/DUJQE+PqBe8VfrIQxWjGLmCrPC
6Xz0inLpisBwcQqqN0ZIR+POaK8Lya6woedxw6uA5ipJn7ZuvHVm9qOYTd1kAX0ty/0arxkA/2R+
p/zySHaC7CTd7wci29meYQKrotUyADVjC7AoFnTlxuuMV5PYRTYOobVIhGhuB7qPTHTc2VwpR4+m
C/NN/Uk5Ro/9RTOhvJMhHJcMfX+1XvyXmC36tgpnYYQsE9mMkPa/qTVequRUnR3iNkWNHJuocLSf
uxniaO8ML6nySjdc4qOSG2OZS/TzQz6+x4hsUCcNcSnwZYbTV2Eg/FXRdAZAFKkDzd3ffP6YrmkB
qcFHxSKI9BkT5sdgKra75kc6eS8yUHazwbWV3kJU5uyOZpCmR5RFYF17oBREZs58CB8spcrMvMxS
R/Fvwyhz5HzdGQSnZ7Ren8fEOGSRyLtbgDGTxHJTJSvJl9wofdpVkVv9EpiHpwnPUbm0n7X60TyV
YYMGJkkUlUlz5Q+yS9HJIBg9fFJuVLTPF9kPolphzFOjSJ+wXnA6yM87vw+evyRAL5mVdzmCSOtp
MgcyNqpNC7AZIN/H88QiZEc/2eM7yZfZdeqMC1R4ie7J9TD7NiBUAl6SF67Pzjo7I0AhqUs25dit
UOy+EebSCMpuFepPJQyRPiyZ1G474ytRYtNq36q38vUuQsvhf9+ZyXcY/sD8cebfn9EWcBeD10m4
5Ixt0ULwoQSD7Ydzu7tRyfPBmeOz2mWm0Gx0CVbZo8gIoW3g6AzdEIxgvP66pZ4euW2g/okZIuFI
Uo3Kxp+Ebw1J732deQdPSxNbdvyijqUe1LuNZaIjiEhWUoMsaKabDWNyHuj5U4WV9KPfG5Xrtx96
0Int8ffesxQNqrwY9te2/+v1d15wJqvlbVlJ67Hq5yYGG0V+n3YQwdDPoa68SmJcHAlyIKuegew7
NvJwLqZCZ2CPNTtz6Izvb2OsUM42p9vnIZSkde67aFlj/nqHs+vdwGUuYGQG4GDzePVuIb3Pakrp
Rlz9eGh24XkpjsG3kxFrnnv+UvemDwZEJ33du/DKfzvs3tqzZjIPeAj5HnoEDTmmE5+hAXAjxyIL
7T2emOwtmrZxPaFdHBh23N2/jK3dFqmMayGDWN26vYWKkPGsn7oezDA6S4Q7eeOXF4kqoVq0pXfL
QU5Adusq3EwM6YDDksnvR1rlWI1dNCKbwqPj3SV4H86c3699TNUnf8GkNir92ZtUq/f6GF9lMEh/
Ns+KdE+Ebgc5aV0e6pPq2MA4CBw56BUg+uQTdideYyNtodlX88dR7TFLywa+KaLL87KyNW/fWBeu
uVW2WD+qkdkhZja6FPWnLtJ43grkC05/NOlr1QEFny2Rm+tn/SmJ06yJs1uBXHG8wevaLaK4iUIa
YCYrq2FWeCo7rp1l2zYwr//4djIkj3z1XXYLI80To5D7oK31waRAbBSERwwvIwxgm08z/RP3FGNa
iwe5J8ekwxbk/34pI3mSa+3ahwakGUiR6h4X3FMhPQd85ygRi9OkiAfoTIgb7nowH3pK9SeuaqXu
S1fcKZxzP3P5DKuCAkuYGIhRNpGKTGFLLD7GjgB7KpxqyAxHZQymAe/ABjDeN9UCfdBydI+dF4BN
cQ9XwwTZJ99EyjfH5BtwEzTokPIFsDCJb/krnqGE/TatH7NlxJOFuMvd6GQkzAWPippMXYAq9BeS
3GIedrMPE5fXwmi6WRlg/GjlZcnE/dyzpfkbT4O1GPYQvTWBBCmyTOVoS5ZkNa9HD/fosyoPUAJC
Cr/rDukFIVfBqNM27TpuptGQK4czsUHoG6eQMZPKp32H0Qg81AAobGUM13v3MkF1ngT+gwFq0RJw
7NkTR2ZjHPZ1FrH4dLr0dG3Z5jxxwwIvro5WB7ef1Ji97E/V99FDXj6hr8SH44fIcW3k3DTH+X6g
I/Y4fSrO+Kj6whXVwGGGodcYCFru3DK9K/iUnQHmaUqDDNqfysil7gdtEbBWYpx5b3RVAZbelzD1
tpE76BDnrjqnICXwCZf8U5/quj3ZULUlgI2LgKkN+dYOgWqSAGx+LTDMAhxWxBEIdnb6dKIp0rfN
Gp2NNgjA8d3GaWvieC951qLblT+AN9cAALL0Dzd0oxILqoiVc99kKy/elOBUWvMnUeJ3ERKA7X7l
eDxkKpgYUyw12shfsJH0idqmCtxTFIY5gsccwmSotyHb4Wj70WOPlbtwIZ7WdVoaWSC4DrwL5oNt
EWP0CkurqFlLvmnDHSy8XBvHnuwBXgQyJZMKWg0udB/RyepMA3538oS7YgptVpWbFD+huNXKMEcx
zFxYLZGQTKfRGFGBeTmLcf1CyQYsD2RPA1swqBjafv5aKb5rUgsEfr8NIMvHysrFY4JDrQ/W8Unj
7tjD2xUOoP6ICSKNHhGtideO5uv1A6SeQB3xG0xKvTPwxq8JHHxL9yn57kXla3ZPn/Qqe1xBLM9m
uKq4VB2y4EHIxTKmOviz40kjkh7hVI0OlJuuWP9UR3g0JqcHGLPcqLB9q2kF8k/ZYFFibXn+Q23a
A+EbN/zi/9RYUwKVzEQcb/uWA1cEzEy9BcS+lonqWm2JoLaqMFG5Gt0q2jIei7yPkmsg/q9bTBRI
urqN8veC4+rxqOxQVhVReA1iETDAq+CiSA8NOmupFOzah9sAXLaqb73BUdS7G93wtCEChvkTWNdI
Z3jYUcRoA4h82eygCD3Ysj76zQiZtaOYDSv+tMcYIyOBmeGb3FLJtA4Mvncw6BcPFL6qrCHC1+LP
70z9qV+2HFxFf5zFsbrZNAHxTX7/JeyjMyPykA8txhqkiujeBErUsGPBJbKEhofdTCMw8k3pWuem
HhKlirNjFpirA13ce9mUWa+E/zncj/VRkdNMDH1/WgPmZdr3bsGeXTi4cxTRHgbLMgqa7ssdUPkF
d3Rn6nssSysfJoB6FN403gKDNL38/8Beic5CviEF2gvDxQOvK5cdEgZy3CiD+fts0oMeMeBGagRh
CLrg27PP7lXCZ1QSEhGy1oQQm1s5i3Aa6RU+Ij9xmutxjd0gxUVBuBt4Xn/doKfe9PnqmD703KLd
8aoxBRnSIQlf2iOsTAjTEHscUGAtNtSUeO59g6bHxyJ5/oK3qSCujELK6Q66ZW0BQIpQmpLV6Kzr
HAjH4fTGkoRMjK58IVa2EJlG5F8WLu7LevKOLoO3CMN8xdOWVYZ1GkwLalIDH1XRjxGMwqkxJGF5
mszsR/weAh1Fgr6Av8vfw+2p5/2FuXhvNgq8Pu4A5ijrap6JB9xHbSNk6N9tqJXM4CSRoHZ9qJX6
B+HYYoe4HabFImDkg6Yc0UX0C5In6YK8LPyE1+lHNEN9/sq41idrJh/s1JQewGGQG+sy09moZeNI
42B3AYOVrtmc1frUFcbEKyAbbj2fxtamzs8rk/jcYZljtb41Fzp8u4keucXWRWWsnKH8fOSbWPYX
lT6AoEDI7utLpPAPpixo8mByxVd+9Kz2qmo2240S83yy5mFte3w4JsQp42EuxQGziV/ZCT8C8UCw
YbkN7lUjJGWIl+Dy3TVttYsBRPYgLZ4GE0y34kcZKDys3vsVoCiOfas7jK9TyZX6H+G4gFTyssKT
0X/Q3VKJhNumPERIoj7OqX05kyKgmvvoae9QfncvvdNWZzTA+WFXY+kGjApGiljxfNYeZjAv9Wk3
pr7YwbJXJJNBmORti9hRWgdk5jVqtipE84VitCcCYjavZrXPyPCQnR5D0wVXv3AyZCY7QIoD4FYc
H8amdpKmPn2ErRCxrQvJ+FgOgBmXG9vh874iEIkIzx9etbN8vIj7z1yHJyU5MHzjmY5Ttwxa4F3q
G2rPDhYDFg+AoKt0V9chr9H8+LByadkBWe1b5UhLLj8C5LqjdmcoFE3ED0UMTlJJoBwmOMwJbjsP
L6WY8SEcFSNCZuQYxCLseVtVRrRiYF9LaZouCnWQzFC1wrT5vETT/HGCYZjqqkZ/0HTFO8Fdkmt7
JVdKQuxD5vh0DGLOqDe6IvRS+ymwGYedq252eAjJqSFK91e3EE3mWyIVK+8AD/Kt+cfCkj59QRl3
i28QNacByNqOBqZ2vURsWGMzZx+c89TBPdqdlzlbTieCnBlhBbVXVZVBsbk6f9Jf0IhLhjwtb8xH
Yx5J4HGzOoozuJJcF1q1OM8m2RTzepx+TEeZy8ghGnd8+xol0LljAqYpLXb/ujB+8te40xGsdtBd
aSYTioqq2UipZbMdK84+5y/hXJUClG1/Dk0eQh74ki9rxflwcicnpPWPVlEUJ821S/hbp1lFk7vs
UxENP3tRYbbwHkQ5JO1deIMYv9YRTZLwTQ4eu07sDZCmhBqeDZg+ieYoLvnRtCXT1hWSKXCc8LkI
X84lGPlhNiesRF1qL9Eg1hWeUBsiUHyMY1+gNe0EljNRdLSelDTwBnoqAoum9Z91xGJv4nLSTEUc
XtjocwNv5+vx6LC+SIojbOdJqdjEyj8tivXz3aD5BAH4Wp8NNMNQeVTBOX08TRRuRHgQx270myAB
1zNJB6TtpQ8dTLSl+CWI1CFAK0z7qam1uHP+j52+drNHrTy7UQLXZFXAML0d7AzEv14G5mhUqBN1
cnZElVJy17XyemJ3IpLIgxB5pem5Ot/grOzdkjOZPQiONYjG+ucp+l1Xhf5NPgxaelrPTON2ggdS
HZSfIG3dS4UwQURFpeq9TOkojDUjsYoORWz/+DoOyOZDKaeWetOOJ2pIQLhoA41dSGOa5czvJdPv
3h0EbTVB37c4k47jwkzKd7cYlmvBJYWhwz97jY/6mCKzZYEqWAc3RT3fc65BjiQvWstICHYvLu4v
pVmZNSLr9muNrYKzop7ITn7A3SRn/vNdD5untX8HGUeA9LcYgZf2m550zQHw5vKdRtbKajigRuVM
5x7h8EAsokgWld5FJrgNeArHXncWxNvJToFI8TV8aPF+SUKjPq5+7mUGASquCqHQ/dQ8o4etzW/Y
OvmL9jO2tdISaOPUiQTwSA1ykfvvwvs+ksBc1WuRSDV0C2IsiwKFHZ/uehTgh9XxueTOvLCBsIMa
IY8imdG9+xX8Z8vEmeAIXwrMbPWdaRQgmkfA6JVxyJ2uTuzPKnHZEDgJSryiyqJS+umbhPgveSw4
o+oszBwKEqVeusQVvH74BtEBVCmRkidS/0yblIE7a3dFZiUSwmGq1V/I/5jB4ESS2cbSuZbnBrgk
tL9hj+Gh1DscYi9DhcEpua+kRTRiPBz50WJHrrwdJkbODh79vcs/VpUdW0ih2aiq6rtAKCLpcn5y
fLmX+axc42dDDmj6SNoBjyvhQLOiUzHq0yjhG/KF5K3ATWVsxpNXODc+kcmPv/8J8D/ZdboQcJpX
7YrB766q0wAKMG8OcpyhQ2qLoe4yRwKKDsdhRpG5M26zz63uKtS1zi+Bmyr8XvlMK4+7ltpBDgPN
RCU39NkR3eIKaWgYCndtipgaiRV6SjyPc/3uFKpVHqsGvXOw23IOsDUGLFwlI6gX1IGTYHZ+uJjD
Cy3Z1DQRvfERiKHwzYWlmBcYO43QqB3lbFTme12D1Z+mvRxdoApbepAWBPbaMAvoH5oKrxvaJ86p
iY1MOOCDZbe1pCg/p9e7oq1p0rZTGrfPHymJbTZyaAddJOHFRFDT+yexZrIJoyTjwgtcFbzSX5DS
Hs/adGXf5CjiwEyb9YRnG2Fqap2/M4ZPFvHOlOYEhdLYKKvBqFbz/pHUUsti40Jjd1wYoc2+zL1o
4HPy7KWV7GLvTlazMWcsEgNS+Sf2Wbk7tuaNPPiEVxIfhDVLYBRyuwVPgs/2nU8dmknhZ+50+v0D
B9x2B6aeQec5v5GyoncLgVIswGt/xzSPQ5GJdB2+Q7GfoXRPJFYCnENVbWNs3zYZb9v6I8nhlcF2
tF4hjUnlPD6OL5r5KONNdrPcnbS0c6g2L/UG8DUK5aBkzAK4+2FEOXCBueuBnZy7glrCboUKAsVW
+2QaIAOr3q/MQcQKTQJiIBvEn1JC921chq3knPc/IFHQgkTdi+vTkTmDk/x15huk9Wu9GNFnz2KR
2nFHg2hTElongjIUSA29vLdE9xA3gtqNlpMf+fKVlNNN7Ohf8onXAX87/LSnY+/66cy2KpDA1M07
mEO4DZY71UGBJgYI8zKxmWOknv9X/A8CqL7ANizIGzVWOjDou5BKOl5hRtw+Fib+BenxNRPbuXij
R/Vi0doiwKY/sRqCVH2rMOrNl6qtrJ32qQZNjD6XQdCbo7c2klCqyChdVMxO1WiKAJwINID6tO79
zJhzIYMEeGzQoJZOkmJ0Qhfeqax14dLS+Nru/wCIQBX+LB2ROTZPKvApJIQPzVl/G5LVQxO+Zncg
oX0xbJpCZP9QiApVkPnZS38w81qxSyabNTqyQXcEz7VcTf4jmiTye4ATJZVb3C+epQhEX9ebJMIk
CCWI6ZdoPS30zeB6FhnvBexfhGT1kW+LVf+EuqYR2qne7s6j5Z8ih0mbDH4iddkHkEKrQpoD1q47
2Gqjl3DY8iS0vcYTnecfvhxi5J/Z9UttNukKde6dLBvWCJBzMq4de9/32fBBMctT2qHUSZBG4uwi
WDNkXrud96v7iy38zYn+0mtRVVjTakK25gMCvSYo0LcOny4P46dBcnWa0dNIf2cBOK2mwScjgyvz
FJLTDQdYDbu39nRSkYsgJVLl3vXlyXyZzrpmUztrOYmgEyNMv9WO97hCWI2Q60N7kpOuvIe6mxX0
oTE4bkWuNmyRVKzQt+0vZwMZX96U7LSR2n3HbJTK5gRjNIqV5b3DyDNUdtKqnlqOQTZ+pDEm1ubD
NDpMIs3fJM3jaUg9b+4WegZZHkZfqkh8UC83oPXxpvouNsUeHEt152UdbhdNK7DK5fTxK447a6O2
8s7BtIIAAWP1h9yms5pgbfIF03cmt0c9bgatt/1sk6dVvRvfbzJ6cUiaoPk4iMrtNSmK+RLjYm05
ner1Il/B5IYqeKmeOtMHIFssUtX3GlbJ7Z2esOALpLWcIbm3BGLv/p4iDTHthDLGezl+7zyUw15e
8v5kiIU1LvlpYvwTSpQT/qi9D/To8ELtK88n96QjgnVc/vuwTJb6J7aL0+m88XMl+V7cueHwANb+
F8USZgVbfoXFovKPAUZWA8O/TIpCgIr34gj77MfUHuYvL/iHQsYomluv742gMyMoTTRKOkHJfkCE
H/KciL4dESMCS4S8gkDlfZPXwher6hgJcTGTejmJ+W+sPJcEjGyYBHM0DvVaGCahr0m0CrevGjBA
wFjEPKrTFIGQWmUFG6psIrSeIqO85HSmyOdm180DSVMWaKDP9CBmiGbzF4Qr1VSLC+6DYwIJiv8Y
WwZG/nYK25i/DYeq8b6XPfaFAIpx++TcsF8PwXyR9X/Vu7wWzMBhj08LbeWA57+Kpt0FFPEH+sWW
vjTOC4d6EWj1cayo+etydTmQukwLppZ7NZiNv//O0YPZNV2sJkPGySpSWLHyq4x5E9Xp8/TTWw4l
WhTcNke+zlt7DIwlASq2Htk37XZjDZq7ww8ef3j3S2VPnRUPw8o2ZpMbfiYtR7lye01TCG8f30O0
ECZ4wlkuvcSuuFFSIB8J9kMG3jR7/qs4YKEmKnlundY4eqTu/s3sJm2axC3rYSxONxwKfnMFQNuu
hVEmgnhXIum5jjshBRShpGgL15SBTZtWDrP/5r1c08zaIiNe1QZheZmKFRxXcn2ep5T4SoH0hVR5
OThmfCRUhHZsfcSA4xHffvZvpQXWrC5gR33yMvaIDrD85eQpm8wKCU4QMiWRVJfjl47PH8SDQkOf
3nj8LlaONmC6rv4hwhksnMHuCpyruTNU7q5br/HT+gzK1r+QvTrxuJ4eOa4KbkSTwbCqb+Ny0Rgm
UeCX+9zRfGwqmtqp/po8lpi/FGbc8WuhMO5uAg5WDsn5M4qwXM7UKMA10GJAY07PADZXeI7SSK8F
QhYg1GeWjZV7Whq2pBKvQDnLBZZtXvOF2xFS7F3mi5u/62tHHBP56eAUJwIWiVSnxh0gsVZB2g89
4apx5yw2Ng6RJqGCLINd7O011NIgh69yLK30Mf2loEMrbEdcMoFly2ePLaa54uDFZotECMa+3kcb
rvMG1HtRKIjhBWmqrmUy8SjZfKhcYDMw5SVHXAfFCxM7lhQBGLJSco1lujjCy4uXN3hpE1aPgtkq
QinlIwV+dOX7EiOrj8i7Y/KxM15lG7S2uLTXiaV6Y6/SaH1HxgDz2jVfOvdp2MOnfGpZH1xHaJEd
Pj77rgqXKO8E+tLZ0DLPk4HF0qN++nhehsSjH1ysnaXz63qJ1LSoKN4uTLaQP1OHDTf5auDZNT9d
VUaIkCcZq+3cJbTxWi5f5OSOOejna5EstoBnQSEUx4x6i9rz0iGmkvTOSfVGMiIuLhTqsfAzBfax
hp02TNxsOB0pnLOshLYaNu93M+UPQHSOA2v2v3lV28EKl3I/jEwbN0jm2raHreNx36dMkmt88tl1
q037QOyfz/KzQYzBJfA8HH9IJisVFYeaGaQsbteyh9DTC0MI3Rm/Sj4STYtCNz4fu4C0ZR3vfwr1
ar7JEsIV/R3tq2qb3Bvlq/9xwYHpR70yMgBMl1J//KRCTsfa9RNXwFT2XPICxVS27WMgAN7gvdef
KfjSe/895s7aonZHCQJcaE7N35cMjWTBUsw/9zH3kbmeSgRG6fbI8ofnH8Nskj3X4k+r0s7PhV3W
J+MNdxhx9VqJnQJvOPAT82MasvgcdxipnixBih//G7vSVIT6AtCtaGMBy/TX7SWG/xA8esupkiOf
g8V8ryu+DHKmK7z0jagtXL1WnhDy/jLQ3acM9aec5KlB/0NcIk8u/ISpPb00i36xHoU7LZ0N5lrm
PMUiy10g3QXvngKpyVHeC2Vk/6nze8cykkcU4cCdkBqaj7YOz5ggSWOuu1tkGQu7H0TC2aCGopBc
yKt/Ayy98Uo2HtLAv4w3KobheEHAxvXQFtSShEcUAOvpNEMdaUpmA0iQvO7fS+TBoBm5tp+hA5IB
9YibKAUvzsrVe9L/XWe6ZWDOO0TqjbrkKGIfmI7bQ4SYitIwaUz0WMjw5upnlTcQRXppARjlxRuY
eF5ZhFV4eomOWEQypFhfzkILvBSnAU4B0aYqWmboNoPRw8PpQihHEps0ZaE8T4XFHEZjDVzqandf
Z+SffpGeeGZHiv//lpqnnN8HAyqHHmmpUFz+5mtJ8JM+xK9mM6k9kb+4NJkhKtAPDqTo4LXy+1FJ
uNnH7oY8hLo1wXl9ZHhDNI4ubwMN0XVj74KtQBfekVOsKtkxLVgjev2/CXWz/2gOT8+qY+VHdc8r
BL0tMxspaJ0DCdsRWdPY/RnPmOkGw1bboNe41kstBJhEqE6Ou0d5Iv8g9UbEVQWKfURMhMZE5RO4
LYtdj61IooGiOVK6qOHeUfff0hK7wwhOg+CCn13nfyRjvqN0W69vxt6ooQ2p/i7uxNGQDrafp7iY
PCKtcnLRGf9WII2JwO+Eii+VIou5+CgcRRP8mofpyeRWjQQ35YCSvCb4uzMSB7ahltJSVOOsJOy+
362uxyvn69HgzKXNLopUkRU1D3wPcUCCRZvD9r9cNrO0NmglVLXbzpIxahzVaqiraZvD6FIvcCZO
iiNCboUg9amBkwMYBvahxE73pVEFQ8za1GIx7AhORoKGnyo9+bwmtPZhyTEvgV1p5mRdiyJkwjlp
PNmcuj7HoD3uArEtBg2E5HHhwqYhSj1YoNvLPcl3xwDetKD4gkAS4LmLqJ4yNEiWkK9xAXHtNegz
IWyY0Lw6cDrQQmZpVu7KYKvj8xg7R3itlV9gKnkGnctA7GFiRwgU49deylBtx7oP8ePvxy1LRkCG
zrm0dJBE7E6nJAQZEwyqorYilIQ2XtCE8H4pZVvvG1x6pQYBzE0WlI2n3qfBecFFvZ/hq2sM6TAS
6BaE6N+uQqfTaYY5OgmtC9KH5Zs3CXnDJ+C5one0v+VxsYfxnPoEezkcNmIRQWXv6lTmdloOD2vw
5LxgvioxERgVFeo3uwEhJxaNvLLLh3VxqbytW/f2QAniRRGKrO0AMfRHoR8TXHUxWl1O9WtmQomY
a7ywn3j9wUHcGDFXk5Wr18uZMmsaLRyrCVqfz3Ae5fVndNpECeeSe/Q781nF9OrYnxRXnB113hx/
S84+yMntF7okIRRnfoy+8R2TI3j7nqfX23RcvX2fLzhRTUgmdwLs7JAxsSiDApmm/k/SvE/xPxHf
JX1dIDO+NQLqfcB2/lne3gglHkVzxHgvcvPH0oOebz0lc/u009DKN8zLprKZRrjVqm91AyoNhOl2
maA4YoJ7IMt/buFccqIsGrs7Ztc4OYI8DbRmwFKaDk2uLiwfCHLUU87dnlcttuSLxa2N/k66pPeh
Hate2soil2d41g5cjpTMvzk+dN2wgO3w0s1cp+504o0ZeYiLjF0HtkCDjIr3uLt4ozRVxbmp2DpG
zuS+1OJfoEg6qVRpje7mGlm8e0LnLzywOfWJMa4YmRPcVWN+LyoNdAOLg2FYTUp4T9eeSeEONO3+
l6ymsZfCcdCTfYFmproHZb3rm/yJPHnALCJCA7yif8niuuZXIyTjtZrOPhuww9K0f5OJ6Wl/GLfd
k7ZexvAyZM96XhBm8R6EvByRS4KaIkSYonJk2eDORBWcW4033/30nNtsjddko6+TmqBjdi09Carl
f4K7DZXXF7CCEnZEItOwmoZZrABnrgEArhC/4Qg0Ft3NgKSXs6FbbaJ4RouyJeduS2sDntwfgnPl
ht9vGGwIJRGdol/F7R5hkNK4Xxb08ELPSOexwe4nLeDyL2Badc4ts6a5pLpDpFhHcXOa/M++v7pe
buu5aMtNbLr59j70Ag2ifSd695SnsMpmqVx2EIJ0bdLRZC8Xcxvuxr3HfxnjpLFqXnFgI8hktbFa
81vAbyUtMC1w9xtobsw+J2KRbOoGFIL7Z8nKQdxMEic2weNkXg65p6ijbKJgefawE6m7tnVMCBV8
rH5DAhlP44Jqx6G596VgKKDDO3MbH+pyiAeGnpkRpK6SmQPAKmhTG8+Q72i/Pzz7uCLwj91aLI8y
Zga9eKYYxKpI+ej8OybGSrYcXFeaxbpeMcjA+A+YQm1VS5EUkJSX3nW9xiikcNRBlTLkYkuNT01q
Vuf41Tl189alLxiFhE/wCU8z7n1taq08YgtW8PsB+/Sp4lxPiEX0JSMmyr43r+sW7LgV7avdUjmz
KICfgNJN905EFHOnut66al0cMn6d+FjZ9IjJJHSZlgVxZ1/Xay8Vv3Jqdc6akw4QBpMdw2CF0SPL
vXBEZy5X0wqf6edscOf0jn6mpdvhmIZn1O1JlAtldN7pnDfVGO4KSDzdUoDqRbNdGF3O9fj5mYxA
mbwuAKLENN4zlP/7U21sKpO8v1I2+f3DUD4lczDB9ekC6hH9qSokbh2K8UmF/1kLhDDRZTu5o2nm
/l9Tic9aZ95CiqQDnlBBq3X9J23s4Mgf7ZeJ7M7vxuEh797sk43zQpQrqTIlRnPq1n7bPfDmRIUF
2rj4QkEusKWwwKHzmHUN+SP6cCEZX3m1ieHNG/RQb4YBhbojFj42eAiAxXjpK4Tgd7MJzg9bqr8d
f2yFq938Wipi93+iNUB0WP7Zvd29LUTxnYEu/YRFkTBpq8bC0GVCNmARJDatJEYxVHhGE/LBdIy8
5Y3iGXdPT/gGKDEry7y1Yms+G7Kr5fkEm7boHAezvANYDDoNDx+w0JLjc/K91qmz4KH79C8OIgLS
fY3OrlTSsnggpY3g2LnS65WZr5i2FzLtTVgcxcDx4iS1IUjic9rk9UztcyUTRDzuDePlJztINs5t
gT7+kqjD5Y8TvBk9p3jpLgZi69sFqcZB/Qj8Bi4Hau3T8gFu2DW8jB62uokN2qxuxv9E9DllpmTH
teQsSg1Aiox7FO/C6Msmta50fHSJOGk/LUEmRxTRIzcckQA4N+Iafl/4wxWk6wI3UwIJlHGkLuCt
0YTPyALZehaDQS5UmtizoWHF6bRjuU0qVNMgMX2H3JJqEB3UB5nvbZ9ne9TINADCCULD3PRpBtYk
fI0UsbftGZAcaCRyozL1CFmvcX8H8okVsubrjYhWuDKpsXTHq8r5SEs4GXWXss6ILimqFB66kGRM
2oDJYawA1Odfo4iGp2QQRomjciKQJtvzrqQwwj+HruCh5czYKCJyF7dOCFDI8Q/RHAAACmKRPGyG
Cp8tcgWMyA89c9VdmObaT33E0l0zePSuPlpKB/V1dMiTpl4C++zzr9+ofM+2uM7TAPkaE4HDLqrH
Wg67wCrPTO7ImFD7rb2mTd0o4XWlba0Xg+mn/HQzZD2BxueXXHApAK8JWJBUWIN8GtFAruEfxUug
/46m4m2rD8hc6vgnLz30bTQ3pOMYkKHK5svKM3OnTHI4SCGlOJxjJrUJb7vKlSPFCJ3m9r15AQUl
lSEnIMbRYGsMXFfPKbcA/KQ9lZAFZKiv519VTSZuOYi980NTf8UfdZX/1wPL6oLjJU4hxq1iAz/I
zfWV+yqLwyIbYlltODB2mx/AQ39MaAV5r/UVUHVw+V3WQrX/l3lZPmQUl4gdyDvk9o0Epf5T2WVI
6yqZlMMQGfsguzOlIeB0V0gB8WWIK6gwTXvHNqEI999F4yFgypsqYgoJwmCfQKaMH6237MvCyKGo
mJONMQTVi3vfGn7+uW2FGQKG0YWWxu7gkCpMQazpKOj3x/NsUsbp3SICkbHdA7rC0W1HROqsMtNR
O3Pf4x69zUnsvDMk6HvprIOqkCfMfCnqp5d7y4t6Ctnei3A1O0uKcqdQxcMa3Ixf95M+K8p9Hx5q
UnKLgf92tBCJ1ZKx5IXxTNa4Q2BZMNqjObTCMxaKIbruWRfg+4/YkoGyrkbRkUuHa40Ixpyin2I5
9MAWTVyts0+N3jE89KQKQ3WZSOF2Enc6vlbxHVQRtgMzg3zVv8hmMVXcYEOksXSTi29oAN7c8QzE
9qc5W7sOC6vvh71m9+CiWBQE+rOLuPH+mdhj8Fr7h6nSpnTnQutC6FENjmTWU7n+6WK+fUO34voa
Qh/bO+q1VZs54oLy5SF4bzzyywUkYqIdzAHxaUMbPP/kr5QbXsNM+991no2fA457LOEN65WITTOZ
RCTrOeIpl6gK0xAmpGv0nzBClZRH19Zp+72GEzlWbW8PyvkWU+4ORaNb0iVPKYbHr7TSwCQl/wFi
14aM2PN0HERn+lDBVLDxCQOBrEPRh83NnH06Fiyvin53NMtpwnq2QIJXub9RORnEi7jyR/ZDeX+r
z2suqLX/LEbx/C0RZarfDnKiFqMX12PelJ1O9LOcD1oSRtPxBK4uQmcwsCjp6JdAsl0ZzCNZr6cy
8WaOZaqrbdWiH91OJ5LIsz7SFRlSKt2GXJTYiF3zBQ0kzHS3wqSnPt2TnhPKtGGK6yHUXJh8x8z+
bYs7mjZqDDp3ZiD4v/PExj9mOcsqqGReb21zkDeY8oyCHiftZ1IHZC7gJ34mwZnqPeZEShb9qEw/
Jbf8E9PJKVhAPbaQE3kQj+2IsPfF8krCLbDI9WNhF+9c3lO2xHb4wUNZQiSp/n2E3C2dJG6hMLOr
DotSEgkL7jfgOVUtH+2CxcStD7rTpaVJcK+dBz3stz00EWQVSnANwQq47mvpumeWm52UsiVCOIP/
CybkQFCXm9SS+OhZrytE3/kMwkFn0Iqh22b4b7ItNWiCWrh+ynbbYzDhiJg0fqUleiOzd5ltMB+X
emfWkI44TtjlZ2eoJSAxzJzsVw4jnpekwCdiGb8N+JmBa7N4nE8QvLX3KLY79AbDnlmIn52hg3iz
exxLbj5p1VoyEpZTXxl2uYcWSLJBPbD8XGvdov5Bpd2yRx6AkHoiSIWScYG+kwt0foJoNhqgyTk7
wLXRZFjjRenuLEDAEt1w8cuQ092UpB9crElGG/ArMU02Oww0w8k6lxnjVKQQcwfMvJwNFLXnRJVI
q7bBm7/0An4DsnKlPadaZi6wnc8hHk7E983Fendj0iZDKeDNqocxKFZQszbuh9dVMp7yTUTR+lQ+
XqmtBvIQlSNbR19m1mcvQ5+vgo9DXRqycTxyai57Ajh0z1Ku6AwguwSTe3UGVuEzpODrrVBR5MIy
28/ejc/hF43dFzuPuI/tx+72R0qoIU1AmQXzhN9F0z1X6cxK/FNLJIYX2HuI2IGb+lNrPyZEeTP7
Oxke9tqsDPXgokrAwjNoXjbj/jjbjME8UXAwZOO8SKxDDhGF55dS7bvrXKvUS/QR6lygkxdKn+eP
Vq6V1hXZMvEldvyDEu8T/b1gZihdwo+VxysW0Z4pb+YXFVgLErJtqmgLMuKx5XxfyoqKEpcbBRQ1
hDiQKYgrJgfAhEBVj/PBJ6GW/LuNQ6Hx1dn2eU/wsaoV2zGujRlDqqGKGS+KdJdbv0LGP104nwqY
hMTRA3HVNXOIn2oPtjnEZVCyUm9CImF+NQZx6shWu6+QVPrdKsO6Has511Ws43khvSvnI7CzAxcn
+ZMnV0queBr7RDYaT58pJh0EGlB+E+hVFz95e1ukd3CQvZvRTITnA/vpmUIj5jaK6HKxyzBGtyNr
R1dk0nucbr9lZSUvWnCqtQjx65ewvtZ8EGRy2snmkwgPcL6YZ3lnLS++FsngYy5QnB9o21l5Sm66
mvj5bmm0U3/2MErYkoq5QF1o7BnUe+7q2VBdZVfJ865K0MsQBcNptBRDJpod8RhBGRfSt2kasyeI
CMSNk669XZdpB3ZiSEzYPPWswAsJUwktJSM9zHnnvdyBYLDbBO5+04Gl0UoDkLCWzkPyNqDOS594
Tlv/Ir8Xfel2KiMNR0MR2shpIxpoMG7eyAxctTsHk4jSAvpYyAWpzk+vH1rUix2cK7aTO2p0sHu3
YfA8sF0NdOlnibYzb5oE2wpLSaXulxNCBVI3aiorV90j3iq/IMQ+a0CyvrJ4nJxjJhenep35FxX7
yAvP6Work3QjN/2o+Fp0ZUK4H0RSWTcL7Et5GYfGZTqzPTgm/1bqBpKbUABgZPijAaz/KyBbcdpy
Gx8ygocD/rRlzTpV1gKkUhI4uJsUGgDvQ93A56zpc76Fb7plXs+wO2+MsmDJ3xjK2KQYqxdMFgZm
k8APcjz1aIwLDziGCSaxzpmfaGz3kL03+e0aBvr+ru4As9VJ03gO1q0dbOTlANXxQyLqYBh4XjiK
j7mJvs1IA3eb4qc6x1jM5D+2KuQO3iqnS3uS0anRJfzfK7MJklHf2IIvwxrAzubo4ZQtSnSmkWpr
GG2yWO0dXTY3/+/6lEpJkaJyM26zxBu962POIIua1FJynD38c+4zdE7nDiqzbKoSptTtkNdLZD7j
7PHYYZKtS7ivGf8b49dA3XEotxAdQVw5L19JMfgfk75Au0I1QaiZnEcx5fXNNXSispYJWRI8DDKF
0rUF3u4a3tZwNQ5o0MK8GKUC4t8Ab46SGLZGsQ+wFc+wdtaLafbJLuINBxPKAY5U4quRugAA8WZU
+7B6mp4nTPsHyS9vziBGb9jpuDnNmccONEfLANXiN6hHzFjTgjw1TjPlor7jxwK4Em07H8H9kmu9
chDmjgzkiMVO6ASCB60iqX7tQpP9uqnj+QhOdPT8WgHjcgH3Mk2RwG8qISmHwxQkXvul2/JWTzOz
NX8pwWjxK2U7zegP1AJ73O0VdC/utvvl1Aiv+IMze+3e8AUHyJ2zIpqNvg6BsH5r7CpV7ZImzQwG
a4i4twf7gtx2uaDNiJ6NrbfUvjPo4F8S0vi/6HW5oM7BGMrQg0SANl5ABXy5n2kbPyE9IUiAAaQZ
90Y5qFoWvoSHVn1CbhDXl5R45AvX/m/4IlmJmlvPv3iHkk3OjXWRR0ds0HMRIo/zcpLs54ZYUUg4
GsQbPsu5ML5mXpg22fSv4h5vrkF+7f7rH4DboCxMEjC9oqHL71Ww2OxsG+gXpgL3yYhxcUEazg3n
daQVZde8Ccm4tTUhAI+VM1oAJFDlh761b9EoG4aTYBRk1UlFduXQatmCkIK3xJEkPUtu+ug3guHh
hYsxnZikHUya7bQza1NCP84Q9eGKsJdFec3hZ6uxM8L7ZPjFuJcZnFJFFrf/uucaxafOzsfjFpLI
U0NLKbor5HZQCMxQyJq5jkW2pliyoahCio08vICZEhVLVEHCObEZOghz6T9WYYBWwFGgmYhwSbAF
dnRo9i9QXzUpWGQXVBm5apYeQWHSL+E+dyE6wjLEZuBZ5SUojbhGhxw3fNAo9BB8X4FQn3r7gc2h
y0CsJl0LFxphMWdLdWnh+XGWj0knyAAQoRv/X0tKj/iQI2mGzBIq1DLcNk72tkkhqCIql468dtML
mX+T4zf2owKxawsbHRy+hqFxrcwXNTla+GvAtAadOD+3JfFVPSbf4BgWVGVyIpIZjemumBzMdO11
y129+F/oI6YCpLnDfRF5ILDWVtKkrO2P1nc2aFYtB9y//nEg5hkUYsEinZOpSEeqt15Mh4iEiKAM
sw/vFL5t1ff6g5WjmEU5JhB/+ESSf5CRcqXq7SJyBQbN6zpcOrnVjajjHqa9IL3JrgoYyTSsgbCb
9Mj2ANQD8SNZ4YB4tS7U/lya5Gqe6s2PdnUM0ZaRtSoEOUUafLHD/dz57Q70HCDEOejjvrbTUb+i
EBu5vIHfJ+wXQW2T431DusoMqxr7ukZN1eO9lz4yE6x8KGENBUaiRSPI226/gI5IuONk9yYn0yKg
RFTqhpbvw/cWsT1JK3r8EAQ2EU6DbgQ23qWo/I1NNpYZAukOsdb19oty1DwsO+ORCRsTbkK/pI4K
v4Tq2meATvhE/AjHehxxC2cEBKZrzsjKh4N/N5mwMZ5ow4q2EtGHA0ONWVqXHUnPySgXuLYbBg09
NgpsDrP62+nlFWb+ItVhDTr6cxZyvpVJ9/WG3XNXVFGTPpaV0htT3VjNEnhT/qwsh12Q95mDnKmd
qMusZ2iIBCLRkCmUlapeowvlMXq20IkvxYDeP1Rza9ULNdEKu60F/kyESNfQXSfF5tl3XMdMgfq5
XhkAup8SG/UslX3TUJxw2GnWr8BIPR9eetZPJvS4PaE694sN4vxX7Og3t7ViwFqmll0DTiEcQjQ3
oOXQxZ368DsamlepsbqFdKSgg20pZuIFcP3Yx7a7w16NdQi7XqSkds+IcHeqjd5eirbZ9d4iJnpS
ly2PdbMsocPJxeREHhFAn7OdPP3SXTrUaBcX0qLsNTd1y78YETOk2B03MH7kzros0DgDGHJ+W/fH
Ylsi+h/Tl7qSA+1LOApUXssu8O2PKAyae1meSwjjRLp4ciPsrUDNeuPjpiVhqw78toPbfKUzQKLo
zzW81hXC5GDrresmReRcjciN2dnFswcVYaSImfhKyibZn1eU+dgyRnJ20eykDdarhpUECevFG/M6
wr6XzECzVTWByDK0VeKS6r9Xg9WrBUFFFJK/ySvTpeSz6c5Jn90JZ5M/DJv5uoPa4Ex9xyxLJAGe
wL8M8+mkGm/joPaHdOg0g21hkpkREc06rbnbybawHHD1D1rvUjj+dE8ExEOzt1mqntPx6/n4yWSc
v2uNh3wkTVkmbq2kLM45Sa4jj7BYEKjVntIJ6Gu5F2FFTLJjxLFqc6VPoD2kUeMF1UYd5dipVEF7
Vi7U2pN07ONcv5Ea5H3dMAyv8k+hsPQUpGKr637b57URNuUKpV6/J9QFFB6i2TKk1OOXs56jWyeO
+LP1o4ia2HuPv4zi1sWvHyp0piPgleRBs82EI/RB5Bs1lR8zZ4U3B6MZm4fLufATQGWW0dAZq2Ul
81g1lFAJJyOaV1zq7bAENJmfoGmpHLDMB1vFH9l7O8N+EQDNdvBurCb2ionyDhoXneEkh1QmevVs
O7UX4aavSi+pzSzRFqQZUdNK0bvJv4kt4Rps4cr8OJuJrTZUHId7tzyA9D91AaErK7hCyUpvuH+C
UInDRHKndpvfF700hOuoPWF8Ut3Qx6gjinXWQhAdRtwnQykC52tSwY9KqExyDjkMMgmNTqus2Q2t
dfwKofF/SGPI9a+mEnWH6I8+9h2j/qhIEKRciFNhB6Wn+B+hWO9b4VpwCRsFGJBrY5oLha98/N1C
OfLOdusdZOkv4pw5fIEI09bIxesiekfKySM2dT+RIZ8hHvRS0eOdQrfWk3ma24pFnIBpreUVdnsh
D5/CRVTVMD/c59HExfm9S7E6MghxAqk6977hKLafC60FlszPuODHdDws0KSRK1oa3LhqpCMBrnEP
REsE8TSEYZG+cMElaXL04RkN+tz+svGaxwlpgYmcjiseqjB7I4oQNwZndWM5NNbLyu63f9FiBcRO
Sd0Pq3RkU9ZqqO1JybyRVPrjDQ84f6nyFT8KK5xgH2u0lqMaBNMmvNjOk5wd6g0PZaDYs8KrLmDE
w4PPhC/vi6pnFQlU9jfJ+HeGaXdkAjjuVPRf4nq6XwyPxQ7JbttjvQe31aAkGA1k3m3EOq+WaslN
i9q+JtnCZwxVwtRr08u81qiNN34cQKSlWRIU15E/qsYo0HadKC6NtU+Y/fi+/uivCs569ELgPDlY
pIIlFDFlhTkGgT+zB92N706z37+N36e9v/6qKgzhGZAEyg8ii8zX+bd5qB3q8rC6IqK4WZXAH99h
VRafQM+Z8ot8YpWl3KW9Y1zzmEyFX49HS463BZlk8NaTOMcFtoGGpFbgTYYUp43v4FfGYRaer/y1
fWVlHhnTG5Cc3BRG9lyKqjor+BXGV6O4htMgNETjZFnVLRnYhie9OhBas2t9TWByhzXak6KtTKwB
/ZzdGi+uONtVTsMKNX/XNmJprwhSOKla2m5liGJsg9i4cxjTHNsUUlxbWMzgjW5omGlPRQY7SzPS
HcHI1diZncCYVPKo8AkYi6jOaifJIHtuJylrUBhjtUQK8UNs8DomlbttuMPJrTavbY4Vn+09ebmu
cY6tm7aky6E0w8+Hk8Lv1SkGCQq+RP6DnD5XRvRczXiIir/cpmnUUkjxlbW/tgxFbeX5TVRAlqZx
C3IiwHhS1dl/IZEqiYg9J5OHO0dTS9lN2ZThgImPK5aHGO3rCHfxXYA0refMTGqJZe9Fv3x+Te+E
2pAAxGHPD7sJsbubc/Jwlt+CFkUDeH5ad2/zQa+73FLhmHedqrJkeLbbqRv2pPlquzv5JnYuxzGI
wH+9OBDbzqMQsY7bKy/42xXIfCzxqzgsTRPKVRzC46br5kgo/GzzBMNY4UCCUzPPevnmT6OFYwfo
k7+g+NRbIGPctso/syqwJyIJO7mHWnGwOdGBpEe2nLKj8yJZHOThBJNrHEofH74HTwrLuZ3qc+76
jsfwY8M98rAKwccts3VcTy5RRuznB7QTPwZQNKNSGHtLIDyqbABGoTWSoNWQ/mwT4Olg94p1gpO7
sqdDcMYEFVf5/ABaMQ8sqOoIDhh4VClSRhfn/QEPsiO9krnKDQhJKZmsp4QCjvq7OTrZfmyrTn2c
FtTvDORgpIDgzR/i7xESvvZRK5Bc9Ulzb0ZZ8bxq1ot0UALGY8kbZ7Z90HnYlMwXyP1r73A62XMw
dDRQxmbsk3aeJltaL0nEtuSf1ACEq5x1AEHJM6daJXQgI5gkibiYsjcOxMa7QmJeItDPzyd41MyW
Iyi9dXyDpwtVuMJSTNg7jLJflN8Vgh4+kBB46fsunYrYhaPoMGooWJ9Qb+WrvGEs5gC3XbmKjuVV
pII4dJq6dE1tnuS3Hzspn76o8tMgOkH13ga97+BCq0/ReTm+vUYcH76zXNr9Be+SxFMmCaaY4K9M
PpMh5tAeO7WOJzBldVo8vv3jVzS+AQSGSAQZKskcQGxbDsyxtPxFYsATyr6uY02jN2TLwxrJBKBX
hkxkuoH77/ufp4oYghi5SROFLaNC14B0xcgBoP7mshZb+iWtBbS9EPioJAljWCWcAUNlZQIgzTjW
9J3k+Fc8pfFYemaWJpTqIDvvf+6TXflapLZ6Fm2Qumho6WiT5nh2Ds3GSVvK+G1gLNRdwY5BjQWP
F3mj4aLLEqdCWprmb8RKpOnbuVkFxgU6Zzy4DDPp4F2EplEVJ/ggvOlZCSFlsxZTlMG0X4pT3jxS
+b6yMRTBPRWCZbUa0aceI7qDm01Z3R8tdfmuE20jTSfqpzf6CQemPX7r9h78XUxnqGtRxDd56RzO
Jzyhg/80R5pRWwk957EPa5umPHEWHApN2sQhH49qDgmfKjaef0EZH3dcty35SypUq/6wBhYVcJ3P
3u0vVai+3pUJMTxflYvLBRQMDYG39m/DQX6Wjh9Q5pzdcHVEhx5/DUSol0jBkLq7MN1LDJlCaEt0
Db0ce40+MQc0aBI8SUn6HvKbvm0/8l9qp9NI4m//NBVCXWq83PR4Be4rYA6z8vovK3H3+7+R9pm9
HQWePglpsQluUCATbblEfrIz506EU/PXos64EmPLBCoR2TIx2nob4XohauVxtrhi/YRw1j/02z3I
Dzu3iQau6VoyfdHlZfR5feoCsyMdrmAZwkGv8C39jrAwSNg+aYRlFf1pEvQB4BPlyckOfgiKUtnW
/mHdwF4d/AmRa0PuS7WHCJUOdJ7UZTEaSwE+evrhqVB2REzK0UAl1qqi9EnIJqDPtxVcEBkMFpuo
hssOjhnf4Ldb6xpyZpRPzy8jof12L7PfM0EbvWKepzBmJLhAVXUKClRUD2kv9NjnQ/+++9sZtkbo
YDQPUH5Nbh/llRw57GtuWB0QHmUNxr8vBYA7PJgDZC29/tI+HxTpraY824eHKmlIAeuJqzozl05N
lMFOCPxW5sNOswzf3kceZySWCJWvKUIT6slZVFPwiwJtJzClvrijgvomipAZMkOwkcWkgGO58u6u
y/OIbMupJxW6867b1BajahRdmY50kJNMiG8dbTVDqQCac1Lnrqf/oZbP2fP1oDClfRL5UwULU0CC
PxQ0Iu8aXUBawlqqf+7LD1K3jn8tdXAewpIyHyiL2jT4/yJQqCQtYEw8yS4klupmsIssoB3cyDrV
mCRZ/xYUPzZ5W72WBPkWQCIpC/zhNx9dAkNM32Wr8kftM0mQGVyCk20Lpd75UXl1JjZzghOwXsdb
8yEIhw2CFLsHjhuDE8qtncfEN7IgptiSG7E/FlrsZNI9pO5Fg3R8jsD4R2oHfSi07Q2C/0irTFAB
iNpAaUYnHHlp2nNU0d2PgBbwLN2j/4vXb8OQ4KhaB7RRN7HTxzVU6mzUKR0eeF8LMDC436XgEJmR
yVAaykXR0DiqUL4DUB76lAWIr4xKtg/eFrwtWCgFjS3PwCrhnzs1vas40aMSF0Oe3AIHVQ32tfA3
8RSRNvvJ45Vc5tPCwhMYmETHy2ONHfsv43juCXliO2WG/I1fhpX3m04jABC726v5BEaCJwu0cMMe
Q6+GMb0D5kXbiffM8Kgic8f0Hi02Q0ZpR6xnp+vQGdxvCJw/tQadqzbPv0uil+RYtvky7AMu94nA
F3LxYQaYV+iRujduP0eFc+agyBS6yfUuPF18e7XX2sJql+GHAuYWoLeKOfUvKyU5BoOHD13hXjXo
svNZXSIE9FI95FM3tVhyJdCCdEes/RXGl+NOZ+Yb00mkOB4Uzy0aKVGooaKJ/jeU33/hCE8w7E3k
hmhK43cyUxo6VrSfIH8CiDPibXSRNuc5YH8bLiN7XCILVT0QdLhY9VICgomdjNEaQ4wJPFEYSz9+
KfVnql2Pla4FUdTvpHTKaihwcbfNUEUMGxyFch28rQoE+ShuCHguDpo76y8/EyxWQaPXr73boLfN
9f0C6bF7oSl8SJxuNl5rJ8leLA7U8CGPQrN4/3E0JP9LNizd8rNssuwv0dGMZOfB9Ko4JrZj9u1D
e62DeQFUO6NifJ7C1tD6wDgCIMwC9BvuG0YXfBKUIJ+GAq4JInu4nnsXwKXavW1M96qx8a3IsFl5
M2jWxioToIADXHtA4uhg2wpt3hFey2P23/LLYqMk4nydun4kSgNAM5UBm+wzDtmvTTsRCGmBzDps
CKArTi0en0jlOlJGDpAYGulVHJ/jxgt+OtrCds/G/fB8gwGUXTh8BupMup817yWAycw2bxMWNYtV
tXf2IYKrckfuFQyOc7iQZrBiIBvwkn/WP8HunUQwmNUnkYLtQemvsagmjW9GCgnXkbz1NZ2orkUb
imElfw+QgfGG88Erlev/5Qo0NbFuHdvoioR6nLhGz3+A1aur2qRjxZGqfRhZoO/+4BYyovz6CF80
mMD+lLFhC2TfL6KqxOmEjHCy9otbNzdPz263WkMPTqNFeljfvrzZRlNSBhxo1Kh4+PzTziXlapBV
fqTetcxVH9iGFIwIkcO7d2lEmol3CHyggblQY+GQaaSe2fc6WSv14H0m/K51qzU6ysf8VB8hG7Mn
NsZbw2x4hNEHtDgyB1yczVvcSX0rS6S02kOnJyZBsYAcOqU8sJxEkuV+8ikR/0v2uA9JxSwL3Wf5
o6S3g5Lmp+Nrb0eSyF5Kv0uCpcnAmsll2yHGCOUA8llUR4iz7QlySbiUaG6iDa6qMbvlyc9zwKdK
cjAb2Z24/hAHJ2i9MU5VAs/82D1oNaAxyUuGjOaMU7dbWxDGd81RNrEqRIsN/toz2TbsRJJkhmT7
vhnQuhCe8HnHl3VqR6kfjfy2HgEMefNJCleHX3mgC7yPJ7Bl0ApjvBWTRC2sLRxs5MjC+2rQDOtY
zInI0gSUr1Dj52665rWYzrKWJGeHEImTzurRIg/hxnpVucUf7gg9elcNSEeXBS2j2jyZ8RiFRxpo
UYTCpBBsRAkPFSLHpcUxvDYlib4yRsG5xMd8k94u1KdQ/NDEfCTXNME946LGuiqDnGUbMWMl+jqB
pTwHfS7rlXo7FrWqGtLQ9maeSSdOoiwsRxBYgKfXD6pdtM5cVnD3J9chdSOpIZl7067Fev4MHtJQ
fdXsHy5n8mWioMdxdhPo0BZ0fKvkkMiAzZWU3DqewXsGW5SfDJVsaUvDuwPrInPb9ZkKPIczuVWy
KmyXSrm/3kFWQToIV8iemTie0sZNaWOdpZAzyTKCW/kO+WddlDMO8HfKS2KN3WBzfxEm+34pZ5Uf
TIupcaOGUAkdizFhIaw90mUn1DoWTcr/LPyA9Q3h/coHVsqSnqoH9mvmWNaO7Z0p3rxxvp/P8bJB
Mmw76fwifhH1s0lUtfoEuRoMVCGrOPPFX7eTAyuTD4y/NTKSySJnT67me5uegPj0aJtxI9yXoahu
yGMq/z4p45/SYBBTWrpPkMkqxzj8iJTSvQxPrN2nYzrJx2mAS6sT3qabx33JgLN4kheuJcS5NdX7
6utXSyAf0KHq2tHUKP0k6m5LDiq5Eb19AI8Ge7IiKAde82ytSQdSbLAJiQsmW07OKIFJFFq/9i/H
9Qv3i4bRjs8sQbFULdCbDD/MIfbB4zF5me1wgB9c73kRYMK/iGxHsSTqHcHw6COdOfLYVDbJu7QA
vRQK/+xax5oWvJc6Ka+UVgyEp4GF8ZxywbPl2MMSzYVPHlXp2+JoZhBrzbHpGdzJa0k5lkkWzxlc
7GbtTEdougsEWohYXvD0VEPzRXskPO76eMB7g4quUCMzDlKHvmUfYzTOV09xYgxjpjvbn8y7JqB8
WbPrR+rKdJWyQ52GOQFLJJ0tcfn8+35g7yroCalq4ioqY5u4/8wOlXVOuoBE6kCOXhytlprlsI2J
j8N72vcpSdAM3WLwbUFnFV5AppZPDWStO3W4NtBKcZqY8t0r52urCAVkDFxWU3av3i4BBDT88Jxm
2FVp2B9XkPknq5/I91j5Mq1nfF8DW1cWSm4YeO6CMsx4B5wEOZgeEo3XWQgnZwb3l0+h2NuA99EZ
AS/DPrRgv9uJJMFsiPmtXH9bQOFyWRilAm98arl+TPX1xg5pvER5uFA5HIgD1lwHfgEL8NYMaOqw
u79i4l4Osp+lEYWx5aGbws25UWEDj3UNCfJZIC1FJA54c7UDDZAwQuggenJ0Vfso9M+EHw+8uZIQ
rPKaZdPzFnH7YNreVapKoRdSe1XASXLATrXsOsPj1AgcUOGeEG6Iytdb2ZZKmITkHEorvhjRkz/W
DJ0h2MQ0KGpcpj3iojlJOpP1h/gMJfx8+iVhFBuMLbjh7us1mu+CoiFzytAyaC0gj0ak4+ffJidO
kPlJm8wWEe8oDqhngiB91z2euFh/3z3ADlcLLbjWg3bpG+aFoVQWucttkd280jApR/S99n7qpcXe
uksBRtY1vHAaoYvanFQM1h5+riL6f7/wBohXcvLyeddqeNwy5HbQpd0Bat1OJpVgJNTMGN84wNap
iq89gEo4+0Bs2UEVCpEjoQMeZNkpVL56HB68PmqqaC2o0m6KJYPO8OXwUeINiUuKYnjOsIKxydc+
PXxb0aUqd2NLGU6dQLkP4+g7k14EGgRky17WjELOss+Jh4HSCwKOfGZ2h+yYZY8jBRg+iaUWqrgf
q0loP6OGb2uTqMK9aIaYuRREnGJwT1p5RKCGhQLQ9b6xkDEUsV8oybWbijCpnJ/KB7H3g5ItdBbi
Jc8B6J+h9CF0KfJ07IYG6OTRAkiALZ7C/wl1/tHTrJShpUhbY/dUHVTbbkGcZZfRrDX+BzKd8F3m
PaNW8nKmHrr5ExKjk3SbRDspFaCS9IVRxBrkb/4zrRi3d7SRL+UXhE7g19kmSRr79fzXnommam7q
2rl34h/FspZBobzdSWyZPKJifJY4wnxP5iHMTRTY02WOj2uBqtHVu15gSG5Wb+a+hCn37mwM3eBw
U/DtP+6OmeRJgQmN1TulVbOvaQnu7VrnJfm4dWd4eCE6KDAdmTzFM17A6+nCF0fZ6ucnH6UAS7Wh
d1gFvraJU7dMdKkrwtaWAz1RpPkJZuwlMV34XDI1cubbiymbtyj8UOcxupywXzdXqOaL/aNPWdLD
r03xXjYvv0T/8SSpUuvcYj7XmLpajIdQ6B4BLnu64Qur1NorcyK+wveSpxJhdXiDnrYctSQrxZdK
xZnovKsjYDfSq+WpizASuuwi1LYM5aibW7pAT1Y2Sc8XqaKSpcYrruxSC6PMShwhulqdwKqgbqcB
3bcnIqN2wXERRjYUlq65Ggki/N7JEkGVAoGftFwZetDULnmD3mXclu0X+PBXQBDaVK0NV676CnQp
wbvyy31yympzxekN4qbWv+8n67dhGuOMEp2cpkDJy8EkwOuUyWFw0V0cI2qW9NKLfsZVgPSqUk8n
VLspEz6rzfGqe4zvpuE6dfuGD/Vb+mavvK8+mVDszuVnQWYm15q2BO3buugisgOWJTkpgI7q5Cre
ml5SGunbho4VZ4UOvLFd6wIYFDh/sUkcKSnqpcZYCOLNLLe6EIIVRLmhXEEjStMYdIOqMdl541a8
jfev+iY1n5xYu4EQeGGEQz9kJ5L0QBXUbeV9rR+JvieB/cT3AwREpRzftZa7e+2+dwSNnQGr4RPz
dkX1EIgJ+KoSm1zv0oJuuSckiGOEelPBPWWCbA4qesL16M7nsVbGTKl5DVhKpJsKgJQlLP4cAGgS
VxSEuIpYm3nisX7a8rRfvqnEmPA+ubjxkRhI6axO32wfk4q1sVGvdNNuJnUotnxh/DJt++LWCAMx
ZkxOAeNdHs4cuRk4WYNlJ6jUoQ0oe4QcrxyYxQ0MocezcA6nrKWM2xSm0QThXo9aauBYGILPkj7Y
y3gHwIJQLTWFvvU2cJeb96SSYLn8nnyVjA/Nnne7JB6HnulE2SrZRhQ1rxZK2fDMI7CwaNFePzag
W6kH4xV2HcXJ0zYOYKRxA0ibwjK3CAq4437M/jH3ogj/I87BYvPBtfVz/mJL1eysUjMQ8eHM1cYi
sgM1IgJrAcbmk9VKFE+Wjq6fFla3Hfr9zcCvhobo8SuLRZvUcKAkPeEbMO8iVg4CLF0g6P0L8yvV
oT7c5Prjvui+xnwRnaq5FbJq2f4YJgGVqzIr2kgr4QZBSKkWWUVyMjrNuynFwnRNR7CknI5bPYai
JB83g/jq9CEubL2J8BnSef6dqSNMiSHiApNRHd1ay1aZidS8WiQCOZy6A10zwZTqk8j/dcjsRbhL
+lm8z0Z2YrWIYFxBPrazEu+S/6iEwzLPWHlGiqjQ/u7BhEkbDuUf+zXfVLeuBFeRtAo3ktEY7vcm
WTHCF8V0faistU1zi4L2ckHJB6Vuo/Wy0ubbhfwcQOmeub+hXfW17vfXzfTlZYtG6RxPe8Uo3HzR
b/lKJt+Ie0sTYHBxWOEVRUv+HS4DlxcX1/z+nX9jM2d7aOmwLpy70eaqeX/ONI3YqGO3JtUNq2eB
QzUof3MLpz4/aDsM45++ERdy4zQ96D6kfUjmHBrrj8FjSwi3569Vzv9j28UgWug0bF909BYpPoDL
HuUVnIFTR5JN6fJwlF68R794j1PGvEs2wFXPCV4rliHyyUhu88MBAmYJzHdDlgBrccGjJoKU97MU
aho9u4JJy/t+GKafMnLr/fW3tJp4bwg6uzkYxffX12oKD54vAnggai5oMVE3FXdfvWCAjdOF4QeH
Dk94Uzp3gSfFbinxNS+xFKOzyyOpObRVtw8FjEHTZgJHu30yufm1oiXrht/vhNxe+96xuAgKVMkY
NczJZ9xHoJY3yaRj2ODE/rf/ceQRZO7Tb24gqV6uE+yCdJ2k0VKm9h9etftr09BCiJh0ZVfQTJmn
IteN+RtXWADPyt+ftfgc5n8lmWzfJZT4xcfSman93KWe05Kz76AnVz99V02UqgfFc1BLo/ymrI2I
tWdABxV7qfftwex6tL5TexS9KBUfRdDTuUrRZK0huGdnDsdmweenqCiwG/BVVNtWDnt6RxBVGi62
Fs1Cvz0kkHVzFkSApzJFILDWum16YiQyr38rugEf7lkRLF8rtGpbwZqADhP5V33wdhjncDAIstTw
UQL53OyZdWpzqzxBadaCAxtAs7OJYhRCqWtT66c911GuyG0rGjqgERlPC+xlHqPAqSsMaEM7i1SR
vKr+l1RmYLk+Yq4s4WZ57M5PQVYs2oBLZRzLmxVSTSznR5il0L5fWPDZFj6jUJk0qKJNmRiEr4Lc
xFmUzkAl4xzJDj3LO/VPxNZGm0UfSfcCObyLqjwPVBFMNpvU1OBFdZooj4wlkEeyi9d6FMmP5xLl
coL3SiBs+WXbKDh86srD/xONuSl8KhZCtRYEUeVrjjyXkYD5weVSPCAbV09j/fO9fCjV3ojosvNI
tw52D7gDOIHwQyDKmAvWZy6SsmuinQSXsxsKrNkh+VfX4Gmllg+J50AmG2cZ2nhUWXo9TBjUzCsR
K3yVPwylsZG0rgNBtq5PnwzqNydZpQMVCUKHrUABJy7yE9HLduVrmk7AeE0i6zXWuuBG3NqxURKk
IPVIQxxoJFFFtoZncgB0Pp+I5dfY7XYPGaf/fdYjU9xTOEeipd6NQyHBpy4hM5S7fTB8WDXKqFNp
1PCH6NBCEtUiXRVgZlBZNS7oiEMX21GMTuOgORgDxd7zf1B4n8uAH19seq2/QffFmA5usSVzLNqz
XBDwBI9737ffG6jqXxdA1nCYT+hwMK1WpldersxQp63LhfyHnicofpct6bcuLC3uRjlk+8f9oFMs
IBynI5r3I+f/L69Z5HnkBLVoSdFMTJo2F5A3sg6/YPdzsPSDjuVv83iPd22cHXeg+79krMdXHKDo
q4ZFxNQZkC5hV/6CLQ0qga+yDj6WWOUvqiC271ImBFZL5ndahsEetfCrdkhUwJAXLg2kuFYYmYXC
64wwS1p7xTP/zCV9WRx1nDahUHhppHSEApS1Dd1i2zAGWlMHlKJeKT/X2u+iUX15AyaCca7Uuikg
s1HQXSy9wcITBO3mkNotYNOWUQhqwh+P9/Ab39A84qxyQxvHmoh7PixjQ1Kzb4U3RQBMfWKRMie1
afKB4myCk0A6NBULQ+CpMZ207eC1XXADqNbWVHecNQDVT7Mre1Sd1RwX7KQ2Kki+E8d2WxHsWR7H
r8wOTsXxAA79cLO/4CSXEPacP4sKv9B9QXShwViZe+VN9c6TfLjLbZ0l2a2kC8tHuqRUbryqe08T
k3Gx5MQ2fH49vWnhr9lwhjZb8XaXak/Kda7otn2g9dTCmjVJNf9IP4Sqp/bN0qft2BwwQv2cH0vQ
9X0Gt6/rBmrOZpkWYrpdcSmvAnRoJYX/yS6zPlgL/i85fkZV3GxmNK+gdIQ+Umi+KcwHfGSr748E
Ar6fxfcZdexK/VJiz2Zvj1UfzR1v2uAWfigVMfFRMuYjPirWovD7Qx7mOFMecBUKce02PEoUZyYu
c1vuNKKOe6D7hGRoQDwY97F9xOEJDMdl/RRg1MJZ1LbxcMeh7fvEJcHVmVyUNLcuApZi/563gvDg
DyXcqupNhyPKfNhB0bymuJSF1xndYiVDuvp+0zGAHaaKCX13+hotRMwKG0gM/iWm2WSG9zEs/iiS
kY+g7wHj+UP2vK/XML5ZEDLS/qacp1PjUDpWLQahzYb2b9ToP4W7rMy2RR4hBRzU6ehUaC5atdtR
SycSggfOaSW9Cax9NXoMzn8eNFL11wyfBdC0YdWXmxGO9vjs8s9uaqeFMAv/u/hYdVUZ9nngwStt
FEtVbuOe23JOOW0Vy+M1/Tnjs9onQhJlku1nesUXL7TbCYFfM+8uuhvjU5otpYyLpACNq6w3Tdo1
+kwarveO0kT+FZwNEkjz9HAEjoFCNC6kIgB8FO+X9NJikjT1lgPBdlDe3iSjmF1CIvdiJhYK1Sdx
9sBLxDD0k3c0Nv7Joy0hnYnEaYWMeXehB8+vrZpVaHI5j5X+MoR5jkGn0tiNTjKrFe7QSAx7DIxa
VrsRkQJ17E7++BttqKhbVcTV/c6cHNYXVbvl9CavhxWcKdKgUlYY0QkfCXXEvJWdaQhhSBBlu99o
zp4X/I6r++3iWFShcQdlWXshcKpysDEN1w5yVgikrQ6r15bxaxoPUjHRWIQbTt6+8otBfpk7ov80
FPWgrq2LRPrQpEiNBvWswNxRIiRHqxU2Op0agflui2JvZvuAYTWsf2pW1dyKMive6JRploU9bzgu
7QfVNpGLJpbFTFjFSpMVd0eaYXpuwYrjSOx1ay16UkJufXJcDok/Q8jd7OlswvU4jllVrAoT1ND9
4uiGl06OE4Z9rw1TkaIXPYMJySpFyVIuIaeRMXiGAwiiJDBl0aoU1yBRws9VKdViVvEvjCqflAhf
0IEIniH+tnDq+1vqRbVZPm87te8cf+2Xhrz7IXFXikzkq3ug+BsPaBGfOrzvRFYswAH5vTk+6CLp
bRCtbMBy4bcPhjWCGA4mox6c2gXCblYixGXyIf3PjoJbEht14kFsc99Fpa9mYJrvoI/3fizgkpAm
j0S9+vGYN2TOTUWmst7eHl7xaemjvNCCca0Ca6jAeVbx/0pFlS3+8PYvri4miK+2o+I0VtCRwA5c
VY70THZKqPUFHS7h+XlPtQ8pLeuvULkUr/fnxLcAinXLTnpQLimMoPypZg9lIG6ea9NemDUCJQ7j
Ugq8U6eGp5HgfuKdZ3W3P+qIY1ronCQYza2UCyR7PD8MkSNQGa8TQwyaLFNc7MTHKQoUimFgi9+4
jTF5dKnwxlCact7xAjXqm/E2QtqqeQqwc5UDCYZfoNO5Ndkk5BOg80h3g00jzH02EQ/TUoj886u9
PJIlBNT17XjxanfEiaxqnIG9PFoeHfwwFrSbhvlqeCzguKGsWwyH/M79XzE6spymoQiabLXOg0Z3
XgGMxQCv4vOeYACKiNu6DMWL7YQT6WWPm/NWN8IXcxe8rir2YCEjmA2o6rhbnOt1DAouyW7AejKt
KU7+3Bdr+jikcZor81+AJNCOzovaMp/veRMV5mhiO7DL6jccqkljhkhds1SbZXdxYImEBqhM1pCs
cFcc4B70O97PuyxGf6KVjSecCd08DHyzyhDdC3c3NLKWIk5o3JTqQYRpycL8H8mhzfYYXapMOJiS
uinojvkc61v6Sk1p7zHPSUmWMq6u1UdgbLtooMNZvAy6w0GfINzLe/E9q3sQe5PBaDdTq1PsUnH+
KYChQVAMB+64otZlrF9J8EaD5sZUTpXtAWaWy8CvZTXJfC1p8ewbfoIQ9EmMViEXtzHlAQqskuaO
puffJzm2byq/zvgwtuVDxzHiu0d9K6l8I+M3YMA7HoAfj1W9SMROJHJVw65Rr0MEitZNwR1Ybfs5
wJaXm1xVoygy4SylSBMMqqaZNPdms762I0A6DiAfJNiFa2yOHdRTu+806lqI91KQ+j8mMrLDZYEQ
Ar82swIfLWsWDdN8KOdUuB0qckHyZitngj+XZiujM4Gsz5+9K8Z4rY2FBnPfWEg+jciwP00mNVEn
+3t17PpYs18iuj4ADCMti2CV/8J8XMrdjEMC7VBKXk7TEBKwbh4Ck2NNuG2CukxrH2ss49psYx+B
RY4JQnb1mZUiTSdXyZHCTeksu4tNESz0NC7iViJ0Dzkv9EykpmdPN/m8kJv8aYx4oQrpgx0okmCf
QtdbLse1CJGucNQCeiRdqAeqaY6s5idoLGU6Gupztq7PX7SZnXn1iiFyGMPJiP/LwZB3DXjBBXBG
KHM8AuYsEz+rf22DJ+/323hdtkVFDYuU74GEzaPSr4E7I8hbDDgzEmqn2HdhvfBUyNPkjWTDsBHJ
s9C1tYlqf56UzXhLKiEUSIH7i/+B6D0UZjxftaX5QyZgpNOiAnf8jaBWOi0TTWUOEuBjCJTu4rb2
Vkl/vHPeXO93OJQU1PEdGqheNqRTl/LrYxUcledtDxkSQGYBlcYrGN8M1L/ULqX1aOuycsQMBHal
3+nxDe+JXnXWobEDZx5TeOyi6Ifj8R5lTVq0RJXHvRfOBJv7l+fMwv964BJyGdM8+1OHkOE4SG1I
PX5YYtrYDxux3TtBifyBDPisYjXyGDOPCmHUTV12kDix1a/HyiN60oRIu++7gBpDL9qSdOuewaqF
IZ0ywWeCvOJrIhUADZU36cvSN7p6ygncgVJoX+eu59X+RL5mx2C6LoDj8XdeZGLWoBBATIfmi3Kv
kViW8CkwuTMyEwZC4NdRMSFMPjcMd1hu22U/M6OfXM4P2xXOdiZSTgAhQspOqqsBJynvcp/MIrsn
tIyKIqxbun0J/lemunrFBqwuWkRBWZv7zleSnqavE0zfR1aZaoHwbOuAU8EhG64RLyET3WZVRSRp
vOFVTwBXGENf3tmD6UtfYEkvoGKzWaoXd6MjPAtzIiIMYPlhIO1/8P2+06f1fOgdjqYaQ6MckNBy
G5auUXq/9AGbvGwApeVJaRGuc7VGE8YLbl5YSbkAVwWnyP80D74NiWM6iU4KxTOcyxGue9z6N2Ha
FRzIhJjlslv+hBWRaNPgKTSX18V1g2v5X1QGSdu/vQUZR1Vk9HU5m79ViPqWVbqf15jRdE4HRRZX
Y/LG4M7p0VuSFR5pzUDYKuPpaPsNjizKEnFi1sE6jdzqswir0YQrL9VMiROorG6MmnrHjBHQ10gu
k1z4a9jrrtyQzl+7SaFjllmphfMEFKP7u/7NthnJO9nEz0sw3VIz7TIHsaoKjWW+VYs70hGRTlOf
vsacJLuVHGQf4Dz3v8c/II+3e5dPVulGMqeQlVrIA/XZb+YfyX7zorXjSM2hDE+xJOnFSAQXpzsr
WGZu+ja/tBYKIEbbTeNrc6zloE0qFAF5XqRMNsMnnVYRcwy4HaV4Y7f6uCalo+MJ0OMQffPKtc+U
dhB7xTD1iF8AFjqeyV9KPHM8KeU5C5FYzGOJsgHQv3gZalRLq/t/w4ys9i2lPBQOdjGzYR95aLEZ
X2hSHqVpog5D+cnPHDHdrDF931DQFwEX1PGOiwDGEU1lYOnGYqCUzNRJdqbGyX4CZvKZIv4FNXTI
AbInVDh9DfFOadmoUC4dzewHPddgPFBAkMkYwbwYsERLJYyi8o6FaGn0SKk0hggikHDJXnYBt/S1
28VMRDeGAzbB96ulFVcsewil0ZSoNYXA0uq3WbRVA1ApyYzC/R9ibLlHMKynVLyhI4FhIpNcI+1e
JTnSQdI9KolrpcOMLXZMLldBk81AqPESR00atYlK939J20M2FBoEhzm3fa5sj+NPBweTOXCqIxC9
h9WEbOS1mZhgqm6+K8P7dft5eAqbpyccjsNXmKyeJVgsIrfL4ZbBqTYuE+iYtqNBDzAbKfSvSln/
GAwO/yZx8rkHUFWGw8DBx+0LpOW6eDb48qsAtFfreouSsUTjUzLcDlGn82zkYpuAA20rPRe11yKZ
ADEkb/77JgJaS1ITtm2yFYqUtF2sdFYcCdq40lZYILso31+7Xz9C+e3OO8SW6KTY/2dMB606VymS
XMJo3UZQui3HUJPCOw3iAz3Z6mLUVt7BRRC+DOwx2fAorVIf4frWtcMZ6r9YT75jBBzmARidwNhx
aC/8hKX3SWxfB9zJn/xcTmXUiSXnxf6cM77PEvJC5SBmHI+hxPPexYOWui4dVHoihuas7v74b6zK
63ZbkJENCWijS46YvCqhM7lKQs8OruXrlF7MO83lGJIUlT2qaTcj+oofb3W0woOVspN2vNB25ls4
YAq/5ZKiHVLgiGQvnIRWcBLzmk/VLAkmk7Md8UBFgPkX8YgoxsAfKEKyFoNFvX+xBPdxBq/Sm70U
9ZdibwQ8y38OkeIrcDYSpXz/HsFshUep/6UXVvc/WMSuFJKxQjcegP9lUJ25YRmv2NxCeaY/1IaU
6Kx+EB+wrUFLAxsoHhi+gOCuXvejFSxu1ySnx8HKwYA4R4W1lY1viR2M8PuChlC2nF33ZVHXJ2nQ
DxarSQnqlpDvrVKLkU2no5WIDQVmbynt8DSAEWqJngB5ZQVFTPDbPjf3OOZnWb+g4ylAEOal1IXh
r+ahBktvSdSsEAC2ipxUYh5vhu1j+0r6OxU9kBmqYhZBF/s74/sJsAtGTaDVGape1/a59ZypC1nQ
a4D88MU3fMEgDrq0KgimV80qiyoAPyZCyhwNF3cNSAwyqR+CsVMcIkkiGwcGPnCdGLVm2FusRjW8
B2vMSrX2MX5TTJqpjhQcfRdfv5pu/zQAEnVSxZzlxA9KkeurwNCXlZH9NrHf483tKikgz82uYpcr
zmAqP173dzzYrKulO4X433vMGW3EBZkHDoF3OL2nH23aJzfyF7QGWCQPpQQEUdhsxg1x+qA6dwQV
m3+P/8NlNIJxzxtijOTfeJfd+nyUfR2ZCFanVjxzJSKuzL+Ct1zfEIR3ffngBmiuSyRUbU5bYQRz
IA/4fNLcSS7HcLapT68DmS3fX7pLI1HUuNDBJgz+k6VTYN+0acyYZ3FWskY2A3HpNtvN/2zik8zT
sOrrenvlS2J8NoyzpLHEbSeF0JF8jYJMPOCobq6j7D0IoLbYOiibljzBYuatKndGDJDPB+++UTuJ
y+GSDRe6P2f7DIAVe78um4Zer6v4q/qudlM3gSdq/mVXxUU5msmjvaXmA2o46Ez9uyFccZOrHDEQ
EFaFOh9cJI/8L09LsH3BU9gnTzzpe3Y0D1hpP5YfrRGI1pLdw4yzXFKfnHEyE9cOT3hWlmMxFLSP
6xo2+MkB2vhVC+Tq5fOO/otnFzBncr+pwQBjXDvLwEm22FtdlQ+qH3fsTIW0UMYVEV/bXwN0NUg+
FSe0yQ9TfVRbenHnro4OIizPQz66l6HvZtj5Kj+I+IFtpTmMpGCf4mY87j5pHG03Sn1c5cys+ugh
16d1BadISCfGGGHOfOn0lIAzL68iqa4mvxE6ls0GYHe4/ymZ6liKE8x/37jip2+IovIQmiabDtyC
3Ru1E7nU+eBK01YnsUxKHmKZPfvQpMmGtfN+aQPq5woabaJk7J5Q/eb4kUFczyux1u10U8fT2dG8
Nqkd2o5wN4oHfeq9lwBjgFOnh9+ei0Z3z9Rqw3zd4uMZSC7FAqht4ztzl/ELMdIuBxTSJ9jiUASe
w1WnYXBc9X+EZybEnUwa4ZaMczdCqWfvQOR2HPnAf9Zzt/8zyXW3QfJXBNDHqr5zLsh+fAoHi5aL
6exI9KLDetduu+CAaCC8xj1IDKZdu/QDqxB7yed6jOSiTVIUUer17bE5JwtDElWwpM9LRXFkNhj0
WY+RE2IYkH/QIwHi2zRrX8hL7ief0FH4m+MaJVXMltKIxM+Jof3IX4tyryjg8pyFE1QDmXQXeGij
Ns7vatC0noLvq91xL+pEOCRIUkyrmh9gw6r0w5p5h+dwmMahv9DNDj3zP8ZvLIo86jhKtpKvPKd7
09EPCG2ELXFpqIZx52sT7yKI31aeHcPZLyR5qUbSpdIuHnA68X0PpQi8Wj8jdJlbGOsMNHRITdCv
TOqyiBxfRy2Msv8F7uVyRG3FMzIxYkUfM50hLEsa5U3kiD31pXL3RwXJ4aTV7UjagZAg31hB3Ild
R8u2GEXmePCvaPYJUQKS/PSFf9n6gu3Y3Xx1yhQ+WqU780l2MklO608HvMmeqIIF2ba1ZZlgW5F6
6R4EZGB3JzF3PFttbqEwzjArAreaUVIh53RvKsJKyai1S/UWH8DXNw0RFueEO5h8DC8ScLyX5xgr
6pn8IOo8TWqxOLL7OffYMIBTgvllZ5enpdzNAvXuHM95eW0sUOnyMI9wR86+m1mH1W9Z2CF7ccOM
4jmjwPE2pgnO/oPnZlFUNt5OcMMSlscStgTIBc7vCbu8QHX7Kn6fqcYD1yqzNfoJ9k/68jmPJ9JF
ubiorVUxDc4NFYkQYg1XMoBTYrJgxUuwUc4eHkK/A9uYzvRrTYKo2N3lLWdpGoD7/nuM+8PvrlUq
sVeDz/ivIMG61J+DruIquOqTOB57hODWG3k/dZ7Z8jqmK1q7Vf0zuRkRoL7T1ArTKz5ApG/i6kx5
yPDD5MnVi7RXgoa54lfAtWbAOuD8AjKX+bfr0bGB4MR/YitnTd/oKVoVY5og3Y3tP5ClO+krsB0U
VEqZuFcS71qdCihUmMh9V1qg0cCxims1ouFLb193uyUr+ZwIP1UdQvF9gYh1nOKlI1a4vzNAG7c1
q2CM2NyTi3vRy/j5k1lL8ASWqIOZnvMXadqZkHnPs79OEOeBsy+e2QlQ7BjWBLZD+1Zou8o39J2D
ZS01idcS5wxp/OVmHgemnovw/1EDeStzjU/3yDdY66DwuC9JFHJ5Rilu4GT3Wpurm9USlRh0PYw8
4W8Lwuy9mAq1r864Emp9QafoOdRLyxMd+SCwFuHpe44o4PEyUziPk/E1qx+rPh4mkNq/j2K3HM9e
ygkO6e2oZi3tC4WL/Glnf6H4MzdSKBKc2LGEOhLAH5Qp6owSMMiWxn3qmXDtVKiJVhGF2okvP6jD
iv8JIE/cLYY+E/ke4P8OJpFkzQ5XLdiptkBoEi+IVo4PcU8GFCk052KfUWriliMWlS64tYPVuXc4
btUSo8QEuJseZYBdeJfVxyf041ZjjpPqXooo0UbIpb5DwAeRxwkjI+WG2b5dsvdNaHdQxCYY8AT+
jdKfhVWgS/F/mRYSjGN+Ii90ZU1loCr206UmQaiBYcuJ4G28kqNU84ZSMMfeI2Ha5kdJwt+29u2U
zQwiGh06Lqjjt1CmwbAVkwNib4NM1JI7VfUGxE3ze4TBXvScJaSVNM3nhGM7uTtr+jFhiPUYCoUg
OhqgqJxoWbFyh4dojGcgIh39AZOE0QL4cNdkBjvmCMFCh/ODXqVJMTZmj0w28BhmYRSufA3Z8x4t
X82anIQeAm9K9361F75Auxyqyhuy50tor6mU5FzVLJ0P2E8EdRWIP2Q28Awkai1hFUbzfSMaRWMh
/9Rl5ajLhoBwPBPGOXd+66Bkyk7KAlWlYwORkCNaPZ7N7Nwv2KWsLv4wvWP+NRY/7iB7/wHS2BzW
0I8n8H/LTzomvpGhndanUlOo1fzPEwsCxyhKiv1fNPVjGPRWy1DQmzfh677UuIV60+b1Yq1QNhd+
A4aK52YMVBNVQDbA6AcQ7UPWJOcWdL4sIRy8WQaAFGpQarZRII5rNoegkDyW/5uRgxFuBLamNHfg
yys0iN646sR2VHZjqnXef7iH41VfcqxrFT/COlqZWD3URI10w2efrp2fa9MOq+c31i4nabNAqn0E
AsLk8MglKsUVvrBe9HwiKgS6hJUkHU7FQxjVd6axw50GHDzKflbxvA79pxL+8c4xpw0OHPeTZjJt
lc/M1EgKXMMFlWPqKadxQgsPRk1sf/56YXa8q+JLUtLxi1TqYPoLhngVy0cLAz2jWU/7ia6KMQis
9I/gNrcDj0i/cS2zckfavnxdCQFnqAkodHS/K4JnWWvrWeZkR3yzrzlRVWVayVG+2yjY+qjjfHJ1
liwtLB1gyzoyRjmyahRv91hFAQ2FNW7fixjrnpUWqiUJ50GuNJ0UHQSPdwuDgx+/1qPF7tRDniY0
cFWTppHFTsYu3C0XfOiW7kPQuDzNgHvr3znndPrj902II2f7H8z6sxvsy4goC8VwfbBGgC2ZZXVI
gs0R8bhss40ZS8TOpQu1s25uAqOAMShokL4SzDu0CfYihXOcYunTloX4OdDtCWqyNrg5gC1KOkXZ
jMImIMxrpamHFmk19lG5ujK5+XhoATjBO09Ba4ryH9M27mPOputQ4FQaLnR1EqTOJIB4Ac6UudIZ
YrkDMHwazJYGIISjn4d51xC6d85H4YwXjMsDgUgPuBaq/6zL0J8XNrCD004rxZSIfs60JgJnO6nk
ew5oTCycQydceRErbNJMhk83DNTZcJL7tRBe0yTCdBp+ARYgOVKiobd2XrBAuqCwidvCwqAJJ0+2
DbIr8umW4LlGDVFjCw195ionMjuVc3p7CewrE6bPGjrAo7uTmjdhS4n80XH4EYz57NqWSLPksJxi
zKZEQego5efST8JJNksgIGqOnMIc1gtjmJO+51dq70sQRh/iXMwanLQJx1wdZ2S8ZLx/1oJCJ8CC
3thQQg/0wUWDzVgM4Wjp51wbYZyh0E70b62kbBtQKVfs2quYDOvDajg+Xh6l54BnC5oWBteK6xLr
hFPnMyFu5beCDYvxFz8nA4TVoqR7u1EwW83PgAp7Gpwby8Y8Dk6CH9ayO37Il4TElcSSwQgZh/s0
Qxe6wK/1hx/PNEPXIpr9wUEQ6tzm7Gh2KWGFCi4LnV3HgoU3DJILLPrd0/8oP15KxkFJ4mFIzhaO
MiXEz6BLLpQvkQD5Zvk5O2UwQt1I1K6KHDgI2RYuiXjdXAr+guayI2RcwOECpmXqIHd903xtN5M5
MQRqLaiWPKofYXrlAnmGOnOykrERifgNKEeStUtFp92Pu8lqAcN8XLdeQfwFB4fEOkhcJLfXo/q6
/yZlU60KSaqbO5AcQpeqkRk2AAv0YHthIUFNAmcMh4ZK9c+ou5CcmIT3g9xBNVrBy5qBACa008HB
ndFG4zMYNf55I/JYjH3qKqaH/bGO8bPXG11x9X0uea70k/yAQXkHKvOUYOgln7HQnv+ooaPPUE10
Up9q8PzbSJ2a46YJeOHxdHZhzs2VmlALkymXe0qYVpqBojS0GWci9WBGpiMwGVhRJxZK5qH9kCFe
U46tYpbs+eB+47hE43BT26GAANsit6+hg2/N7tlvxZR1Mxn3NAKTAnJk1Rw6dhEOymVrH3H/sPtv
+IGViMVEtOtHVnLNh/1mDIVp7O6NWdVeFKlIA5agBsTbLm84F1NQ6cJeUfLcOZwS8jzgqhKDcpXW
5R0RapE9nb8+X5oOeePEx6WY2c3/zq4nXMZMV5plYpx4dJUekfgzkiOWEzfuhOlwg3l6f9XD36Wh
0CwFqJYeDQHEJkMrEP2ngAWsZsf4EvLNVQFQHHvhAi8+JUc1kJB94yz2zjtj5gF2rDfj+Vciw+cl
vu4XR41zko7yk8xq2r5CRAYgKMjZZgDLI6fAN37aJpOR570675h4PTe5WzBKxVtDmi/a0Fil1LTd
MA1xKXv1Vsn/JKS8cFOlZSpcvu8Jv/geN12GVYhTFW2GGNfaer41QROPpaDV+eU9lKzIQRWikUu8
nW6224v5foM9VkYgmaTKKBRFc1YpjBgj2Ls/hMUz9xvW5QpZ9Z2uzoPXLcpww3EeAu0EOfiL7Xik
PIp8t165OBIV7gnDpfbybrwddZyPlhf9b2yw2ScnuIldYocYohV6CTCwGUkZf032s/ubfDkG3CWP
U/DqE50Y/cgUEbI9V3DMi3DcTfn+tXHPQnCczlP0hhJnNrbGSix9wYHhpHsYNVyFyx/He5PUDe98
XK4IYAM/qwIWY5j9X3MVOzGVjvLPflHQC0XpufO41lWrxr3JO2TNZPIoWZx+LUmuZJajQqWjaVH9
SabZJ5Uoi353tuNgdyv6eBtYkSqSPn6hmts4SpQYf8iojrcpAmzrJHxamxqBeZr1cCvrVh3pgMCk
NkVH75ulR45p7VrM8OAk8ToeY7xzr5rDj2CfWelqE+QgPIfZVCQGdyS802k6n7Y99Fz0TGNZur4a
LEXT5bYcxs4lOXfhRcJN0eqzmI/ThDQMFTrpV9xVcXOecCzIpqDdvfKzxmUHUKMptLzyJ4kaNs2u
gxboDbocjxMJ8Ypx3hNT/itzVXmHEnsfEwQeSoQtLNeBFWP3Q4wkpFk+NKFQMU3eu1ZUPQdPLfpY
gHnl+DVeW+ErhqwUE0CQBmWKUfZ8kbWjXcPh42rJG4R525FUqaCZbBA4XOq+i01s07/sR2YlNjxv
5HeXnBa1W9XFcc8ro1H4kF3Hk0j7hYM8JcDa0MN2PrGEfegqo4J2UOGQdJN/2IQpa2ZCbnsF+kFV
9MT4+mp847QRT425Z0zt7c3W32IRGNkOzgRIMvW4tqSDwkEzUP3gIrePmVSBEYAvRF1oOQf3vUSr
9AbOK9vL94siJ4q7Bn9NvnyP/Kv1aPHMc43lHbtG6UwS1tGvG131UIBsVsI6tx4J0tiTNtGvvaQr
DyWCM7hG1UEs9iEoWrTwn14coYG2souQvXtPmWRNJpHdNAvXgxmqJfCVuPY25jrO0jxR2iSXzhXZ
R1rgefkpkYXtA7cZhzGNxbNF4XatilgZcRIE0SS2kApJ+D+0I1EYua0d2ypk7ohdBaTCdHOE13qS
kQ+xNXPU79rJW3XXqKL9pfe4IVs0eSAeCNeVGdkfr0uTX8z9vDwUJk29k+JmhjBtbHd3I5NFKmyZ
AGaRXwKJPhDTzN/gAlpUUjBml2erimqNbrGddvkkCaFylQoSa4b6cZk5RFSBmWbjSN9WWQGz+tCP
R/itpil2wdAv2USX4q2CY3pqZYdg11nRgtw0YT432Ukdh4advgToIQFBC3JX4nB1lVDVERE0PuUc
3Vho2LKsgWMhssHzLBKkFHFs/3kpcTwtxnpDBE2sFnGBgjB3eBlmx+qILO8JdjPUYQ4qvpuTayW5
qlxWf4l10JHK5OfoBixDLLriqE3bWE65m8w0geQ0USeV9sm8YIonOR/nYB4jGIAeMMdJmvl01Mhy
BGeqU6SiMV9prts33K7oMACYEi79gVnskqiweqUEsOVDdIuOCDjXqq+hjC9S11NRMxp3Y4nzxuzp
6YRcYSgSZom8KARNnu9zkdOSyWHE4jhYehLOxx8qEme3SSKjI/1FuQvfMOOEyewPVj2E9IKGT73P
S+J/iohHuWuk7cKlr7BbNejIgTkB+W9nXNewB5kQIiVtefmvqijJCLh+ezbF862lXf5RPCQF6fmu
JInym+zjO5WCU0ZMjYqbdIxXa9h5ZL3EYlZYdDYmAuzfh2y35yr38XY42NfUFj35/l34mbdjOyoJ
02fUX3QFDIM6grZBhlHs90muYZFKRMa7L2KrmjmbeilaUVaHh8twnUmO0ehfgJQBQHrS+vQT9K3q
AYyd/EmbpZDUJG9pgq51wltoXRD5TkTSzcIx6kXDBOVmohdMHmA8h5NizpF19QKjbGNHavySr3jh
fV8ahO/ThA0fQoSY1gf/Xz2fr16JiM6RtVClfyp6XXCpQbXwrtOw6R7dkEmKdbgh/uAPGzyPRtVH
mnUg2vFNkxnMFPeci8+MJJGvlELa/EVYO/FmrmTRTeYy8Chcak/X/gvjQSKkYScbnqzCyiszRENf
sNkntAqxBN+Hto6OP/3fToRI3VDHcgpKBQqHKwqGLj0KaTLue8IStnQvIZdngX2cPK7EkxbjpT1T
y1WjXKkqK/D03x+SvdYkoB6tlngR1t0+UeB3l9Df3IgDGo2rqyaYnT1jun1skRlEATCxHjnP4zUD
WgrvEF9yK8M75p0V4izNEk1JENFrYSgBHi2MHY/KUQuTxddizRz6lajeRdc5VMmMt3eJsnrR4cj/
cpcnB4SENBIFbNn6sKid7wPub7JHv0rxNtx7TNZwE5svnuko5I6D1lcidf1k40YZ9aW4+3IHHZzq
malcWKU/3aZa/uS9g95D3ZdYU+S2U1qXdwsqIhI0+6r/zHwtDGsdgebytGdezwsySgI7DHT2r7Ki
3ZOrSuAO69jnFQZkIZx16EgXSW/uVvpRL+h54Lomg0EekcHKJdeTQDAv3gIb5N8m9wuuPYXSi4WT
yV0Tc7P5JafQDprhyPiJC2qxU9ACkB0BMl/Lju+PGnoxZghR8wkWLYtZv6Nj0uQKl3itgXG1jpRJ
5B3z0cKH4nwdvwH19ZwoahMIh37DXYyzDq9bubcHNycXkD1e21/8zl+ubEJdXZQ8FcbF6MMuh2OL
EzvtZUpfiqhbWxpv5K5cpdI+jGp93jWdnMiX8dSW2/jVyGq1xntYct61M+E8GlpNu9/lMumnQMit
1Iw0KQzlXIcrM8U1j7ZNKbTh9YrDvHXM6b4zNQYHKwVdS1ptyzp5cHT5umT1peUmSPo1FeznfWL6
+Uw+H38QrQPRpSAKGVnamnpQNJ0B4bKBv94ROv4fd3/S3Lg6X4BtyjVPfR/ljKF1gSHFaAJefKPy
/l4Sn8p0ZXeW5gJXotZ7DMBuPFGcVEwcaen7tirsXpjRlcML/PDiuYo2Mc2gN5vdnvecpy6b8odh
U0TenaTB8oCS0wsiUWOR1dncWObt2tFuJU7tIRPBoiRAUrFoaZWv7BltlG6c0XvCNfrU8pP1CjIZ
yQq3d/k0FlNOM9tb76Ua6wmvwZTFwP7xlVPG0YF60MfIGHtiUz9d48QQgKmR6GNdpOCsdypykwkO
2sE07eQ5lEMXWmaiIOZhbl/s2OXxOwKDhNviL2K7poVNHEPwUokPa0tC966i6hNicI8LJmwz5zcM
NtFimIhQPkAWHClabpqKTXOGENIAh7wyLWPC0SCpsKr1XW8WnmeqBbvDGAlnXRjK7vHD24Ra4nNZ
VBCUgvbyubgx8iuk09LkYhneYe0rHy+uULF1Zcsplg27QxQ3rGqO+VNixOnITc25dgsu/PXd50lT
0ZBBQTMToK3qM1RlG27b7YZ4bvzICM/3ol8ir5XGh+clGMdJBSErfKaAb30cVyYgck2O2dinctzX
tbkGdK1tXULdHBKMlrjiFUREjTDue03RJXY75YD5IbSiyPlJ2hGAgudvyoAptytLwEhSDMt3tVmT
+7AP7jVa1aKUXtfhFl/CN7KhMkMHFoJ9HdLNWzdqeUHAJQ+tl4jM1p7yOGpEXDSSBQB/g3HIe+lR
WpVB5xN1QKp5TzEimxsG/AGWE6i3c4IXyzJMxsCz+HZG+e/J/KLijk0H9jt1lSgYAUPLHfQk9zPK
SVDItu6kiVJELIeoIPmMG+ZrY5qvRweNKVEJH1IYhRrMqAtvYLSu8/awRx20rzY6CE9sW4YLECmf
mz0TUtE7DVPjS9hQOyuSMFSUuevk15/kSZLWNVSEBw9buSTL53uq0792fxOb4J0VPhZiKuHVW8g3
fSU8/x3wgH5X1qqEAVo2gsVcFryJUKPs/yZHB55kkJzQ8qeFmRAmYXx3XFbKhObp2Kv/xF/k20aV
BLrZ2imkyBAMI2QXByjy2JXnDO7MGPBeah6dvHEJVj7ZF5n0D+Yk8TrUplNrJrkWnlLNMj5GPdQi
Ids2XJxet1NXHT1qdapov82lGJAA3mZGBk8uDVC7qVnzxGcIB74cZEODcO89PPNhc9ip2x2Yg9eJ
OWys3fOtjvW5xyl1pdI9pKcQL4hBNjyOfb0Kn/zwqMheSWKvNR0g3qHTWDrB+Gfc7fmq9DIre7vA
QelXtL8Vr7v4E2R72LxVi0tFL0QP2y0wEGiFlGOJiuU1HOepD/BSdmVRpktrdqrkRN6geUGK0B3s
CQr34k3d2dWbZMd3Ea1RnQq6Lhd9z7CaTJsTlxVqdeCkjZhxZYvHuP/ma/jn1uwudOyozCU/RW/j
BN0pfjdNkeqDg2gjmnWNwTcIU/cUlI0/6RQAuSCO7cUdK+V0KndkzIOeiT8l/6CtShKhhcUA83Xh
3AXRA8c41GTeHyUwOWaRqwBhhw/oPB/xYkSrPInyepS2o40Yy9Ca5rStGxj1NeFDL8ULS5coZXva
E/UAO+Rx2W/LQczutZAQ9uhMXrXuyVedAbN87WA69nINXtxLOXTOy11nXAjMSgmSNngUxzKDLmvM
PPhfaoG/8y1ZSa3JOGBDEIwntZtrcBAk7SZcfb+J4/hK5nxu/HYRY38FW1vXtI9qYHWJCDOrBGUU
G36iymA79d/AvKq0uvzpCDLHv0d6pNCUtLILTNFCpe1SokYnRK9yFAOYI8rZ1vehpGngFafEHSd+
IefRpvtFYyg6ii2OYL4VTgqEQ5sjlqWHkSWG2uJga1VH+nhQk24MolvTqvlHhHw0Vf97wc4XcU/O
KVSOKJ/Ry19spFZ0Xlz76NsEFh4ynIMiAX10WETAXEbjB82pYH8n0NpyWG9RJ5gugGIOC7yx1TQ1
4VlhMcziwSMg/eki95FZEVD2NNYCl0i0Hh/jyGDvFQARYkpvfg6SysdaAfGEXGgAUt3caNqnvRJF
FNYRVpE8a4pjm2oExESrQWmPdp/K2muwm0ooXAFVhtJ0k2rMIwtKEc65gRRx1kXmqVjbRRPWkDg9
rm+EJlFcksw1AzuxoMqbu2onilAAvECazTt//TONCQqzJt70KsBKuz62EQ7/L0Wf0w1h0Z3bgzMG
Bck88/sxqtSxGy/moFP6gRAh3xDbPudzSedU9MO0DacguOq+IVEUq5Tm2b0DdrpcpO7XNuxuUEDw
bI9/EfpB75GSOt7RexkRtApH8fvmry4FwpaunS5EDS4Mn/Zmj3bCjsbuMzzfFIE7dfrfq+8Fa82G
rOZHc4zlzYF7vNwuSewwChmb9V6QMdJ2+sIcjmsx0lGuHSFDSXllZaF7Lu6Y3o+TCa34e84e+wLH
galZiXISN6xFi89f40ppLwCiRuw2Jhq47Fw67FtO4AGLLVWc+JFtqztItY5T6ccSW5GtVNeNbetJ
ZOTWTGLUeBlW/TGHULtf5CegHujabj8px3gaJpd5tf37Kvr0fZUiVkUnRH4eqZhQJWsWZ6N+YYT8
77lsCQkrWDwzfxscn0K/GXw45z/vKp4VSfczJD8LvK4U5xC4Czpr+lxZ2XqbVbs+V0/gPZwNijuK
r2c6xoDqYQsoKbheagZOcwf3jsKrTFTJ0Llguwrnn+IPuYtbRVwF7hi21is/0TdE8PREgXFgHCpz
80LVMm+DIO7wO7wkqliWwmof2KcHVOkl4UFy1J4gPvEvpUwYex5Vmw2r7FrzjLnVe6ke/gxMU73o
zNkuut+cPwPcU94dhk5ELsMnmiclRwHr0jxNnb+MrJV2YM6yaOWNUQ5Y3ftu3QGULlM5Z9Rj5y2Y
UUUoWjVSg+IiSIBNGOd3l83e2/+mrIx6zCrazxMrsxOuPcSeSDH5/YxeA6ZEEGzpAfmUAmsRbbTF
zCrvbHvfiDZ6bZDZSVhqfHofVWBJtZK517Zv330wgMCQd4/rqBxdPJiujDrrWcY5w7eJJHUMWrbf
iUVc1rngwUQhozhMqXes6VghBb8SDvgB3Sar6PNRrH6nM60jd3xPmHA/OQIipgpwBEehiXPL/l8U
YOGulv0k4ad7nlBLo20o04+51XfJqe3fMFuPLxAa9hm5c9jJIERKfejF/4mmhyUyI2ybjCIvMHr1
ZssmZ/HoDL9+R7OOovxj8A1Be6T2tvD8B1xW++HDvbBkgyevM0vbPv3DZm39F/z8x9C73cbgeNL2
USmUEu1imeVh/rGPxXCAuDlOKMnVKMi/YyG2OGJWUdJb6ZJg/lyNr0noYbO92zdVfbpTEWBji3oa
H7CO4pd4okMRXQwNxNr5HyDjccrKbJLvRYEB5vJMLEgvpt3H+CKP1kyfgBa/iH3UzaT9f8Z3Q+Ye
Z9FUbAvucYbsqftGDvoMLjHPtdQ6ND/GbgtvjZw1DaJWH7eRVj8vP8D3lhufeVwQ+bxSMLheCShT
Y7x5gtGB/ZpNvkUw4b9zNWXDHuSQRm2NJOHMAO8Ek1S34FdSob2N+NksF7X/6BbU6WpsXzLXlYdc
CGsiv2ZKgHRO01XCPmQsyyu6D2GliAzCkTXpY28HmGbUQ2PuF8xMC4gBEW55+xQeIwxGEt4jXOLf
x+XppTextgzyIpIdRCMiGpe8JUfjrWPnBr4JWkmZl71XsvE8/TFZwMRUN68pD5j8IMminVZ3N366
Dvhgp/8GIaQjuJWnOmxrA4dGsCCYCsbZxYwgSS3YK1T/m8PtCWEdi0WzoJdHTP8IJ0T749S9yswi
3GEoidw5GebgWjfj8ENwvyC5p7u2vOLJMUdOvMHINbMXBYBu3HhwFW6MSnCgEmaNB1aFgGqWBZFt
sQlY7Sg478rInqmlRLtvl7019OI5QmejvvQFtv7TAsa0EpDO7zRdX6ubZMD94Bn2qbaWnERQF3IR
dUfjOPRU7za1jE8OhUz4BVVsuTloa069O5iBQGFZ30os/hcadV6vAcoOGlWhBqXvNRkygRSL/m3V
Vu+VMjGCV2MHz3KOg+NfRQGswTG4qMZkhjpA1hXpWKP0Kl//UknI2TwoWv8c7rhWE01lGm2N4x/k
ecYdLfMDq/pOpdZxMAf2b2un9aJI04gKigsuUFfop9Ndg0E+e0AL7L6vm4rgsnqzMe8gxx1YQRAy
Dlt9UOFM8/9LCN+tqXN80H/CHzWStOnwWPUttj1X0pt8yis7kJk+rRyIaKlweX6YG/MNWMulht0H
AfR8JKGMy3fGKiYv1OyT5rXWWGvs7RbvS7q7OZvRwZaDLqXqvPh6pJjt8kDV53lvOzxnoXvOmnhu
TpMaHoLIPz9bLEatmmnP8n/kvkMHUpg5rM3Do/4/rtQxt4YI2IlZp9+k+CVMRWkFrJOhDjIH/U/W
gW5Nu84GDujyysAG/7vhksHikCyUmWxAwpedDTie8r54P5VesbIlV1OWhC6vpxTD5tbV2XDF81nX
fS3zAYj9RZjliPyYfjl7f0mQd5Pf3ZElsWopof1DiBd2ScJnaG0ZI/C4VsUHz2GBlPR+RAStbSHd
MqGRWX8mj6fOsyh83LaYiXbNFt+FdJlMCaV+rHmLMCWM6YLgtqIi0FhozjUK4UpBlwRU3GEYIjtV
MqxKv9umG7o9npFhaeMynI/BtnPv1vdDWQwSqBKbzdLkl1UkNJuPG5xT/LYPherWKgmGA91xxKoB
ysVCocoEPBVQsuRTkj2rG6ksvPB/rSClHkky5abseDiit9gzuE8wFDbrmhSk6tzclUTX/3OXvVuT
4+xX0hpX5k38hvwNJuQ1Lq0Y+hM39rylGx2FU7cD6jfHjbu8nwDWuv5m8pQcGCqRqBi2zddZB1nv
DHsm+nWaw2NVgZRj9jukWOx+05N1KElDTiAGt0PJfYVC71Pnt2Hg99W9dn8S3CXHfnhnuXc34q8Z
Gj17jsDCXmZV9IEgcOPUup18jY5n/KgKcC0qfqpxMAGp1mKjnpQx2hKi5aGETTGk6G7MYR4hEFjn
oOKbTYlYPiMpeNNhNSe85/AfF4c82B2tR8Oui1njMF0s8uJnTRUe+CaaBdvOxu9ianfB9qzNVSkS
+/+xTF97PbMqGko5C8+I5hA/sZO1hLPaR0TxECY20Q8fefV2t856IfxJgYk2c+xFN07qYhzwEgXl
plzMoh+eLK7bquErcBb5oVM0WEeRKIq3EWEaPfRXwqIf7n6L1gjNmiwB2maSlDAA6KxYYGT0BrRc
ajBaE+e653FV2mqIXE+kyJ79M1T1u90/WWqHosvCwhbdobuCvXlU2tEnMTcvAP2VhL6z6Q1YGS1A
ExSFBkxbHtgUKEXMS+hmj7Jm9l5bejy6ZtfMYvG1l+Qt1dg5QDOpN5r5cjgPeuw18ndWFKrqpiLL
chMxaFe6Mw1od5Hx3rkkk1Ouqv99p1m51WtpegYgheNZHls8FFaKnpmJB2RazNOkztO+4gHF6Nj0
PJTbCmSWO5mV8FJQDM6HAsnn1ahEsIUhQPGI9DqxuUR0yq9vkWzdOpDJN6b6lYeBf5kZz2V83WDS
EPs/RFmD/ewnHja95y2fRHo82j0X+bxHyvCYBXnOiYuHjkHiMvVTXU1uVTtjzVbj+vjStMzN+6v1
VADIshGETMhZ5WaVekAq0sfgTc7wCcwimivDl18irwz/9lHsG4crZgmmCB5aWkaFUIWcQ28U7f6k
9t0iGt/OSs2KyUcVDxrnSglRWfAluAMRop/FKFDMGXHYJVloL5Zh3V/h4OSf6R/PU3VH3IAoNQe/
/iasigl9YgFWViBbdbhk2Fqi0iK5ZJa9y2sKIFMGnoaJQvPdO+gMkjWav9Cl5E4R0Ztn5OuzN3vU
lbPd5VFL6naoBIsR9u/gbaefKzXtvw69YCciDM0zY3+C+eZg8H0c8OsjlMITO42PzD9IFM7p+b3F
tPBDoDmwgjmv5TapvwrKn3AORmr++JlTrJcUV2VTS9wXUIFjfrT9DILCaPJpW+rn8ffJXekCUnk7
6mVbhHUXF4XlIzgRruWv+gvmx+XRopfqEdC7DxwEgyDNdyL2wSrQn6ZYriHMeS6eFdg02Ss3hB21
g6HRk9olsnhhhHsfxb5ShzVELj2nRXePHMeG2m6BmzYsFnrfyjEMJYMq3EDqukZDhKhBHJpbVru9
j+E2z3ODfUq8ruhrBjPJTFAqJQ4UzDbGonI0jzOXDi2NRJK/EbABeI+PhSEXwzpK/V7B/WkRtYpk
2rs/4zQNtADc2m3XbS+uBxce9xJ41MeOvs4MEWoxtsWtZOJOAioeIwx1BXA/4T1j+F0B9oVl9swd
Ecn8ZtReAXy5gbg5oodqlKODGOktfxYgOv89yk7HUS5bOETiaoKFwyQiNRIP51OwynOy1HxxAJvv
GY7/zWQnL/5hEdsoTOCvpwI+fGz8N4uhT104egaGxm8VNTwcNgtr+QtGRlR9e/ZXlBHgg1DJulgR
tLofmwz9nTcK71HEqK9dMJvHXO/Gh3bM5Z1006hl9sUgS/dSdf0pWwpgM8M8Fni3eW+d2dUQmcgu
Cg62SHEd7szCHjqszRbnHzGb93M904usWahUP2hivWivG02vfJaDsJesjauCj+oZZW2o8Cw55DCE
u1OuWfNLB8wYUAAbjS+qvrZS8vBF8BEGUBJW9b8yCzteZ/ldkXFq1Ql+K+2xhbsvxAQWJ5PSQpwt
kLSOtj/oeGCbNpoEN1Fj+fMPaLgIudgr+ZfyV3G87SUUtu05I+T8yPs/1tbQGqX8qqIqPTc1UKO3
7AjSXL6sTyDRkdIv5h0fpIim5cGl8N6PsAhvhMu8cYpYuAhlbzwSXYzqn988Eeqxv3/nxulLy6Tg
48HIXXqrBNiS3h+MPkvktm/WE/84j/3/bQ8Y6iyaRa6NHqiTIHVXCj8yJtvcEOw90r0C1yl4MKvS
nUMlWPe6i6rHLi4zvxPBc8heCfZvVr6prbLpnC7Ru3ufpdPA8H1MJShaulaEEYsOsCQX847pyO2x
JlbY2QP8IppyKXlLXun1DegPIimm5qdHB6FW9ymgoWsbWA+VVBnkiOAGE17oddM7+WPHUQl7AA88
QGm2mcw/WwZt2kJVJ8BSWZc2GDByWU7wYEZJ2HwHDlWBJUPNdN6DqcS1PtY3CRJozy8xYjh4B9Wo
VTeOOE65TlXUfkAc0s9aTWhPRz93hcb2X3noz2sxVbetcgVhINCieHgBb7WtBxTBgu+NzDMKr1qP
Rk6bC40Ql5/r5rAIwUtgLZlBNLmuzQVR3vf5bvvkj6+O5pgT+zCwZCKfAzp5VJQ66nxxdHrmq7B7
1g/EkMLVbZP/cu+AX0B0MzCp3JJpNzmsTMPExtptl7ZzNMANef8sREQjH6sgybcMQOVv5vmqVs9h
qKDu5FbNKV5Pf/g14kHe8DvwSwQlgBOtdEkTxWYutWaG3L9JiGT5NdqTJHzCqAyxilBwJB8Ab7rl
3G1dYuNaemU1Qe3NPfrU1TRHBhjoz3xVSAjaUwQFrR53E929D+rQU4ETP0mpPa+znUMNlfSHWKYz
L/KUULiUFUhy1z0OfiSHtXFH1kthQAw4AFncP2/j5QYNpuunJIo7LeDjGEu9h9hEAzpd1f3vc/aX
It3KnfPHnOxFDCV0Z18YNZFmezDby1NRPHeY3YtrSxbc/hqN7Ri6KBrfqitwE6iYpxeAL2OuSdxW
ThfakPVrI01fHaZsHX5n82/GyPiiu5kkFlRVs8+MCpH7dujNf7acp63MgwWXfQlhFjr31ABK+B7n
kpgq0XkP59x9WXnmQwt5gCh7qgWaV5sCSCvDV2hh4FUhxIl0++VfG1Wvkp9IUbZgB/f0bHlcNwE5
idBZAsq67vrtBcVFYxqS9r5JShdp4IhLWQOjTcQfrQ/PQopKkGE3Kiwwb+rmb7AmsKtUZoUnpWEJ
nyTob7UTvwxllMx6js9vd7Knr5QW/wmj6llZFj7dcTuRWfHKT5osO8BrXT5vSAFwpgFvFFrbG6oU
ha/IrE19iFaEGsjZ/l0+/BJisobHk2Rz18UrGEpMQgqYwJzSt3YNj/6GlL+EU0SQ6J1b0yMzqMhk
Ki+HUEblC4c1kHpXznOzDWPw6lWpowAB+rVw7M+eTjuuhNxcLA1TOHpYG7/M+vGl6ZIg81flaCbs
Ok/GE/yRx6m9Zkrx05XQIFZg5H0RQ91iZBlPiSYC2+0fEtx76VMOx4Jhq637OcYwTXa3EfBtHLfv
Ov5Pwe/h/BBS8t4o+i5GTVgwOmxOPzp5x0zyikXGoPIb+qjVCUOSGMHqIhq7frHrnY78bKzwkrkl
FwY1RlFd7U0szgkFHTvjlp/2D7Zc6AMq1br5q+vfljvfpZRFr5pkFF1ltwgj64AD+w89zzBrInoK
ErX30GRM/5bQLqkVPOKs/IN3odSUYWE3LnSA2EFXuoOUmGz5rK9WoVVZAeJHHt0nRS/94GojO6Zz
Dxs6iybKoIlxfFypwduhegIf+KOoquAj69CTtoj2pnU3C/FFlOTOUCb6j0DveBtOLevYtpw6km/W
lqYdOgObl3d6+et1O1WiEMnbyTsHQ8oBUipKSjr64vSNkQkKuqmPkOSlmIaUO0vFT9PA5DtqPlbX
1359inrLLDyW85QT4UCEILtSGZ4U/TSHL43EsT2d+M8yrqdd4uuNiRBd8BUWvrsJTghGmu8DYaxD
ODrMWpL9sHCdBBLX9Jj8pEAdqvJFMcwKVr1ltd1ZtRieFuZItvmrzpGeQkKtP05CKwbLgIU3xSkv
Xv3jK3+b8FbNj7W2W5hNGMl7K3mSQ/0az/9fwXqksKcuAqxjK96xvZGCrViCsbT9YW6SAay3/lOT
eStfuejkqv1jSXCz3il2jLwNFSh6FkYe6THBn3DIE/aJuSjOeXv5MzYk030lZ902KTrgVI7kr0cT
vA4N5OMBGW70gZ6eK7wHlRr3YKscXEWGY1zAcJZmB5uGKXFA2zKkR9F+VXWkcfElK7uBilg15GxR
rnIODoGgJSeqJaJ6unL0tK/Z/qsjfDipbzkb/x9ABonXMB7hJPjTidUiRxUB+Zkmml1Wt9nu2/xG
7X5MGLVGYGB/ix8DgAUr4qXYGoPJmTUIaRsri0iq6L/UPSD2zGBZOH/4fD53zcdWusr1fsw3wwdX
sihec1oRJIpQ4LoAlYvl44KIjd1+otTQeZdg75fO+0NYbwZh9EOXJjan7XYxD8LHkCRgGk2/jaC6
vmEwdYK8a6dpo9iwVf8naw7sgmTIKn46ERwy/aoRWKZop/L0tyRsCg2r16iJkqm8rPXLg7CWlos2
Va/yVDYjHalgA28kgzEThtqNG+XooeO0waCA34KVvy3b7R6e9iV21eoNFj+E+9Uc4HpoqhSu/Fn2
QzTZF2EeEGsZJ+KQooY6lq6GLzH15pjkPVROvjzGEZ0jLXO1rooBlwN7dQSLgVh+alR5rqguYeSp
a/1XQH0vRCrfF3blcbTwwx9X08y3PAQEC0//tvtf45ipH028e37uIsOHH6fr3qrUULtOVDGlYx5f
55rVcUN9febPy++iw7+819fxElyZ0p1JR0R2EsEB/QOd3ed67v4JPSld6CkqZnOcPQQpRA2t1qI3
f79QKcx7GVXx4UnR7HKt8lCsAGjlpGHMfNeFdYTl+lyT1vEPxZ+AoEaMkLN0DY97zyyeYBOPjRkX
MDMLADU3gGY0BNOWblPfQe3/BIrwIS4atNVFax+5UZXQ3L7nMDutFDQl6DUsPJ+fEM8FItdFLqC9
+dmqak+Z/P7tBgTLFRow04UdtoBfZc++S11K78w+/B6m0mzEhUkGideHLs/0JgW46Z5ezAee140U
PbhecKNEMqSM8T5h+jmXT70x2vjJLrDWUWCDVV3a6jcm4YbPM7HG6ooxOiD/FUgULze4JbuB3JgP
KfDugW7Gqlr4Gh+JfjBpCCWL9Ll9Pmw3F4016M2JuIbY/AQI6WsomAyWRdQ/Nr/sXYHpAsL1TFxP
UQoqgFmtayZKPC2O8Tk1KWd729CYi8dHKpZ0jfcAa5biiY79w88anEG4mmH/iTtgiU1gw+TC9QGS
xKf30pmLfhPAOMQtu+ZfN6dmcobEA43zbXpOk2gh26hYcSyU7owdca9Pn9UQ64lktyA0lYRCUN2q
80lMlVP5RxM4KFgpod+Rcl9fqrZP60I9F7vWotvEb4nZwbLiGObFQ8DpIcLupGNg9KTynZGglN8F
5mUocXUCsfbKrchJ1/653kVJH40tK62nX/ICi4HqD0vrZLWlKGAFTxmhNdxI5kMD8iuC5WmED/b0
fxRQQTfiOaNwZxkE48m3AbngTnYudtwr51ql03OoLcRBH9oR7nCtm76aU5geltL0DVrgfidhP4kP
nY3EFc542nVPbEpRHbfwbDkGAbMpZtNk/OJv4j/dmwBDD8WBmkYzv4JwmKHTh6kQg8QXSBejTjTu
FO1vN+b+pTggOC2UVkUKeBSs5atppAtc9r2xbXT+zaP5UhI4olRJ1iPiHkzV4fWrMqQ3uzG3LL9D
QbLEZjPyu7ywKqL/bX7IDXlb8Sh4/tOJGZL0r4LileGBktVPRUvQ+VGQlsMB4Hy2ywGPL6jiOvJu
gfygnG5mEnyHfSV4qACl7fnUJqZFd1TN0DAST0mVDvgWa6iu2Y7w18tQLt5z+RLUSDY0qb0mEG1a
I+O+GCFUtorC/uB+4VNjpT3rkqZjx5aE6n6X4hjRziJiMX/37v/RlfpHJphvwv9WhLp7Sl9pfq0l
PXY5ApO6SOSu9oUn9Gmxpo5YcTW1HdvqK1iDiVI8s8xVkQAoBYhDJexXnE2Eb9hGabevY/+kazqx
p9Fw7sOvdHcxo+NZloy8FSe3Z0Yc676bcQ6GwfI6WofI5jyGoLM4sNxrCUJopV9IM1ebC3qCf/4n
wOALx7Qsrc3e64FcqxudYUNUlf8QjTx+F7bcK5muL3KgfIfkRo+dkBn+K1NkPVMZNydN2hPC18xm
zUT9KOcMC1D6OeIAr/4GFUxTraLhZMjwgSUVtSv9vRTOKBYlG8GRZwOzEfF+9uPlDa86jkLuHkV8
qMMCtxoq7vSjZGeJspS4IqavQe0nfZ1sEgA3hdh5a2qhWqNUmCvWqy6dK9ZJb1q8btStrXUzSQHx
BBGpnrwkmTlNkHnqFdnVJ272W5iHp5A6TEPbUMEEbxdT7HY8bKVQHgGEJ91zJ7q2xDeD2fa87tD3
8Pb55c7qwuESlb12B7f7qy3lZpNHKNh++md8NbVEdrqHgC/oo7fk/9hFKOmBPs1bML1+pOMRiHAJ
2/CFB4QC+8TzWEBE3z3WrH094C/B4eC2hJeZ/R76Q5EkzkZh2DTnnctk202jDK2rOHHHG7hC63uJ
+i4DbL5yGjcQUR6crYEC81aAXSlrEI84u/TPJ0ovUvbgGqPLef5hXQrQSeksF937P8PQWIjq3zr0
MGp/jRRZlqceKLodpeAH0gtqzVUa6ZosiYWLL+p8KjG9Q5SUNYkrkwDT+iV29TMHu3Qs7KRPKn2S
/aKmjax4pK0w0DMMPwXUT67+Bb3IzBsMcjO2g2tqZHvOJKJrdilrfL3/qLhAaYD0KLGCqu1QXEBS
5zHrgURv1XL5jK3VJagG7tJ8+edWnAmISD5iwmM61siIvVPwdLacidKRtgWy1HQGGIl0O6VaCqFW
fPGW+t7ze9hmmOacdD+rmWq6b8nRk4WHCCxDd7Tefe0e3IZB9XIWDIIM7pvy8aLPeUnt7I5GQq2U
fX70qLrtHR6UiQeTqjCNtaqH9v0CfLBENHnJJFh5vCtbFF1JHt4PWQz7tDkTZ0z5t5zxSiPVTOMi
Pg8DwsKyu8NrNfmMek9mJyc177uCCcHlST7vg+dYcrUQRkOj17cUAzQDcA6EbrT5gxWMBkQxZ9Wf
ufdi9IqlLroGamiMeIVhJyhaLLETDr5zsANaGp3YuZnODesiWqMTxDFjTPyrZGs/RX9H0M/DuzfT
ZMOcjHOp8q2EsYMGSiKRogcxYsvRjkAdz9ezO+iR+OJhfT8vSQLiIkY3Mo9rOvZWhTLfgAz9HY7f
J18RrYqck39i7McHq2MrHs7Nbma4zbagYY64DfeyNcMZ12RNBVuO/mgtQD2aZDA78fEOMBRyCH1l
g+OH0aAdUnuC4N4QY3lI5lu+6CzHBT1vyDkLGGv0xAGA6sVci8cw0md9qFwNfIqSLKS6oGCofhmn
Du3+AGFRJADwj3QMojWf14C2XCeLG8VPIgFEZLs269saNUPMOwYZC2XxuOumXU5a2y0xhEorbOOf
rHyHU4zPRqt0H7u9ezRS26TieiubvhRswfZpcRxUZyfwQvg1WvOlFF8bKmUJ1iU5zdv+lpNr7QYe
KCLLDZB0GgjVIXgQCq5Y1O1TNklGrowoua8pxMatEZV8h7yFQuBqT3xGOBSD+i2u6HPig1rw9QHQ
aOW1YUtZ8F290ECg3P/MywCBwFo7cnYAPNSYuUQR80H8p3b17GC6cjiL4kP4EFziy0i+OG8GnA2Z
+tGXqDR726ecxb1hijp2nlN5WbXBA4Br5gLIQNk5JoUANYyI0TFKajUN8anL0YJDkXQPyeP7JO7Z
c+JhQrh/ookbm3QPXmIK896VS31NnUvmPl6KYtYMy9nA4Nd6nnerXHgkpizHTZgkCZ5ToOuzzb5O
jZsYLaU9mtVvKKaeJZ7YO6tsiGsGfDGcfj5Hkfzw3lbZ5L0+A/sf1APCLpmwtjL4qhlNfR1kwK4h
Zx4lRQ0TqDWr7QMyLeNTXWdmugScgks0bjhX8rp4FWYBjXmhJFaf08kQHkW1OFQve0D8wukxlEWu
kW5N3V8lN9DMReJDhR/pgYpsj8HrcPRD6EVK0OeLjqv3kVRHuEr4QDCcFVtzTgqVfnbpeiTAVNla
5SxFSlQSewY1krLnnInkP6BcoSiK4+O6toFPxGIQOkqeagHr2QCc133ATKpHYGh8Cj/7ZgmkPQ1q
VMYQCFTzyZRyhA50mD/wRLm8vsTBeuLlmg2BIsFlb5mCCY1K46nu4/nIWDoUxnPOrSCna0H3Oyvf
+9W/D0up/RdjfcCa3iceO6N1ZWua5uWuIbmwtxL8p81FaUqRJ7MrhmNwHnhCOYhT9YS3vyhFRWdo
Ht0Hq0b2flppUyAv2wpVgyO7Pn2n6tOdUjw7i7NXXVfgE7PnhumF3d8jbT0any/wfSsWvGWutysy
zRNa3v2PthUiey8Gs73n+Oww7VWqe2cl5PFnHXb9TpI86jDJlBiBJwzU0clHYxn2tOpkwOoiDFuV
WvVhYTGDK79CKEXVxgpC+Uxhe+P0cwcHr0z+/qrtGcGE1+qhhoC2QO/tkLpic2yZj33ExzZeaeLm
2pem0D22P4Nzj4Mb+9oGqQxa0jifMN7IMa+qdLV5PuSfpV7QzWfLOClGon22vtWXt+Ym2SKQBtd5
GlfLEZHwRhVeP2RDCG89M36MCinjBJvwb7E9xXNiBmQdJ+nZWI5R3tIEOV5+mjGcOIPDw4W5qIjl
Ee76pE979I4j5vJadDPT1N7tCOA4FnDoNUFUpi8MFq5j+O9UlHZENo2XRWh4SIAqoauMlJtFe6dB
Z8l1m/aUpjr+//yxGM4dTUCYOcwPGG4U+r+lziVQzKXp+cmfJXR1nsRrR5Lf5t8tSNgQfb/aF+86
hlbXzih2PFujf4g9DBvpS0pUufACCq6q/L7iUZyKBJ1UYTMJ5XGwHiJei+22JCa34MdcfbC1DSa1
fhABDCiqKNia2fnCsfoB1ch4etH9SVes/QhaZ4HzrDmE44kvDz6ChfySLUnF5jzUZSoxw25k+L5I
p70eIRYP14S0S/CtJJqPSEURen3WEvqyJqLeXw/gFYhvqou+U1bDZjpDG2gj5MY9W2OS4MYfIjra
WuSCFPYo8+BwliTtmPgxst2YearOn75K3h17dNItsDKa4fmdvRQB4jpladikxQ3+nt1QKYG9U6LM
HSs6JO8yeFmCSKtEzyZaiCebFd+PCF0pfo9WURqHlHT6pf+A/uWjsDuDPyxilRB3jm6OCy+kG1ef
N1UxZWj4f9PJwSvd5wq3QTBHSfbVM5HUqdsNITlBfZkcHejcMgPRnehzgAKnSlrGzKrcXNn2Q0vr
kSCs2ALY7liprjTxXxYa92y/CRVcMpvEXnpaotNHhSDvIqbZeYldDXObmzgLNXTiULVcVp1avei9
ftHy5idj0hSVHayJbSCRTMvdQmsgBW11Idl6OrxjqYFCcn0WGFup04yqtgMzVPXhdHxZkNPYGWSR
S359zPbiQ1KX1zwW3Oh6F+OI6B1eIGWBDGYNqyxVeqY33AVvdAvHicCpfBXVET7F9aDBsQUSMLYH
ijaPTdnouo5sH+VmrAC5HPyZ3NLU7ePLQfbM5D5IKnh36N/gtCrQ1dybAftTgqicCZuEfPh9pr+Z
YxnP4DZ5d9KGbVTNrPw7oQ1Wi6yFmqhT9Z819DmdNrMShbag77rSdB2PgmW42d9FB+yb763UBkPc
p+ssRT74gj3RQjwJ/BDOZVlXI7+WNGp3CkV7jpInpniyYhhUTDnS2whIGyZ72xUGowuNs1VAXyEi
PGdm97Ry/BSaMrRCs6ClUexRJgN+Hu0PYdfCntK1GydwnX/WuSdLRDBWSLbJSac/hYj1xCWOb/tX
4JLFlGNFE5fhckWhanvSX/DZ2A0OAciLfh3CYnSOWvHffXtkGzgSrXQ4HjfBECfjBNLQIX9r3uPq
OU/f8poo+Y8ujmsKqHWQc1TUZzFJBDMINjjBdmm0fnfQqtqQBUS2ykqrMmwdK/0pqksIj9BNWnE/
V4g1JiK5mQapuUm765E7za4gIVegGKne99xrdF5a6srNr7V7ufgeTwpU8Ud/NhHB765EpympST8P
Aa+EDqsZ+eFPMGhEteXJS8U85pTjQX1/MEH2Fm9XY1EKwlmr47BBRc+yT7NUEOiEL+OXeAQyOCTA
f8071WVvfX/nJfpXcyxnfIdx9ehnj1JW6nVK1LLBgE7WP883AEoRMC/NpwZwos1ooXA18nJqOyNO
IvHKoCAD5K3PXxCnZdZXL4mYpzb7yrJoqczO+NRtDB8m3YgW5wsi3OGzWYnUEb5TuPQdPFpeRCZW
1msfYAM2zIG95WOahi0Ukq1El8AhXbNXqKv/9YFibIuIAC+AAAtvZ/wNoq9PW++6qQS+CCt/S3Eq
MrH+fKwQlZ74ee3KnzD541a3bWWGM3igX26ziq07gx3u0TWI+nEEEXbUMu1ZINr+wybrstGxizlw
FA05FN76MWtBW/MwdaCCsFEKBeu8doWs/eTfMX/w4deY3De4CmRGozmX1jixvucTT51PuWfbjMZX
nK12PzfXpIU/mw3r4+lx7Sm/UWbI6mMxOCz6zgMcy2bM9GDl6CJW6fzXkVQZpKB8y055MWtfmdd5
4hcltmR9g2o74DrElKGIObuDXZ8Dwgr7PjYnIAstWVQbI4E8u3ZK1/LQm4vD8i2HK7MtM8GrDjg4
oBsL+3c3zWPyW5l/NipvQE0w6Dx5H+XVjQe5wJB7EkzT/3kSreLKLj76utHnTGJsTiXzVvE5a+Eo
pCsI1wVh/EwXQEBpScyPup5YEnhLcra+ptKHj1/CgXb5ooUCo9ZB1vljF+F2L5APDHHKdq3A8ArK
el1jtQSOh+GN+EEJL67F8KVjjJwUZkyAA7QzJz/VhLcG/rZmLzaaDvfWha2t4HFDXj+fEFZkWwUU
KQTMXVvpdv6BwZmT6Auy1GsMaz1ny5dSOK3EE+RimnqXn8mkHlI4gQkcVMSXMx3fdgz5IUnYoV0s
iz1XuWrRJK0Pty3CdaP8a3owo6fsTIZYZCIszMGz8BVOnN77bn8tBqxCfii8xH+qsqF0CxkXEQOm
cKTP2HFsJWQpKepZbenWwBhd9w6WBVwubgy4z61idhWhvC0qhlyn7XKCOWd6LzAYBqz6WxWj4hwL
PsxUSGYW51yV1wVebtjPGtDQSZYntTkoXwSfBve8WiKtD4utaM+hloB5afQjYF1ufbPXt5me0gj0
H7DDwbLK5BYlO7IlqVD514zHpc3C/raBiAG3ShnwvgfCcA1xxHlzzxbmPS+70fd8xT+fW3yaP2T/
M0HLKRVu0e6SkO1+TUTYG/MAKAHO9jcLaHOcYmM7CEMwE04nYw1gqMf6F+RENiO+eT5ZWnQaRZVt
J0il55TulgqcObo++jgvStfeIxEBTK4M3rG61g/YZOZ7Uuu7ANQgw94q5nqR2fpjufRUQNqTRtdO
I4BFjVtvbAfX+CtrVJdBvAfpRtwcF+YmAoyZY07DvBr1I75tSMjcKCJevyoLJO+aHGXSJQ1LzZbD
1OGepjL+3yKhciaxwNCzWVkN3MJAV9OfKc5eTaGsvZRBxwATemMYqtWC7DxySEnbFenRCoDtaTyQ
Ll5OzIQfB8XSSuOXjkCg0ZpECbvF2Ugm8QqfVTUZzBncGKuYMP0dhZeX0Q64Vadr62iZLUb+JdNe
yjv8qPN6OoG07r+fzlA7Q5/c/f666klzW7MWQ8u7FHE6eIvSZtrwOn4UONEJubLRcjNfKAU7TXr1
hQP/rt0yGCZeuNquFeXoliewNJogIeWoU/+8HE1JaKPryup0A3sjuYGO2LdQ3HjBG0yg1DWNYCJa
FX30HZFFtYmGL3BNxB1TGBDQcOfFeJN3U7R2gKmo68XKFSkda7EHiqiNgQO24aG6zsjQ1OUNm5wV
W/m5WnAQ6qRZbdyiRvbOacfoQtlSJzMyI+Ag7a6M3JCJj/zVUIyr2QD9hzbrBMGS+ADjRdj3KL4K
bwCZjMIyfEG97M+hsOPjYOJimTZr3N7zaD4buq7ILxaDrLTEHqktFeHK+R6vM8pikMojv2W/FuMx
6NjGjrYrNj8A6jQFA0tTxWVReyhdb2mOykOjksi5rhZ1ozwlvXZ80fHITJOLkR5NJ76fjkfwB6KE
RXdbtppbbCcesoIn4WtGhWDrnvENae1ifc6Y6XIXgHmID9mwsQRvR+1+zgjO7KFGgF0UfnZTmpXe
aZKH5elTph8RO+nMhkMit181nSYqMRk73A+/O+F6q0YU1SdriUr9BFSkCM0tHrDVUZwPjD7ImkSc
9UhnvIgKGg/Qx6afGvhuiCVd7R+o8FDyBJGtX9W39vagmdjWcnXEIorCC3ON4kSQChkE/wafQMAS
Bkpzf3Mep3ItcjZ4hVt9MZIyrBl6aVY9YqOMtNADiaDR/EghU33GHybUbZFT2dkzHcz8yO+9ZLh6
abihUwL5bRBiVFrmkZm/Wxfqa+Kd3WL2kAX4lJa+M5CP0W1YhJJY0G/mTaqkl43R5785uRqcgKNK
bSpUKi8T2N3FAamSK4aBK5pYl/nG8LvapmCmPJmfxhDoN3jwjyqSc/gDc5tZXmOf1M91UFIHB864
NpfxbQ95UmUfBYF0Awyd6s/TNP8L83zjJH+9hjZ2E8YCzwNvdZjlvsc4xULDd0ZSBvHikX/eV5KQ
1OpfpyjFf1FL+9k7wmGkHmz3Yzyx/QBmBMPJlLYQCXTxI1+7cjptHlmk7OAn+5yNP1udSzWiGdrL
rhyU0XTuEkwCIrJ1JHeoEcPfEYYv5vzVEpgGhC8DUlUxC0j7dw6rb0c+M6fVNUkNpsjNGKwwuM0x
rLSjNlLOrVoZ5h5EufJT7zEZraef/9Dxr++s58FHefRphtK84eSZS60Li56HcABHh+ngEGwh+DrA
7ymBpFxShrF/2PAAeKZpDet4VHxbpSAC23RGkHwslKCiUAqZdWQAhP4QQo+mEEhojISOyvc2I2bs
o0Do8MsDY6FrxHkkbgtD3tUUprDfdgv0nqlFPx1Oe5TRdjgI9K800ihMFRbXh7BcsqVFKoxscrlW
mnp+MrsT59tHR9rZjx1cjxFvUYopPbPTsoJiFM2KtfVfX+N/jbfyVcgqy/Z16+wKHLFT+75QSUGv
ro5wYJJGevohPtD86S/6cN/rUYnAkl+3iR8idLIQKHhoIWydcWN5SOZvuvEbfz0/1viy4gXRx0HF
cX8SxGxfAErXpV1LyuWZQgwzL+GXCg9Pa2Pa6BrbkDir3BLJ2XD2vfshFvc2gJaiHA9B2ck1F/Zx
pINgucK7eorhjlSMEU1PImcD9tAF80+fbCBOUTF86j2yShw3NLVYTASVfw5Hs24zAabze2pSdKlA
S/cGmAYD8DZv8tSyH+hwSU0aAiE3D2a+3x/GbDxcB5XnpBt/3aZ9yLiFrbyqvEj1kSp2JKvUmkYQ
YwuLwg7VPQg7g0jSpxdIbnE72Cet0L28U5P+rxVJCxXHw0mlhONJrIfBOw4f8YmI/rLX8+CJlJnV
IfVr/XN77XV2R6lbx8VkkAFukIcL26QEXUQijAhoaCL24PRNQIww3iLepSy4TiLDp/wmtRsL2hNT
e7Ax3/F0lWSbzw4U+lovmWcoMF5WVmXDvkjYLw3LFlVyktTcmRkfU330TKXiEQYKEEq83T23krjy
3ygvw4mO5x0g+vcJWOf8p9biMcd4rVaXOggGv/aYRVcWNylOGcBu9k7ZJiWHbYojDqbvGaPCHVIj
tz9/UPpl/Yu1XBbl2EFLsNeG3N56bhVCbaYCeP0B9t8EJyCB2UimYAdmYXEOC0HhKKdhGxDWfb8B
/7N8Byvlkx2P9NWZ8RiMBnC/xY6Z9qoeZ2ICmhnXSLYjKA8BwwC15l864fK7j4rnB0opSk50poFz
GrRGtJtDoOC8/j19utS9EnunnOPe18OsBPeslkBXJJamB4pvvVPwO8P2G+YGCpc5xGcIFOYOqtMP
P5Yi/99gBdKk1CVGxP65zGqKCuZNoos/Tqyc8VqkLC30HFDs55m7zmYSROSmAFqDk69q6mLq820F
/m0UWL2975HvxFKojGxGb1REuirROKaNZfJO4gMVU1N8lIC+fR9FRp8i0pcl95spjd8essRXPOSJ
4xmTGXeew5OC3C/xROWD38vetjcqtyEoTNS8wRrgg7CQv1beaZ1SAwJasEt80Er0sphUxaTi/rUb
7OWAI9lOZLxQpCHZXAd/FeQ/Et4r2oAYbqazEuIm0QDLt0QvckROGwn38UiECyVmdr/LQMQp3ZdK
Op/MTwpkZOr9YdxqRisLv0AZCUZNNuWJEi0ajTWI2muINYJrY03AhefhvZSfhUIxoijAgryPdYUi
/sT0l77/bKXL1JtWrwAJkh3s0VS/Ri0ZRQYD2MBgektNU+l1+1/VTU+Z9AD2g/oAEalh3kElcUQb
5VbYOicKx6rohet3dmeFBmsz3QX53ANm6FqKg/B3S9z35apt3kbov59fY1y/s3qhjcAq+XuLOReX
9ZHg8cUXmedKjkejNTUrV4OYSju8Yh/hMXzf88xauco92/hL1nODXmwyPi4wDQLO14RCMmjjDs8z
GFTLIsoWz34wE0epEVbDNY2hurIWj1ThA+jF2uo5njhy1fUIAnw0TFC19n/QTjgQZMCcU7oo/VYB
wJWn1FU1tSOQXtzE5ULj4YELn+O5LInBH6L0QGHqP8gYRA3tZ9Jmotz6bES1i0XTroezgSXENVDS
9jVMgkzpj+KTBnxtE6q1PnHyopkQipyHrNgzU/EYya7Mhyhh0MZG9phRpAg8iHSYPSu38egXwaOF
os9IiC0/pVPbPCfwISkpgDCFNXuF3/Lm8hG/2IJOq5+3lJmK54yRwLCASyH3Q+cP6xz17aNky3Hd
Z0otPJxfySdCr2eVZ/d+e12J0EzXbOknhqCjXi38xmB1UpCzztB/AJ8x+2EXTe1jeskl90BmCInQ
obfPv8f2qivseuu0CaL3pl+3tKYFOur/pw2b6EidblMf+wf80whjWKAmArxQPLG/zmWOsmg6jIRl
TKROuy4tKX5aZ9JoctCKX7UJL7qe8oKUw3IVHsE8o60Br9NjNLIJytbF7pGn9Cif6x/33CpZoa1c
1WccnzvyrTDK21c6x259JV2rTjrd3Bln+qFQx0VEtiY3ORZUugmPRmU1OBPQcQE2dKdUJmWEuKmi
mLuLiqrEu7pwGaq6B2fDJ7xsCO1Idx6emt0jYQMYpHxmMEXRvIQZyI5kg2a3nuz4KaKao+ndt+TY
JkH+vRUO9n7gXxTPtmHSu308pHvH528J0MEsvCCU3bTeXmUAEH7uVsOMgUeeqAq7SPWVfsAqnZh4
JgtriXU9M3cxHeHTOeNjTdH81eX5mHMuBuTzVdVjbq7EJOQazWMRRAzvTm6Ib/VF7ZQPp4L+FZeU
fMZYPfF9llUXU50lqtJm+W1hoYrnRkiYQWTWhwTcOve33WtuT5SOYNySwNpcG9WvwGIlJJu3D7/G
kAvWkNVffFhkvIlymz1cEKSy1bbOURoybsMxH9V8FWkz2J+ct2pIEJtML/Z5tH9U/KJ223PnMV+g
4At5RqGBQO1ikHC/KIdw25PNHOXpTXPbQlfLGpHqT1LRAp/hQts6I5dBuwZ6o5+tdKWU0tGinwhT
BbGl1tfxL6XbgMxKVn68tdp1rTOr14Nm+qEYkPL1pZflDZN1iqVbk4eNT6wGj0U+DlHuBaKK5vLs
A4BjX3JaXsa2NR2YRcRuod5RAYlj6RtxkGRTqki99deY7QanbHTZ1jPIg7cNE7kTz02QsizI8nLk
KSBusMH6UGk946b+mGZcWyl0cAd3Yeju/qaheBe0+/vfFMcGChUx4WE5EHQ+EPyjxyaL0s0zgywj
GXGeZX6JeRU9pTnlnnvCq0O8flkDNk3+tn3fq1HMqg9hhugWSVxAlaVOkdCUvTpo5eQ+EfIBLXDn
7pWpKkh02vCrkZcMs0Es4yBZtNaErP7E6Vn0m2HL3SYhY1Pj2WGEI1O2mh9Q3sqz3mY+Ldv5l9J2
aYZko8YA3sVFG4RR+yceBGG2o7C0g62PJrogum6S91vJ42KPwBN/nMKDfbfVkNvaV//6KBaNV+L6
mUDgMbCtF1ORMp3VRwPB5WJBlZR8+petTVjkEu1woor4b6735q3N1aogNLDYtEs9DQvwQcQ1S8oN
JkT0c4qq5BVzAI3P43sLw6prccNHm8rSIIPzf0c51/8AAz3BlI2E3OIDB3vFgQbZkd99hAl/oWmx
mUHxKPzjUpp/KiNJqj4mVmlZOl41R1IrBlainHyz+7VnwmMFBuTeLH/RHHYXEtfZ79r8+C2x34xR
kfeKTbyj6ww2EVL3AguIfwKA1KG0HtI2fjfLdBGkmcEVdBzEaJGsJWczrB74g1cm9YwUOw/gn+kU
Y0EVO99+SaCFmHhdeXTeEwo2iUAMU2EWR+WmL2BFYfLsh/qqUGO9OKhv2/DjmcxceWC4dApuZ7Cc
WoRSZi79rV/bhoUeHLk7dSY+xUfxjciMatuVn1ArDYMym69AAflY7YMnWD4lP6sb7LOEIbwgdphy
gxXoWedwA5lQCljkLJIOSMB/I3h+stDHLg0L8lweaXHdShmlwn/1rh9wijhMUOMtjpEez8UNLJAU
fBfYaaSBYhPJllbTOxeF3mccCG/UGuWod1Ifbq9ELWSjZqs3lq5luRv9VX/UP4meuEF1qg72D07h
gGkOR8IM1Hv3jRVfLOUKKNRbzo1f7Fhr+J0mrfHj1vAPPwhwweAvzBm8iZyJVH7M1uADTP8bF8k3
JJG5CuF+HPNg4LTmYYVZgOh/QhmKiqbKazWLnU3IFLqVG8MTsvNyqaw0fDJrHi3Uv9RX4TzDtI2N
lA+nft5kTvX/LvfXsgT8GymTajQt6YiZDtJORlYIMXPj9jMn2Xd9Jw9m75IhYe4N6hCCPMHp0BNC
/yC/m4xrI3S/QbQLuJ9+8gK6B/JmGIZAFEIVLBo4m7Sew0ChRDdO6dEn4vZ/wSex/XUbDDD5yeDe
tmKsTHAvO9bKmboU2NRK/0LAHe7sHYsBXZf2dyiMV+vs94cgvSi2dx7HQJqCPRA2whqCZKJkaClH
PmkZE29aVlUrcNZ/wVtrzNYCLRV+nhOfy2iBwfRWq2jViunen5U/IYkLXJ/c+CirN+azrRBIgMUi
Nq7OXDwpMe2EFWlMCr8iGOgBeA/r44Fp6IaZpcWpxFZRLRIZbZObMBDH/hQpUiDcy/Pf8T71sChm
s1V6FRNJLcCpi9xvuLjSs/LCQkCzpUmecT9TDnig7hnquiYnZJODjq7BQUBZVsLCwfoe+neNxkDk
afBvTKpmoscUGrzSU6Zhtd1FmmDIE5n33LvvVAG2sa9Gb4ifzLzzv7k9I8f5i2qk7jBIUDUQBMwx
ozfZyRJf3SR4bH4gSs0XhTFlD9EAM8ZzeeH2+usexVd9qPyTOPY8FURy10kSN79Uo5dyiSA1BuOY
YPB4QtfV5gfg2BuMQ+N94sF7VcifAB5CB/HzFapiV34dY6ACkbttHxNPOpu7gG2EarAgp1HVko4J
5Xqm0cBoNX+DNL82bmFeZIIpGf32CTlpYoewNUyKOzNvkOm115Bpg60cljKCkvbH3GrEo76LZ2cg
VY/rPWn9hUvdcYNbD5i2RHzHS8QqGWsS2DXL0HJefrgOldgXpKInt77P2GQgNzXykLSiQ72oiLDy
q3zkMZ3TiePP0UXWRD2C+hh04ddvVLcjmFr2AXmYYEhpJlBqCtlb3tB5QBTeocCGymxhyVDZMMMy
FW3AjkJ6kocw6h6LcvcaCOXkSHZryRqUSS7emNHY8exV1MXqVfBbhbCRFpK9cCFbBUKy8xPERDV3
vPtXV9xQ9aJ5Ro1JouABIE9nSL6s03/L8CODSRJV1X+Fsbd0fAVINJU1XpLRSupNelIKaQhlf0+n
BAs0aeoGzgpYLOTRB7DdM8Vj7zC5DiOGlrk7MtoaYpGJ7bhlMg6jKWVCyYkzfCVZlJlvyrpxhNnL
FLNCQ+NTAtOTx+tP9psIki6CNzRTM263pcsSW1H24ad+fHQtALXe0rjfk9PXAxNahI4knI0XIS50
MzT7MF3L+xqZvNUQKnBit5ntP9PJjGOzIxsaIZiy9lokqQf2M7HYjyuawBHEKft/B2Yz+MafRAZj
ESzKDMlsElasLoDo7LU7Nz/HyugOc7W5R+T1ErG/gqMaA9h6k7ZKHVHrHk+otV4H4aySHiyYg1VI
8n9N799uW5RgWZ7V6BdiJ2IdPep7HJOGvtp4F7uQJHoKCNBfhjgew6bMKpZajq/rnHs28yhmXNLY
Yc5mfoZeMwqM9yqrby6bH2G9B/jN8mN7AJcFUC5259tQlH/9TXDv1h/8RiMSkQauzZ69XKuglo+x
q1opttF0PFyMOPv+7RNOIlfz9Hk04MlzO864FrXUAQJ+eMtTf4iQ93euPW73jPSUXwsgrKKtSyIP
R9psf6ljEqgHhOwni0nikAv20AaPGX/736YhUjNB6GqQ8BgUX3W5b6VZ9Mya1I4TDkEkyBd16t/7
TvSSUlGRlE2/EVtOzv/i0x/5xC7iWkF/iKYy/TMrQWL8dy288Jlrhyxb8LX6qMYpOAVlowqBZd1g
yTZ/9XEpnb/isQ1Nc6UL4zki32OfRbzjzvnX3v/on/7p69g68tTGBy3Rhqz5Q4vWfpbfDfDhoX0X
JZAaUUVOq4j5A1Vbd7YjFiU7IbBktjAX3SjpavakGKMDDuJr2wxcLk9TjPOnKd5nnVH5kE2GKqNe
3bQKS/fJgclKH3nxSGXBv4p3d21Fz7Xc4rWSgXv43f+Ui1g3QDsmRKW5AvxeJ8sIP22WhhmdIUyp
taV6teFhvkivGQphq8Er2Ky+wbo/tJ2s6PHI0/jY93V+lOja2HkC4b6Jd0I2FAI7QQ2XLJSSorUm
V+qPI2+oycjAA7uXquXBs0lYIVogbCuqRB6Oq4bL9i/GE0CTeFlrGHL4OI4lItcOpjNVnxQfEvgS
iuymyclV+3CXzpiUEZ039C1NgCmmIUVrTQIv0uAL3uuQSPXOoXJTOw8lMwSzd2RfQGPA5e75N5qe
Q02pvrXS7k/t6E2f+cxP27o7Jl4dbgVGy+vpej261vun65gZEwhn9PLI3/y6xP69aNHkfEA+GtT1
v8ejxrwUl1wTTlVOIVgBAdCB7xNrg0jFlTjk2RCpBnZrDSeANF0xtT0NqGiGDNPSDIwBkNtCTkJ2
0Ant/w7/Hu0jZSoo5iMnbzsPY9E2iHetKPOfFhBt74ZN5p/l0gZ2mezwpB7RxvpvEYHpXGQvKWcq
BR+wpMZxFq+FnqgRDGaJYwcw56j1vWIx2jb8KD64V8aq2zSeIk/dan/Okiv1ZgzgNWr1PBmnspON
xeQE3wQueelZlI8kn/C1B+v50qWsX6k20nHer03Bm5UzbPVeXWlNNPc/JVl0RLqmY2zytyct1YXu
96kKABu7JqZFWOX4O0OVEYUpmLBMLcHIRWsW5rJ8BIQWf4XrdZJcN2zlVdfgJMxeTrsZvxrQ+Sd2
Y6lonFD6l8UxSIBKxfFornEjX8MOcemZFvcf9aXtEzkYa5CUlsbOQsj3Js8W9lCgPRPNU3DSHtFT
dCVbjzgX4B4DLNoQjODq/V2yDJoWyIma9DpR3zDhsoacMOI+7fqI3UTTlyAv85DJt0Cr4GFQ1zmh
b3jxJrjKfEdt8bvhK24BXBhs4N4OoQdBAa8Cdn/8dCk0nH44Y5HB1AqApndAzQPqmsRXEo2QQ0uk
dG0EhegKl86FKRBr3oI51Ab4zXu88khoXHw/A/MeerczwFUfHR4dRYZsIl5Jzm3MF7iZ6a0hJ+ee
gER4XF5c5FOlcxgTho4zQtozDIMgqHkVZHpoa8VTKMGguItjuRVxkU5W5jFMc/yNBG2I9IImlGsd
5BDUOz5A/6GGqApXEa38977Rb1IDFOdTnDsBwfXLHn1IPPmvw786bP1atnBiOn6iz38b0m7cbtVM
LqxqQvnApoAry01JH7cQmFDpSGBPC5RqSjbJPadPlysWRsf7ySwsWAPUN+a6kPwX+3MvgyIIXQGG
KN09NKsGk6afAqk5i3CvVsDURh71yVj2caUl3e+lV0NkPTW8kxLEGUdo76TpluO6c+wYUoLW9xFx
RWTOlRsrcetvpP8VQJtMCGDhF+cz5izi35Xetm/fH8ykaoQC4pmcAtUuW8aCHZYtxrl2PYmv0xx7
sgcCQ+A75COLgdaGqUSvkrikKzYzGxV/v1SeXGg19z/UGBj3+a0+rH1HFl4cjxndCNrH24VYU0Uw
7iOyAgEt9VieKdsEVpHDPVIMuQU41ZzwbnLqi+gTDoqTupOMGk7ZM7ZMAALKWwrzst51dyW73uR1
feK7WOYX9ts976NQfnMWWjfwc6cLhHf2h6yFc4a3yXptIy2dmYi+tVVuhJooBMfGqVwkc8Eg7ZLZ
GNcFZszMZ5dQq9Jzl/tibnFx9zRgHQtfDaStsWDZ5dB+/cr9LsuQgm49or/vesq8kDGx/uOk+ar6
9TNVq8E9QcRGd+ISzOR4s8BljS0CakpllSjHa1hv0IYdyknhWeHmfRQz0j71+EpdBvkg9ZAtMArd
fRIiEFruT9fWOTYD/cKIsYnyQHHGKpa2ixZo7e8On9ebj+kMIfJRPuEZLvzWy2GmP0mK9R0Zkhev
3r9PEWzWdZd3fyrHmy/NKEB88H7z6Ok1pChkQHcZMLqxoQ5mOrgc14G+uAoMhrUrM9Fu6EqzcshQ
wAjOrM3TtS1YNH8cobBh7lupW6o3eyCLwHOsm3+9IqlyWASQ2Ak7B1no8CXrbgmFWEyEfsjsxdZP
WV2tIE/M3iIc9NVSImuPw6+WGCbisT7vXlB4piDqBXVg3rRiHUq6prDMKY3gb/mndx4XGHeg7Kli
4tuO59HFl08aa+lPuT6tbfz1koPWigQLAdpO0Jy0MaRgzeywcE4zILEthLoeWlLcWPjmaCZBck65
wi38yJo7wOa57SvJtCcCo/w1F4Rjep0fBud6AEZ8EChVAOR1yM+0/Q5Se6il+dJQPSj2z1Gq9P0J
Z7YZBxc0j8pKOdQaPTDUfyTDiZJarjwxIUwzZnr9LNc74GUOoxaSPUHQnKCW67Y9Sqp4YIysUfuB
yXPi9X/q+lzgjoh4uY6hzojapaD5VYv1Yn/a/CS/EhWGGTa+n4hugeMSDW8xAFmxm7nPeiIKWjIj
cOQswqQZKn32HZtinijhQpeofNDsKiB5lGtdjavuwuOTpZqxZ72JbYhEuU/JvSu3Aay89bhZZSCu
BpaFVVTs1N57p4PvfeAtnahiLvOHMFQvPAthOAkFxFNpuASEF3SO8zZv14b6R02WZmlHWc+OYhq9
mlo81a9itXcD1e4UXOYln4HWxPK68OCGDoxHZYzr1mRfxk/nbaRt0AFnXo5tufziLZE+pmqeUO2G
zyoNyHvRPKoAYg5LCfWJJYkEhZC39CyWL7workvLXMglH2gB6Mg/XrswhCGBmUa1Xki7bdBjyT99
xHEarF9lMI/0u3SUgeylE3V60MUjnhOaAuVj9unX240A5vC6hr7jMIKsBxDzzepJwjdkDzsLeJ79
h0rtVGDhdSe0N+Qq56E2PkT6cN5XW9yQXxmOyhndNOiQXlrSAItCHMWkWHIyjWQ3Zvf0ho7AyWwX
T/5eDMeG8Uq+ybjw+k8M1VBgFMxdLHG8O3PYs3FRGjFooPoQrDXFaLBo/LFWWeFsQ0cENnRAqq+V
jDiq/xjgsLvzN3v1XhLA9TJ6VD05iaLk2zdDBYK2DZCOgjoVUK2YgSYxgJvGXYBqxAu62Skmn5+C
pIkrMAXi82r/Z12grrN564D1KVP4q01huf1JeV8LZCiUIdYXgOXWRNW2URD3ny2czdXSY8KiNATE
aPhiUJak4XHFp3HXU32MRyDmaqwdtqVMJni599qGeHS+SKE9v/6YBcWnHehko5za6LqeNUWgJ3iN
TXiWk000+ajG4jak2vu2HTnFdAMXwKtrlTIBG1twO9vFFewTZscCvTl1R56ZY+o0hDKGsFbjpkHb
0lMOLiR+mtRci5+vg5/IAY/M80RXF2YGM/kMpUytbGUcj4ibZmko/+Pha9vEpvVNhf4Yf1Bx4YS+
mQBQ3xD0PQnVH3HHYE+yX0IazY9LsiMuUzbQ5QfH+rKnQhGua1BJKl1eHfdT2mkxlcCzZFGstYZb
Wtei+HU4G4vuVy3QryCrc0MU+83AEu3tagqiMWTSUb/peAqzLQp5q7Sf7DKqk9fz8klGyx/s600V
4lYTFADUJAy5SU2ZxeU1+KKeqAtcJ10+1jyHl8LHkFIhPS+JEXOLwC8hQqqJU1Bys1c2j51jiOnS
FIJCOyV+VI7tFLjMLIbTLwbVs4Qbg3zfGkV893HKWtUhRBKmEZ4VZSav0t9pL+zPsI9rRJ9j6LXK
zhMmKC2yJ4wniA/WWhtfBwzPc/PblQEiSVu/GpfLWfEpjG48w/TFN0PWwaI5V1OZhntI03QLujZy
s3QaxVWaQI+8ObFrfiQazTY1pNulYoqUWpBkFRl7KC2rZJe5FOtth78PAr/TSvzuiZDgMTxlFp/O
Ur1Fr3mOoC1a0mCYVw2FcPhv/idKcRcOzslHzk+q7imI/IFauDvsFYoBNCTdpWX2dTs2mtQw2pED
JALzuQb3sJTplSgmAyeRAgn7sm3ch7YZmCzWJlim1/zbMH7utWYXKFxBRs0xC+33weLPF1AmpfKl
AU0v3kCtfe/gIAeqctM9aIcvE3M7n96lcClvTqBqiVynOjKT0p/HObz7qoZbDhgVrRTLlvMbol0a
5FPkAQoZMrLWIvgT7q3pAQm56QqrwvPpHS23xVZUYTFlYBjyKRBYNwrrQGXWhs3Z+xv2xlPJwoN3
I/dVyv3ZVf9McGZ402QGNMkQCquUGHr/Gn/cpsNnHnIcA56ukMD78KbxHPGFaJHbHoZMpfOfRzOt
cPlEKDmjnlJwoe8yDtJolQ+KEs7ujqbt8hvWlLCLHTZZeKXNkPpPywcyTVgGvkXXs2GDWvrFOEaQ
Qc02JXZCME/dpNVgwq1uzrweHl5AI1MzujKixk0Kw4x419c32O+8JMnACG1dgxAgldoC880cLvIW
tIyeFP7W3QSOaLc4Wi9ZI9DbdSylOW9d8/UbD6X4vNzyZYpzzEq/1CUn2j5ZVr0TAYJCNcBh4fT8
Xd2kP+MjN3WYB+t5ABT2RZDM6TFKBU1Rejj4VxV+vQe736PsXm1C4eJU+AoyvSl7TWwB60sQaXZu
uLuZOIUsS9wT2qMTlmZ5T6ejVdCapKDScedAgxIuYUGXvCvrUQJRFBX0yHo0u+hRowVOOARmwtm6
Aojhotm6I59GZdVDKcaNlqoOp9cl5oUrzk8iamtFI+j2IRbnYiPDdQa59//cSgAxge5fD7VLMe3q
iTv4D85kakd6puLuoNguhxxQw/R4CSrFpVVAXMFciULnnhi3g+MhQG93/9aIoGn620gbCUU5cAcx
KGJ5I6X4yuWJARvM88IYnUfe0LflbijBvugAyou1Nwbfr6fn3fo8ZDunyBGmyHvcHWi+TKXnRYWH
L6KC1qG5pQ91dvJgYfIWf8hYi/cU47volRAkFmmLAWtB9J0gJFHQEMWk94/qiszKnkwBH3mQCrPo
UbHNoIuq8+ADmzD1zbjWSnDbNzY6w6jR0ZL4T00lRPP8Uw5K9i3W3GIiwnGdwupnOjTa6wnITRMe
JJIZXjXipDtMymxn0SLS5eVTPXHZSXfUgqzboM2BcadpqVru+6eKeURwU5cgrNvksVstmI1SUIhn
CILL8Cg1d/Y5PNYF4Wt9l5a3DlqIp1quBiZ5Kz1yIuEK/WZx6xbdkDIl3P9c5hB8FY886TrLH4ji
WpWX/C5j7COSycLRTvY7i7LvB2T2o5KvaL9qoX9dVtnfeoF/aF6+4uRZIvigvibD5+Wwr/ayhneI
x1QCyWNHki0PPpdTKqYmT820pt/hno2vOpqA1Mok4eP7e2txFuegN4yuzs18/U3cxaLR+PmFPGd4
Z5Rgi4b63qUSLOm0SkKSs2WTbPUjT0qseJvO5tcVEzGFpLBLUIQK0C4LoQBvdTbkq3LlPgaqYdka
DlQbA4NMAo4nnSrrzS5d7r5oYMcyQTf+0ZPNQtiCz98hlEYI2ZPYtepJ17LbhECeHG/d8Jzt7MbF
5/PxVGIe52Mq8yhoEXPWsjz0nqrIIQXIjfvTVU2BtwcwZNNawHtNsYPfXu9IBqNCG393zzmiul0y
G0/HJTaWz3GXBZpUVD+UK5qZ0RgNe37s7xTWsQcNtPZfLurvWh+s59bZBNxd2qIj96XBjb4w16nv
GOWSfsX46lYrIhU65LTzIkS3cu+ClTOz7tFYQKqGfrRBJ6AbpEdFjs67Nsp3U6x0wgs9e1QAEoOr
tHSQKr6W58tigWAmeXSBObYufxGPi7o7pLTexsZIzGtLIxF8TdQ/XwBTWj94fUugw/gYRZDGEWGK
jQfwdmmgVsPwGqr5KvO8bTCkol/3ilYRktrJs36PzQ/DNtnITlTuRYZ4DnL4jp2XlGR3zVEtKfD1
hfwzsQ1dKeE/nPOvzPL89XIOA5MJAtsJqfPOlY6YcMwZXThO7dZlWIzdpIAVj3gSnkboXmMq8N8B
m7vGFkyxjKLWnwWQ4QkBwEIornZUWD4pp+RYqExVMpf2Dl3LbJLeF3lbgUbkloverclvfTKY8nfF
fDOm2VErR4sG2werQLP6e3LD/TIYNP7Ohl33LNRR4roojTRD82Lugqs0UK0xmGOjlqrLfsrh0ZlS
hkCW+P4Jq2bUk8kGw2bxGaqPVr+NOZe3q+oRlrnFymjFGOj8cl7oqaf3Avi0CLHQQAy3g87wfZbU
oZA6cnoOMr2CE4D1opDHnq+oBHKTk9INx1qHk7p4wdBztIjyF5lffwiKaJQMPJWc83OToldxSWZE
L02qho/OJzP4Wv5os1nlKgFNYyGgTH8SYfe7lLbtd/iQs2V7+rcW5vs5Qgamkc+XBTGKtLpyrBsN
7+Und1UT9X7UDX7myjf4EJjPbNv333CQj1CfzC5fS5Af2jN55uJJuxokLIWMBB+9P+nBbuSaiWAd
AOM+bJrkp18lTHgpQXpdwoIeUl6EXal68qkExTbX5WEMfxFEwpYG88Qys8P5BPjsWNcAe/DMi+AO
flcPUZBQHU5EKtaC1YO8By33l8VEdetaQ8ZpCMU4SfY0sgO5NE6QuLGLT1EN8DDJL/NpVG9nxtaO
tFUt2ZK6ZUCyGmmj4Mm7phOw4VwDymoFer9HmNbHtv7mUJfVURCpcCRX9oEz8mDA9fPURPdDBEO0
XHsyP/xGa0rVUaxxu/cMVfMfjBNIHHAIoBOWCZAuaVIGh5xnQg4Qesc/qwNCfwmfxFXsxoQLmVnt
WN4umr4zF+zo7kwlrLYGWzhaJeI/6mYkPXmEdfY1t7+XP4VYtvyzdj+W/hF7SgkwPcKGdapmImHN
6M+nqk7NLED7X+0bas4bDINHRkNA8sSVl8Sh0lt0B9l06krZHMInBy97p+A16P7p/Pav/IDGmFLh
Wt3pve9XiA4n/XdCUYUpJ0Q228gTy/5gMGKO1NNPEXe2cYh0brwgxnljhoDrcFHYf05o48iK35Gm
0I9yZcMA670XpbK+ORxlZafPOqweevFXHmr3CGxYxhst7ipMaI/fNBSDdoa3AFgtDzz1/g1kNMKZ
bDGqN4NtTdqbFotF3Fnk8J6p3fb8K7J4ZOQbNH7armVxmO/oufMhnPxqNdxEVBX5jKaCKGXjxDrY
ZAU/PHUP7/AcCTyr81BRQZlNMd98n+6uEIdRpzv1j3uZDssD8uvoNnNJt8TYeNTv8JjED1oewsBl
bqBUiQ0IyWBf/wSRSBHQDExQlrx9s69YX5yHCzDT1jCFZn3RddV5plKzHCZcb1UtrxnJgFIcvQ9U
c8wXXFvtPZUyRgiAoRvCgzgDxSWcRtJv8ulbUdXWuaK8ZZtk85a2QolvC5Y+zQu53L7pNe6V5w9O
SiCydSDz/ppE9sAwSB4w2PA+eKxHVB9kOnuOIZGFcef+WjLS+DKJkM5V4hOtAILmDsQVzvut9cNA
0Sn29B78HFG6m86n6YSr/R1mI/1oVqBGG9drJmL5RuKCNn629w5hgjNYIBpW7Bu3qz/Nxo+we77t
5LzAsRPgv3Lc3ZNTbrY8qzJlds18yQAv3CXbkA8+EaJQFUNpgSN+vUfGCo17wfbHcrAZpaUGAuMF
qY9KHyqpedsPdlunju97l3MsiUbh3tUikwVDHT8XKfYZBIuJx6FjwqCwZzy032IeEqtQTtF1/3mg
XKbJ39+U7O8C/TWrSPLBmCfn91GhWjFOfeGROHp5C+Fc3Z04Fi+LfdV4J99rk2jHNcu/l0J2GPdA
FR3vb6vfRcmd8E1+S0fQSu7E+auxlwaFJB76THrJOYRL8z+w5kVE5ArHervlpZQRp4TN5QRhRzKT
pyYoiEXlS4o/KyZOECSJWBLs78/XjJLWuNpU6GtWSdwOZx4YzUuRA1lU5VTz1oS3EevpRIT98Q90
4U2pBq3VWvBok3wA/QkK9Nt1Si4zRbD776nZgaQb+pHSEEKPV8ni0f1WjnGYTDZqqZicdp7A8i+E
3wpoku597y2di41dla9OQNVXwLruwdHg+tQLKOa6qKHMDhKhyGVYC6hnUjlKLSvlaMMTEw2LspAp
w9Xz+LMu/Dh0mI4PHJfWnM4XblaaAkKCs9oafI3UCSYNTEAaDEG2QyjLvKFkZyV/9TnEGdnC8bDX
viXVtubuk1QXKG16bS9xr7D8dGxEUiosjqz5IMFB094uT6L9pWO0DQvchHC7r5v5AHITnhug/sL+
+z1q1EUtJJ+wryvA34MWwMts6YYLX9evJZVXxLCst0gaG3oVj6X0PrjPXUuqiMK0zkyme52eOGIG
UvrK3mVlFcc1gBN2vfP8KyrDhjh47Ivi8GTJe77cUxNZ7QMCTKTOjZhof34KDag9ZluTTvQ9tBJ3
XPj6E5JPFr/IdbMU7Sj8r0UEeh1u+FLdbXONu67WKa9OWU8TIeY5r33iwCbSgLkzEMsLQXyh7Exy
VcNBuvMtARlqFpelbEgZdNHWcOPLgnrptcm/Gg7o5OSwyv0tTnb1AAt8gG46LMF2grnSuQH6Rnvm
o/rrGqgp5hGRX5+TxallveZbc+5gck6WJ1+NPSHu5FtYFLyvjnBU5b7cYlhaIoyLSKw+R27R6/+F
rkVEK9Ta5cXu0NoFk3YELqQAZjmrRfYuzOe4KXU1O1IPigHxffLH2jmT0K+5BnULQWmCLRsKurJT
XXgN7dUSlGAw7+bX0CUxyoXix4AyCsjenB7C+3FmVp9AQT+A6MQPJ6TmUHK+lwFOfcrQvQcgncLo
AKoifYOHlQ5PPHcTGRkCtBKMJiO6YNUxizP1+przyclAjIlk0IJ5PpZiYnq2GCSV2g1WCXFEFKPd
2FbYZLbzTsNQZhYQ48ibqcagbojfL+dcNBDK26x5LGBHipaxKnxMEk1TPQZA
`protect end_protected
