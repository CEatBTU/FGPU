`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oLMxQ/1qvrbxYPVC/PwyL5tU2URv40SXzqSl+pPUGjic7gu1Plz+qIQVVmEcX1Ay5s/yRbdt5ZPK
wxYr71ldng==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ET2DOXpwLr32NW//eG1vNBNE+bhicUBuYuc//vrFQYAKGYST041fW3S6MmjfstgNZYLMXjSbvxpC
hjo+AEE328TRf4A4Zv+GScq8EPTUi97lzpWXixJaJ8JaZJ33/PvQKfMHHXVeynvoFa9IjQFs4z7K
NYqM0eajNBll79+gz1U=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BhKOhzxLviF/SJnJL+pQ737ytznHDmJUFEH5mpC0QFysnXntHYAo5hlNwftgdzBHAnTXpGe30vr/
y6OgRKikFfJ8n9gd29it5f3PFV+0p4b/LkzxEnM6mrRz5SMUF8a18eUrVtw7zQrMnpbHh+5gZ/04
lMlqIA2TGAQD2W1xoSY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UULVT4dVdy85wL02x+7j5fmY2fLnOJwYgBA8WDaWGywtaHkqkaa13ZzEZX+3gXxQ4wKxk4xH6Atg
WYlmy8Nm1anokpjcYPYtIxbKS1fJ6hJ5TU+oMLRxzkji9q8kicuaK8cM7puDayq2RTHl/bvituFC
rXkwrS8ArIf5qYbTBhoxf/upO4L+zWutcwHFVcTiQB01ok7R57z6+jJHMtko/kKcmQKGWBCUFk5S
YlyvQLQYyi4+nft1fnKSnJRdJzQ+gVc9JI7xsqR9ouq5bNjd9AbpJm6sdjq2BgGA55uusSgTGe8M
/WUYI6iAV7tk8PYXwTpid4iIwF7hqcKPYl4Ksg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I3M3k12VwXNmLHRS5YdqmWaOmj3dDbEFGESqzp5j/9kXGYLmODKyJe+mrR60aM+jHkf/JvwS0vZS
M1ukjw8Y0xcx7luEROhjgtxyeq5UUTxFDacevkJxU8/Rby8rvETYhXZ9d0Fca8ZTSiF7N1TYzpRR
tOAt/35z6Cdk1NYzun8JAj4tH9cZtkJA9MRXQccpg1UZAzeR0faN6ewMLyMziSZgDYmyxDuHibfp
WXzvE4s/GBiN8Jy803m3q7EfZmzfgN+vd/c4hvvvCEsS5FF9UuT1eJvCfHd1c4JiI4f/xUXzwbhd
oTeFnK/bk7iK/J4UdxKdDVLt02/lOTxkXLCbew==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kki7dLAignqZuhjmBT6W4JD+gUEbcZlmxAVBOP6A8VU3/ogIq2PQI2WytnUGsVkXq84foMBg/XM2
hL+j98SHnYQTl3R6jLCEadeoaNTlUg4GMa6hjQYZmW0E9olOBia+oNRYiRjHlOmX1oWg21PPfVSY
Dxn9sWblh239lcJuWArCfFUFub47Yi3C1MHqh4TIcvro3L1pNaD+R2tNcqwb/gdZc4K8+goDCcye
L//np3wlkWb4naiLjKngaQTcnBFB7KD5RujfWM/g7RSrKg04nbpM9/R/44wAhPs63CBnPAQnTjO4
EZT4dfE0W3FYnsLJ3X8gLlXr43MmM2DZBeaAbw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
xCFU+YhMkVQY4Y5PuINZyM9ygBYw4psUDR2I0ZlQHksNhLOtOSjMfsikrphsFtwtITtlNsWPFa+U
Ud4hBKB26uXvtpl2x33SyWE98ZHsuRQOd/unErv1RyX6ihx3t6DA/TppTz6slhyqkvT7TlutKI2R
KAZwBgTR2tCa4IQTTzK5yUFwqt6IrePELZz0J0K1H0fiQyO5zp/ha8ehhJ8vaXlEL7Rkcr/5NbtW
sOkIbd9FxsEfCmN0DLvH3hfD1xVQpO6dBKNxQVLLksj+ZUl3SJgqRxiUVUxCB/8MkaBevF+4wwUh
iq1yXm0dXTsPV25OEn85XgEfqvsW1UFhIYW4Qai2+mOQHcIkSPXJi6uHnsq+wZDZr22R+MjXdHCV
JcwvMCFalHb8L7QXg59Hy1WTrl6Z1KReJJKLte8lFdY1ahN53vjKp2S97uzV634RD4MdlW4Sd6Qk
Y1MV5+VgZr9KxwKjf689lgujxsClwpYMzb0itAIU1MgEaDOTWVLmIL2+wl2QMqGpMjvv0zKDwUBD
ZFZHbL4XsqaShWUUBvnw3kXm/NsAkM5YShEhvc5+bpq3NhFAvtlr3MqvWcV+8nI0Dm2dd6x8NlhZ
YZVTI0KElG1IvrUe+epiuRg6ybXBlF9SJ9V7RS4owUOGWzG0xlogrxIAI7ssksSYsXN5G7RGORTY
UmcLsfsnaPCvh50gqzitzFvRUGASX50IdvbFRrIRzcchGaOCXk4RrIFdQjwEwHOF8lSJDc4Hzsa8
/E+gkO6nyyR8gkMnDqTqd2H/Fl9+JEy9RZSaPm7bv3XmyjVCQXPPAPYsEnfPe3cDwe07HQEyqJ2j
L9P6r0Lj/rJT9DuGBQitt69CaN8k/Ja3VT07fT1IawtpopQmjdkbotWNeYR5k1pLSTz8Kr7Ep1DL
sUxEMbE0a+MIxA5kS/opi7+nQblQp+7lZkZzDljG8WJ0lY+TcW5R3O1T0RaLvFmNAc6mnsUk61lB
KOyL/9x7Rylgmie0/vNueIxrTSynIUVYV6YEW6bqfBHJDhIWB7sSAs1D6DpJUpu+uS8qEOH3prHc
5qxlqO4VvEKS9wBq0ugw0VDl+jOZiLqJzWm/hAhiptX0okbFBpHYmQ5ivD1WgrysSeKaU+NlA7NF
sXGpTvsdJiIrg2XYqI5/lN0mlgfylcwgR4D3xq09h4MPlxgslf0vnB8vb/Yfkt7hsGUahzmFNhMc
semrJOULPbEBVK+14NgUvSzWgh8u1qJuuY/ntuG6hGwz9w/+jhfJO8oSM9zqVCIYIN+YXyPsEurP
UVE5n2CH9W8pBLWsJBgYorL2djkR7otkQQplKqjlRxTSo+GiuFBU4E10DEmweqsYySwFstub1JsJ
KFtdlaB1DOEdkHZKxV8TJEKvSi5ESskAwTRs9XDyDAYZG4tvlNnKRYiiIiKBy/noKLOAbeul7s8l
Fh92hq+2DszC0/PFQTbdvrRJ7eNkHl5p+PDNHwef3Yl9lM9w2MM4ILPZmYyGWoQyQue1ltMXatoF
QdNF3YPHO8iBhoHuJ4KCImsBYmhC66oZ1ZIKiDM3J18GkGee/hdZnrb9EhuK44TmiLFKF8oeca+n
s7LnQqCZ9dvta1h2pEU6YQ9K13N1Ubq2omjmpCLA+nUbvwW3pHY2UbBEUi1NLud195kJos4CI2ul
iPQ6Qj86XWr63kDyg9VeQ5iA0jVi646Nr4tvzZgEFwwyqwSKWbZ+hmNdmAhw56XOileHXoT+utQR
lVJRx8evBSBsp+GQlAl41b8Bre8F1ouZ0gD3D4F+er85kUvOrt/0ktvQcqThXhvzWflag+3BxUaA
sD6b83BHOZG2gxlCLCIR4u0bC+HodO7KIKYp5PZ+4b0p/2Y5MFbEcfag6MYGgjYnUGRK4TQPTuOH
4oJdSbF6EpqOx30vNG89ViT0AdZ057Bo9QjEu02J/37GQrWSgZRE39/j3fSzjXkuCoGvvo/VGHi1
1u27CpMUJrUPEO4Uu8CHAZg/lgvFCD4lxMIuCxQeF6mgNs6L1O1L+tmxO42uZTDhnqqbmeXni5xr
nYdf4p5EMvm014dBnOmK/OApMibTuHUfPxbjA4rH+Ma2V9JEIwYESJdrt4ApJ2w1zCe5xhLyYzsa
rvpOplhFj0CC6dHCuYMS9vYTMYtrmCouqPuTvw7UMOEbAUX2FncLGaLX0ubWL9jD3GflX+mNGROT
q7Z8woOM5gbV+0TSO9AUyqvOXWGCdKVQLz4LTRycS4ij7t1avk2e8StIDV4JUc6cDyUNTGCDvMPN
nH5LT7RXD3ZVrS7I6L6yb4RTHGCz0erLehAPZv36UnTkHPSlFfM1VF9y7CUysQsim10SzOQOdJKr
8RSz1JF1vND2g/3g0JflmdGHPr4/GdR4D0VzPqeSOCUEoSXTErQENSsnxC8kgMu8YEmCNQac1YAt
CTl7a9Yay7vIc41hE6goOEQ+dM5x/HE6VvWD0xAr2O3b6yLs0B06f+yOM9vCUhU3cMbeHfdrOBqD
lfYtdxQgQvLLQklDmNOL+ci0jRr5LlUH5gBqJGxknqL0rOmsn3bg+brBQJLd3TKNWHNQtuygW/1z
NquYv2VOxbgyxh1eCGDHaINmWp36QtUK48kV/yfeDfjmBani+3XKTYuWvbY0DL5hqvdHkahYxL8G
+VA59+tKPVwo3eoT0tWu2BNIij2WjH8zTKK0Pw3nnue/s+EXHa4wR6Ba2VRgk+UbRI6rHw2TdmzZ
oj/6dn/fecGkYA3Myv5ryYyU9WNfQur8pwNOh6Za7s92MGrusjvoCjrSRd3HYUJUX9X3RhVwgQPV
ArFianyME/ghlu/hFOwPaAZYfhYSb+S0nksu30rPBXppTEbuOOR2KtiFypzu56skNA/p15Mpmgsi
xi7r+7wOpfDhrBbg8Ff2nc0niim6gklvE9vqVPKpBjIPghTgG0WhD3FluROTIjGEy144n8JyXH7O
fnt9wrJT8NZaEVasNuD/Si21F3SY8sED1eUvPHceir8YSuakxzZJkUn/0LpS+aS++ruzJEQMLOon
E2df40Vb3FcZFKZ2glTcXhs07d2Q/+Uo6sqrOSuC1BN/e/nq3mig6fF0Et3ZlP8PYq42j4vLLEqu
5c8SD7vvyXdQRe9bxXO97kzgg69fMIRvxGPJxl1s8tZ1coySH1RdOkyaebtZrKtGCEj3dR0MYbAV
+nvSXm6B9UCHt7trZzNt/kMb1Nu2TkqLC9DfqO4SUJEEdNHRLrR/1hwrkZXJ8TWRuIjsAOHcDBG7
H/QlB+VO9FyIP+BlYspM88t4VKs9kDD3z/+KD1CfrgvLMz+heTsL3TlH1aEttRJO4e3y1uY1ORs5
gXerw9UBbSq1/ZpKpkfa4JyBqEhdVEcwkoliLwJvYIZk8iH2M37B38p3obycIWPhMth17eK/rhfB
ZxZgUejx9VbqDR65wUwjcpVJQJqXztQ204fyRj0aTejpLH9C/B/eXyRsJ+5gd2KSdzE3KkTetjeJ
3GOxGZaO3+P1M2KHPjA51865vkfR6hEpKmOdjtW/zRcd4scJHIWsNsNN9QtXEXVIpHWTTfeKRU1e
X5xTJ35fqoSEJozDEtwEJoE//q2zBlVdKFXzUBBccK2zHF+vN+S0AWGtb5ge0EMCX0jpPP+1QhzI
S+hwrnxp81JDbQCMasb48tfuMMQGIZRby+G92Id3O8fjsYfCuS/dPPtN4SY0y15GBCT0bMReDW83
BWM5HtDlPzz0N9QwxHrQl5TY/dtXxV2hYvfvDALLtJiM7VBq8KcF4rjjjsj84VY+VHnd94DS6oOd
yIp8sFvaD5L5q7+EDzyjORn/rpTAYbI+v1TJOgrmEXs/R5/CX4xk2+UfRyV3AFJs0xvwiD8jsDUK
V8U9rCUVBVno3TNYP4ZRQOxn0NfTERZ6w2vHV6JD8Luxsx9xDltP+StzDLqbAvnU7rA0O1gzzrqa
0JMihlpYiSZrcri/WhbnCO+PHEbTM/ysOFGr62bGphOjOW8kTRVIy0zUplEq+0iupWtxeDGOUVLu
mXexTotEK1DYko/Gj/51rmFpWSCCjx8tye9Fxw2MkB0HSDZU0JxOahQe7qx1d+aCvOH3ahgA7Ha7
hf41t/QHTbxFfsCYQZEmzXouTxMuNfxOsamnosPtE0sNoBUaMpbbhx7l/v+GA4/ZB6qMl7bTO4Vc
bRVXkJ7NNFb8Gj6Urr0becxFsRka67fK+p42D5XtJZz5+R/5f0GcHGtojn64NwTzDqL38XMnHblW
q+swaeBuP0XUghcJoUiIb/ZrXbbXolGxI+nYwkJBzkZXZ67ItNE8+dv9cc8A1noxYTafS9qWLbKt
tLUtTxHpkEVt3lVEdGKb2QPW1aL+0ebEq/v8sTToQ2LbBtxgeBa89h4tipmzgyn+41Vg03yyjFNl
dcWQukhbbCbexfE5unvdSAk4gkelstxGJgNylBo+E1A23IrScV0ZtFxM5ExN/FRVGNmcl8ZHVP8j
PpAgcd1IlFk5WVVVXk6Ed5EDj3vmhjBDKyJonVbwMWili0WgNpZ7USWC9WIhUunNTm9rzn5URhJT
Trzok2JBi4w5py/2UMAXUiXMm9E1LEGs9DlRnOaNGMpBbc8bVsqmIl5TZ/YeFFuE1WYTpUeqoPeS
Sz8PszCOYH1BNQ+colSAgucK1XQAl/kVUE/k2Tucg3lIGI+I2740AMU7opDKR17w3e/gpF66LCXL
tnqU9KS1lmGY4zeXDzm4NJe8eZKxMvb6vHRzoGw1fzP5nTsmbijmvxrP+exOZ118lGueOk+STN9d
fOHDgVAT2jagE90wjsCY7Anl2hgFf0FcaCRBmtZVknbmWAHsyCnaoA7QvuBIUs8asTpXlE8EGpIf
bmMWfh0MDKYfsg2rZpz/vcorVYlyAnSc4L3tUBx2CvJo/DI/KAUxB+0pVGAv/FCHjVyux9qB6qe3
NofCqt4wTZXLt5yqoXylW8ssht1aJeCuUC+JETasp+ns6TzTjeMwh1BAi+4QMiWIO7qYV7LqDtAH
6yuAEFYt2a8mdpWU3QkWt2Z1X83iEOwVsi6H436DSIEm6LYPG9frvuY3C8+zwXOpmAlB6w982xlT
5aTQ2hmddFpFsQ8zHbKlPIdzwUJaBV1G5KlxI6oCKmIbe/h3RGXfiJMDV6PbAvHllz4YYMTSBpTY
WRzzl+W8ZtoQV55CZ24CJhPyA5cpwdv4FrN9xwRy45qMJjAmwBNgxArydbKh3leQzKn2HJfVH3M6
MJG2NCWliuejLuQrMNY2za8IgCpF2EzzY+muCyaONKCXlU8BDg99eu4n/BmCG4Nb4wBKKIHePjR8
8x4wUY8QR4IdFusXd9xBYcLkm35whACaQkKJlKo27yhQ35A1qCYMDqV6qAmZ254N6itlHhIThHcN
Ig5FZD8+rtVM0H3SP/I3TV3Megcvmb8Du8DHb2aK+rhsOGZQTJ68Fd7qkwAoIDkTxaZOt62+x/Pd
XMphqxwLPVgAcFteOs6zfAyCf3qUClgfHqNfTEbEySPxcRb6SQM9ADeMwvobOA8Pq8vBAp3EA9wq
6/yl3QGopET2amG+oNH0IFXejvTQaKJnALWWEiuUwNEbFa5LXrG/LA0kxuRNAHCWgBVw9/FH+L3Z
e7PiCagekPhShYekOEyw8Z4cFQu/fIBnR+LnIDUA5/vZsa/RseJOWIRMJCAVg0k0Kt7pA0NoROmJ
g16/Xz5eYLI3wT/J+bC76dbi9bua56hdqqFbr1k05mx7wg3UIXaoCNeO6Te7VrkSGkvSB+S72CE6
oPLPDvYNJppFHdnv7QcA4Kx6zyPs+O5HifIg5tZzU3/qIfwQALH0WUmr55fAfy/uBsLaacN6dghs
6KxcikUtTtHPRQQL776wQCQPoAjtpPGUrIt6wFkeholhOAHTCkl2k1I/1mmMx0Ge8riIPDaFiKWt
H/UK7tGxWTqf+F4d2wtKV7DzbzhfWkD6r5w2sDfdoYDmau9qO6qtABLYwvU7ByQIAoIgDmTxn5ZI
oHGCo9xHExZw8t6/Qt/8b6jp6ic+VPP4YPpKpVOov1d2OsF8lKPpueDX8KXQn/jwRGdNfa5DQVY/
PdJMfQmp6RLRnsb7lKrtXlqAa4hD34Ay5NtWBGe3WLFBBOmca+arEy6sBcdPP1F8xtIJkkWnpoUI
nCUkChQHEbdS1BIe9N/hVEPnl5wi8EfszMk+KCMeT0QfMd/ifjcAWFbLcIo1IJxIIuRRI9z1Odzh
1effXfQruVK7QgFDIg9U9Ud20bQFAPGpb+iNiwiYFsg4pGTTWTRIU5U3G15aYDt3wE+aRuh/sKwL
uUYMoFZKNLiF5/TLlgdAyi7Wx25AMVqX9SEk1UXgZWRQV9/CyEw3qxCq0iSNHNB0GXM1o9Hxfgwe
JjvKB1EuEtoY04Qyh2OONJLHP9JG2x312uyUbnBY7MxwrF6PH7Pjq/Ep3ZYYXErsbsJCYVV15R1S
2mpFwDvxFW/UwaTZWkeQrzxRERbPYVLKgcyngIr0mKgD5hTLXeC4/gpqmcqj7/bfGnU76UCBFsOD
+lmhCSo2yMK4VEsuafojo6iyrzhYKDp/sMrq+2lTXqh37sRjLxb6a6SSRl5EeVQCQSIzcKrQlTFO
NkyJJtxBk/IYYw9+RnIWHcYb1c8BhoOl3UmQ9IWDhNAQTxBHFnE6OcF67I2tXKO9gVRy9TGX9RAe
/bTNpBMy2CbrRK6IwotmE4/Mkd7BERk8Owkdxu8d0F521jFGkD8d5Il43Wk9cDlgUuZmx+k7r5Fj
WKtXestcs6ynfUhORzhsXnGKSPdcYtdoRt2c+bwas9UnO+yVf1PyeGgemsaxBf6s1KTr2Tx6Jyvr
SxiVA7j6tOQDhoNmrqEdYLWZQ/981dzyJ4ZF6O8TWHwzap+eJIIP3AfsEz9YMic/mhvKFBjb98z5
et/1g9YdSv+g0h5KrrnQ1uE/ZHO6BVt3DeH1wYAxYqh0Yg83Kw4Ndsw0Vonv/7IehKrEKgOLOOxt
wkwggfRYVyJL6whltst8acu25dpPrfLS9Twh8qrROALN9zn6SOlKlUbIBHHF/Xydu7EuRmAsu/eH
yj3TNPLVqWwO5AWlCyO34/+aMgefZzaByEKmmyjcUosQcREjUV36GahYj2BWKb6Zeu4hKp9whtO9
pLwdvAr1nVnF7V9Iz6abD/rQ+1RAdo5wZvGVQ1OhR/YDABklYg31qdJqKuSfM4T7QdugEXafIqfg
p03McEyGDrLbrrjU7DtrcCS8HvlSu40XWvzt81tWeK9ZE3cyaJWpGYMo0fN9j3Fzd7if6KhnxcKA
el6Rk4HKrRkLwQ0hFhKvGrdISgCMuEvaaWuWi9/7AanyUXE5PHH27WVvUZbZZVEmvOMJiwsrgZNI
+p1zXZXJWB80U8hxfJLusthZ2/tteKbJbnwhzTJ6az8L1po0DSGPazhW3p3ZaKROLwVIdrL0Hpym
hXQUbe3SQjTaw6F2El4yi5UEcSRkn+1fImEy2Y1d1K64zWcEloEnals1ODJEBOSp1g64BYyYJje9
T80cqGq6PPe+V3HUrAlFtw93m2Gigm5q6lA7YRt1FwUUDm8rbchhOOT/AC//m1TiRrHbzudItxiF
d7+X+hfKIcGoi6mHVcM4DKah7BRx6oU3T0HUNcjGJ98SAiXSYJi76pvXVjDyjGgbha+3p5xYy70t
a402W0/drdGt1OYX9p+48cTRhZ4g84+iHe2UWJTd93yzqILlP3ahpfGKeNpsoUPlshS+f00TU3b6
zRy4DzPdXDPs+mCY+5l/I1XXxzoBF/2cB4Qj8q+ahEL+Q8j8j2MBBTJvvSTIn2/p3yx/knJ7tKua
lHzsNzMIZ/NCmbL1tdQ/1VAKMVTn9d74PYNTBAdeyv1RYKvzhy2Ar44QlI6Anj9/wcTlRoqXYV0R
VdbMMSVdCfDe/84a0pEFVo8mtO+vOIA8bVmhmFR/SORpPTpWcT3nhyiK4rXK2UUl3NzZw3FYyu2N
zpnQaBhMvlQ9+DrDShVcn8oVXMjmYvyxPWzwT+5bkxHCgjaZ0ztj3mUfEdhDPcYQoQlDbKsf7A5y
9pEK6wd6IKPR4E+BGbKZOsH5mak8iCPNWVCaf0VmnmL6OUhr8e8l/JWWnmRUbYd7qpmfrL8xuE7g
AjuzrcyoctZYPF9wcGsK6b5jJt1XdtXiCQeswmQTJEZoOax86bJfNwljmdZ/ltX/Uiun1PUjZ1+L
9KCDq/4U+H+8H198B+0tFA4cJs2PL644wW3EDQgyypug6PoU3tbcGBEViLNHSiQXRFHYMafweevf
AuXKFTROrv0d2ElW2R76PL3OeVftDeE2hMlZ+aHMGr3uJv4vaxvcg8Qd+fNxYQ/V89FXbxbIdl/y
rkPCN0MXsjdwyG5kFerNdL+VQPwOHpQgIGx0oft1w0aRnZ8RjnxO2u0pa3J8x8AeBCYFgO/JZfaI
U0o94TfLmWT+c+J9YWjKBWCVOSiWCisuMTdubXCqprArWL+kTx05oiv05X+/sAdo7PQufKuq0e75
7A2EmH6l9+CNx5EXHnbrFimcj7+b95dPzsiCUXqlXuYQ2S+xCgVA36bgZg/fxy9WUepaO23gwsMf
+kSMzafFFwQHd8V4UEPLXdHuUNhGN06WHglkaMDHv7jp8+BHHBlvh/LdtFKUQNu1t1jhKAHo6bNp
/w1zblcdO2YDMwV102cO0SzuIKs1Z+IooghUEE7pu8hoUgSeRhxZcThA/0x8uLOPPGtEj39mtw6I
6vTwhqVgMkKQ4QP1bMBubSiHDb0RLulCJNX9eqAf8XsNTvFfuEMboV/sPF+R2jzp0orAQ1qKtjo0
Iku+gXNo9nEuaNEUTudhyTDO/Q9jdLfZvB13jSp9PkNZdIG/5zbbNlh7JcPLOfNtuuuxf3dRM0Wx
fm4jHe9aHNRXIdZp/KWBb1CBEwLqLABOEJO29VTI8ygJKUIsBtqUPZEjI27yN2ldCqvufjqBui+G
4L3RH+ELsENpAhlxPkGzZUiKD1DV5P+yS7rvtpYB6sRMpUaHPBLidbyccqXcc1zQdyPoY86gzZa7
TInujrB80nGroZouwICt3EPYkXnnWFx3Ukeh6W8rz4+oD/KeBw63qOaq4AFmDpMZMZ/SZlvf5rtY
HNF5xDtvo7097muBigaGZdyghStKvNohhWxLeBeDJtV68LKpa8sbCx3gQ5bNkEy280APGmTFsOtp
0Slo70Pb3ycuUQB8WfRzMFjxZllhAGwh7brQKpMYqsY0uMMOQ9dItJl6vVCQiibV3cjrWhg2c0Lp
eGEMK4Af1xzNijkYEEVqTzkS7EJ8uQSphVAcld/fYWmQ9oX6e+2Zf7PzL5eNiuIMphMgF0xbUDhT
cFf5Z1Sa6lIxIaNY5GbpRwQoE4MYd3TwmP70sBs9rNpQ5u7E/m1NfRri8hxwl93AVv333KawoLxN
4Q6BjaHT44jl3qroF3QyaXPbczqqxbLROYb8tDPxEmhytnFv0FgQnR8wv0JGvSQe7xp6OUdNnpri
IW+ksxVQfJ7MvHqHRnuLz9SHCjj8HtCOcRo4I444aOAGzM6dW6Cud7qU46RxRkwxCV0myCJ4AcBG
Wt1tRaBXRed2aKgEH8JMp+dxTJOhJuf2sc28rmnfuJVKUxnWHrAVuZ3lrXMx+ZGoE2ABRuxPATEP
cDfE4fTlP4zflioD3Pg75lXJ8PMCiYqXJxFnXghjI9sPODM1SCgwwbWxFA4Paks8+WStBQ3XSgmh
DHtUyWOR5CGFGU03SOHkwCUONHMaYcjORhyLgwTtAesdqq3BfVnRMvM3lcgr95W6k/IackskUF8P
SLOm/ZyFqQZChe4GLqkYzA2EQZ/3sssqwHlykTHiqIIqr7rhnyddjzCOkPjW9f5foBSOwqVfHzNY
69Db+xYAI+VOWYX41AwbwTZ9ghnv9hCvAdvzUtjJgsAoD5yp7FCm+ZU4pAtSPKREncs4cwsvdS31
rliKvXjd0uTF0X8+VZVFyBQtQNKdKCPiVzWkget7xcbis7Cz6zGOU3DpFiQXMIvHta31QdUhFqIi
oAspBlyBBu+w4UO23RQAszsnG4NUmYjwCEDSUsTQyHeZnbYDgnYnukBZcZJ6AWHEQ3cBOTKxwB9Y
IKv7Kz5oeWRT6b9zyqn8ATIVfOR3R/gDqGPnM7odsiy4OqHbIuM0clX/x1jRV2RDfvSwhrPg2Jzo
lpSTTFmj7RLGz1nD/udMSPiG7B3vaTyU0Sq+hnHO9hUyZnLvLzxGH9Ftbv5xNhlMT0YdTpYpO7e4
MGrFpa2ZOhmOcNZvpRyoDMtLsPR+NvSOPDiSQo4XvTTOinUFGTZW88iIIL2kipPoxNjuhIAwrulh
peEeTU+SWxyfvU+2P+ynNSMnW+T6gPug10BltBvsiAljbKd+EfuYkCILHsjb6qAi6HchC7PS7K+k
r72klheqIbW3DJILPFfMbaBMWfQiCrSs07gPNmw2v82IbbrMMhXfRt/z13jfoFiCODTQ9mXLLBRV
RCL/nr+2QqWRpdHw3DkRQUlLJw3YQDoUaX4teMvsXRz0NnDFYLpaCQVNMYPc17N2w8VTdhPXutl0
jSqYl5qv4qrD6hzd0q1dZ9EUX/6sO+FL0mwt0gPBrPORl4FNNZglEIzPnNIwMHEnhEYZv/WIl6xh
0Y8+mLjKyTHC75423kWvjnrPXAIugspfOZ/G/aG7mxV7tAPxFP7lstREufbfACOEGimiKlbWK4xy
RG/B/Q1yNr9/YcxOQ2OnK/F+mDxLMPoD+rXH5U2y10EmURZpEsPA0I36j78QyHgtXwcFzF+Oax7e
Y3aS6zeLkW9DMhE3RKyUckRLHo52MKv9Gc6eitTO05sMA10XHv0ZTspUVd+FgSgu/DkMBEHmKgVO
gydzSJvuW9AHgZa94T8quclDM8NNZKgApNtCE77MGMkKB2VGyRql68GLGXDwIupi3JNS3RAELoaP
w1OITctQukQ4cC2qQny+HIlu1Yu9RjwThXTDSmxDNdYxOa+JApJ91zO/hUzm+XDpeXPF+ZSTiHGs
nwKPdelp38Xbi1Bjz7nDrBW0AKXpPoq1nW3Z8zerplKf7d8SozfiMpPRgnsfJR63estPeg6wa2Bt
ltfXQ3Mv14uuqWcuDIydm7SxOd+47fa7E6UgcwGQqPbyluwCVbmcIjLMkzR48JVtclQtskKCKIH6
+DH4tdZUxOF9rXIYwB2K6eOXLfqASfCg1PMf1kZGOfNCERSTj26j76vVpZg7ytQ2A7cKcNM8HJiT
gXlsVMZx734gNYTHWRK6xS3S3M4MuJO4y7rQTksXknknCqyDasBVBvn+jzS+DJz/fkPoI5wR0/wi
+sIczQIHFnL6IxHEZf6JbOCDhzW6uE+Uhkl5bdTEIPZbyuMR+tQY50y9Lije81RsgzIRoRA/eBy6
8P0HNY55W3jfDkSCmjHmpnUDx49+nOrK+Og4Q0o5mzmhEdi3ntRnBn0vsjv84SCHFLvsfO3ltTg9
7/WWEj9RN/z/UBV2AQyyrcrhL+kETuYqNn53NW6mcCar+Hpwzc2RSO+XYQHHJV9JY0RfkHnXT1nR
28G7zOehADoflSZZ/fvxTkkStx1QfU6hXr8xBapsouL0Dknilmj+GRBnXNAfCrLlvwsWOlrheqLC
ycPn/Fx73MC99PpdoDSKryzM+96Pu1RpAC7K2PH+CDYkrCa3HxNP4e4RaySxWjh7DE7XycckPKRi
nIi6JgoVTaLvLNF/f77nSsNi6UDJvRetTV+uzYTW4s9imVIVgIuHZgKTQhtpRgRLXZpDAttEijrY
bmrrmUghReUS0zyr42BVi6eiD+RBGbe6RobSUtOkzlOCs7sTOaJyExaNGYavzGYJtLP1OIvyaNSa
PIohApBDykDuk/LGGuRrxJ62y98D7IFhlK25nMIuDLL3jKnolavO9UglFEezaEodxFuKibcEeOOy
7IFJ1XYjQ82EtDByJICc4uGaznUhwKETJOiX7lJNRlSS66f2z7VH4k2UKjywZtCQzj4BTqUojaXe
anN4qF1h4VzEKCDB9n/L+WGgEsgA3sUnSMNE6ZL8F6bjyqFq6sqPOYX2G/by9wjKOOgyuDw/0tmN
f4At2B7TqvLF06dqq1Whws10st0BSHHMf1gvg/vZmDM0SQ5JHrZfsnN7o1rTjySMkw1ln5/Obebi
VUKeRQRb8fuUjA3AZlZc8/WkH9ogAYBBEvp4+QR1Jd+undCSR5ofnuJPPhd6vtSOnhBLIRAUPjXB
/jK2N1ZR35eAxp/bm0yT7dBQZicxEjO6EhLW/DU8IFQkkp4aWb9q9C1hBvhBcJoGASyfq86bqX0l
YVKg612tBTtEvJ4OWQ5Dl+9aI//bgmb4P2a/dgPD27weq7VSu3HXkDJB6O8pnfg2h2un6FeY5LB3
wpUgxQIDkJJbLY7ERuV5Mt9wCRYu0gY7D1OZO9TgfX6ym9QKEVAdlaTM4Fw1zevSlCuZOVQhc5OY
kJEFKOVUOvGzsShUMKEDea23O7wpRHRZeNT/VNEascNzjYZ4pNVZx0L3hjTAwReeGn/HwqVzyhMR
YoHk7b+Cu2wlUoYPluBgh6IITfc4hRt9HOfw0v5v6dyIkYjyW+sOmtrsi8o5ZNqjL9Ho6bWyk0vs
EhiHJRxkb67ljFaCGqWYxUD1LWi0DYw4w6egOChRMvLNwE5kxiGfK6lXhextIjw1m1HQqco6+qjf
PFa8QLP+x5Y4aqqF6b/sxP7za1ib6Ffb53LJ/vC8KiBkGBmKeX0KwfJToOxpm6xDvKJoe25y55zF
A775eW6Dgl0XgE7z7dfdjPxJTYZadDwKTWhCdb8sELGT5FmGuQyKtULT2G/OtzTTGPLlfXZPVr7e
dSGVt8+MzgPz8MyvNNYExiZUwipipflR5edsK7e+bgEyjSxANzPN5NPD3sma7/OHEhDZvFAYqYP9
mmmnswLSYSP/dtB1KY9c7QlwkUdnfC5x+hmr8csVZPwxL4+N0xz6cygbp9tU6Dx8V7deS+5pDid/
NM81KjwIL0GfQ6xL76j+6tDxK0+WecbL3oDI/huxE8BpE9ZysQv4YAqluoGsE/68Htp16bMfsND0
1POkgMEOr+o7zpIgRoXm1BsyHqASqLZSnsflxzR/AHb3Gw4vv29l+AcIZDjcTFRV7pIJJ6EReTwP
wNHX+mnMzHpDdXbrD9mf797yOZwlrD07TKb9KIYe5L+Xtv8rdtD3FE35GEDN+hROsuymLwUVZiCw
6E/9iFQgtSilJhFA/B89/oPiX5VdErLErVDIYTMbq1A2vN1AYLV5amDEdziABlA8dO7TVDLGpFfl
YsJGapLb7oAvJDuCBAXa+NmRC4qLozLvQNIozZzBwNxbqZKLQj4lQ6jDKaLkRtpdes1Ebcxg+sje
mpV26NuXlTyKUVAQM1SJfRr60oj8GyIkyLVTcVCeTDsrrBTZlTh2U4ftGUsg4piJXuOtV9tOVdqb
7COC+EfTHh0zPVsN+p9Y2LFJACBEH6VhNYo9g0I0rV0s2VZW6kMxiArgr3Ynjy9Xz76zYFNc/fDM
bdZs6hPZnCr0BMExaapVMldOjPusVgc9yyez+g/QVINwobdmXTHCT0ecwPN9TlY9Osk2KBY7WjYp
xOM//QfKR4RXjBfM3tYbVSkCE1ZYE5FOvljtVkq2YK79Xpzd+NKiFhFyPzarpXy/pcFbewlJUOQT
4j/gFnOJyt44VdjWJQesc3h/OdT/6qEEpB3mBiDgQI4ePAsIqUPstkHAHXTU6WvP3U00RUS8ZPmk
kY8H6Uw2nJ98um1bAtW5wwDPT0+AKYjDBNGfBi0UbLBUKBshopkkdXZ/NdHLdAQN4F9G0B/fnsaF
rKzAHMix/nDRS0e9BTyPjiqQlpgEbAy1SMvhRY7im3NUbcYJJD3gtJ0TO1qoKDJPlyEMYNNvkcZJ
9wqiKZnNs7vbXEhAO/7iGeHNYLa+Lt0i2S/zvgXqMMSYNOL5ayKiiqIZD0JZ5TcuQlG8Kw+Zinxf
2q60jvXOZAV8m15KyozRC7KHlici7BedD/3NMeilP8jqzgpCeMrz2SfrOa8LKwEMrbvePpZdredJ
ckNqm5Vq9GDKhll6zUax1I3MAEDtkUlNw3PH5naVLEvpv0f0BqRr2PlMhvPt+25W0am64XGPsyO2
EDyIVEiMtBwtnqXnZPONo08AyZ7aZLIZAzPWpvXRs52fM+oKWPab9nDz1G8rylcZ67fWYdKNiozQ
/EjTDXOlt4X3WDknqDyL3BrHM90WJMuw50UtLw9sQH1/PmyIao69mzuxCt0fTzz7SLldboWdb3kP
p8Wor73DHhLXhddusNcPxgRdkxuxp2BojPK61OZ3LC7lB4wbH4QrotvaS/Ays9tc3pMgRi/9ZBbN
qnUiT7YT1+oIJ9RzggVMicyYT8lY/cvAFcKlHpfY3By+YDAjvxKEVmliEhka1Q5g9DSub5wFh7g5
wJk6vNhf2D/RGzhhrjuHUpbgzWBYh4WghXAmaQYdgdQ4AvjNrbtn8fR0C1/TxeSW0ta/+JtK0Hku
tHMCRxHreoe6wzo3ICuR79tj1B6tVoOhmVo6SEdiLDOsfE0jmymYm0xhPvV1RA/RZ0EnXC5r6Sdr
e7pJQwwVtVhGWob9JjdSBn+WAG+8LLCOo2u5fH1lBI8ZpKaneaucEcjSDFVcdauZvfRS7L+ESEs4
m6IWJRFT6UsnSmKpMLUNUyHMOs2h9/iLooKj5X4Ad7NMr3zApbFY7OSCfQXDflx+Af/W6Sudo0D2
gUUeA56q2S0m8jjEHhzBZnI5Viy0IMMpPX3wK+lUn7clEa6pQoffvV1bXukVB/hIvtPwkvX48Jvs
XxpYbzoEFBUn79UeoyHHf+xEFId9BU89+ywmg2xlU8aEIk/8QzKyoixSOy5YI9/Yez6fR9NWwJEi
XjzdW2Tc/SThOdnORaKhY6TYYWKSuzTYckaV46moHsxtHmbjp/RXZ0YJDXqbWFSjnGzDNE8nFWIT
/k0sARIxpktWmwa5rHM2aVWq9AawIaBMWR4dtzdSHjRWhr68hA/qki+DF/liSdGahwtNKBcAdVem
0F4sRxAcnfQAkNOdtFhNxaXAsQPM7Bnv/2E9ty+8lk4bv//ewgnEswbTkzeGAvfHxl63GFV+N8jl
/w/Jw82Ti6Eofypjj0uqzgCys6NFE44OhvaqXpHB8T/CLYANUeiNKiVHBO3OOHdNKrmCBAMTOZ91
47cV3jOKn4bE1fGY9AUSJgIOHpnrc8AwackuA/xcd4CWe4iR7sOnVb0pjCSel2JOa2IBBhM5ggEz
r7tV+MxdzVCUQ9VHk0gnA7eke+mB4fAAk5JJ6dzi01DGIckwOyR0lZa+L3i84IJgUtTRyPorUtw9
DQWPyS7qU1pV4APdUELUoWHafU6cgm7SwVKPxBxwg6mhbRPENNCQ+jtgQ+HQeFn88WENROgdE9W2
jeCkqWB8uB+MixaVqPkVR22fY59wej4JeWdRcM8sHoQV6kVKGF4tQqbXIzQReLjjdllE70z+/iId
tNiwWkuqk8XvEH7FvfnphbPFu3Vncu2mRsGRTa54yZYVPdZijVasMnl7ruodR0wMoyBzsA22lUq6
rqCxgBPni1FlNyRr3u1AY41Tl8zWmpyD9cCl//0CXEWZy47Ca8X2JQBj7Ga4mMeH/Iv8+cC+zm+j
8+4VA/pMCRbAckHdSuuxMV/4mlo148RZ396YeQtCXVh1R9FzJpHxTFEpgl6tb8AaLuFF2s+rcqzu
hDqwPFzSjEz00wfKvrLcyuNWGhkYLdPv9BECvrXAuTFW7DMmBOqcXkNzTAOEnFXOOj0/c7V2cMxC
CMV1dSpjtxBGHKTPj/jkfER7nBr5+tUuMod4Hb+rsEoHL6ZnCjV9oMdAGgbRWmpGlqVePhhB+Mrl
ndpwwNJnE17JNm4nJhkF8/kEnjAt0xRZyGn6VswNvF+0/uijC6Gp41d2DRe8yyC6hPvTYlgut/gC
746drSOenGtyKgb2IDDPpGCzHZe/beBN8dsFJfO0JtDAukdBjBEJbGV3j0FnVTx1avROJ5d7xPcl
XZ+rEVJBTAj51bB9+vCHN85kJ5wX5mC13q7+OIQ0/7UxlT/A5ISKlBV8t9FDWwvAjZQMpP/CplXj
gFFiBHicvWqR/+ZV3cB8VEEy44Evw8fNcn42HrWnY3a1Ot+VfFuh2enP3QNEtxRjR/H4e0ueTZXZ
9mmWy7Ym/GRSQ07Kok4hj6lqP/21hwfpwi2WVyjs/VgqfVAq+XOIz3cWixeHVvvWR2aSFrI/7qfi
JNpKs62KoLx8r5YD2ih8ye8IbOg1ub2R0NPe4lH/QAytPiGtPZnk/q3RHULjwgzuVEtNWRGFNEYC
9iiH04b0nWkcldYUAQFtSRTnVdonKZFkvXOtGWX9EqdBqlD3z/uoWqx4/GuDR+wUmHuzByUeIu1d
2y94dD77hERhQO3GpDf4VWqWvK5Jqlvdq4EJcchjeOvgp7hCEG4xEUdYFjd+mYbWSO/ZrL22PgW9
a09+IPjELRJQ7RCsYUHugzu0nJ7iJzG2EzIPrGl6f3Z6z072dxlwLy+xNyCWzT3gypIIvfvkh++Y
oSfiDrIVWJBXJoe8cBO5czioLFw2xssQ5C7nHMmqOyPeuHatNJqpNNGyT36HGSHgA/Qczu6AlETk
5+HOxWpnDfTnidBtxKLrXHp0lriPiefVEFnjWchsOX9DL+pSObV+f2ko0jtxzXvfjgfvqB7Dgn0U
Sk0DjNtWPK0EyEvd22Pr2gRe/kpS2Tfk7MfpcNELx1X9tWKxeUZZ51zk05qf6p4rApu2422r6+X6
BAj1J463fIaVbXh3Deyl+dYn1RLfRNSGLZy0Mj7xGCI9m3MoFY6eY3j8EtrBqkySEqjU/jw+FSqa
weDRz2ZT0jb9K4Fa+vxZFGUiM2KyOApmQOyGCU/vcE1/mpf6D+JqjXJaVBo4Tj1KjNeBhMW2CojN
6g8PtRGv4H+a2g3qT+lovpxjQC0P4w+8mkn9kKj0LcLu3S00ciMRcpvinbkbtWbgeDEZdaF1+NoF
ygXg59qdL6g/nHndx/KUcM1g344qkyxx+oIN4JVLJE1y2vWuEVYw2FAaCTZKl1p8h7OA4bX9autU
Cjs6lsfoPrYt5EbUnx5HCTZhfP1XUyVvfU/gVPP3JleC3vF+yHClalWQGgumZEfRma1slF5d3NKn
P6bue+UiTeJyV6/OgmwPWRa6EkYQX83PLnk/Chh0smhalbcsQrC+DXtbiWWbWeQMx1XyavkABQfY
+KEcloPQ6aWPrxOI3dj7eizbqUHUigDKa54XEVAJ8qlIsDMllvSd4PJ8InPrzUHujjwag+Teeo54
jN3wk8Wku9lHhc3ZDYzmskxLqYz+sJ7UETpTc/sx0V3bw1POJUYxmz5scHLefC13F88YokG0O6y8
T/uzaEMWntiPSMbFeFV1oHidReH41poHOZdj9Rlsk38Vev8sI5bZdTZKz8pKiquILg0WKP3VNlEh
9Pd39GPotHxmlHqg2X2pWoI8aveyTAxzEgTKFkvi/IlHbT2ffQd5iLAmeaPSJuR3Rq3I6JPn+THk
qNWpGv9TjAe46JMvz0Awm2hDPViTannIfGZZ8eSriN+KjPA4BP9rx0RnMvQihIRsGIg3W7K87ltf
ss8kOjY7bmfRfWRAb1EmqPY0T4vYzFtFpKXQFZSYvIPbXhzKYdET4brpuP+Zifgo2KF63DVLI9WA
8pyeJXzjD7iPAIXUw2mJFMtJu+I3K75meEKRdLbGaU2oQ6i6ieOH09RdtSpqjTeFw21zMuhJkkAf
t96JpnR1d8/iXwsiyXZYm4e8yeqbJY/2Sn8n/DjxLl+TjJinoKOza6fRBmIGxEoCwKkqbXagsLMY
5fPdXzV/+Tl5Ay0ExywAwj7VDIPH+UmYgAQGCChdQxoOW6YFqg2GRyYbRs2jvOHEF4t04jucrhrt
gEiNqSTXkmamkmjGifM4UI5j8/XVKRezxVsArJ3h8S+eRhHs9i2uNlj+m7LCGct3kJCcSfBzu62x
vSBO/IUlzFK8Diu30h2I9GMRhOfXbAIn8YhXik76PiNdp7LB8j0WPgrvSo3gCteb+OxoClx24E7q
xI48AjClsxLmQapvq9Wcja2lXsqR8jfmtzjgwO1jUAy/WELmu6D44+MAALCKGTOA3tsllhAiCpxu
ZatHM8YvL2Ortr/3PPLeLDsTO4imn62u6uBaY5cgbOP/xLeVEOmmRZWsixa0OTSPCcbEgxnuzfeF
GjCGFFRQp2He1DehF4iDrOM85qaYKchwjSCmGDFuI356Zy244qFgBFIfgnVrI7YS/NUpeKOpkTgC
Do2HmZvaso6SD0uJeAbd8SKK6Smb391sYYGOzR2q9aTL8AovevleIZBBdY6TFfC1YSoArWl9Jkp8
a0+tDGBJ0b+eIKrqXcOOC9LOi9A8AUe6Wpf8cyFauIJRj+T5CWld8oyr0ZbjZIEQw98hxGBfCVyN
h02TfgVwZui/UgoFzFhaox45/lC2pmEBQEP51nZmTFqn6reUkeaNBcpxsrKETb6aIWJQwdcV4oAX
Fb48xfma7bveen2ZeGZEZ7ftGQod2LaI7HECfBKS03DnTxuoF4i8Req0Ldpw1D77+10TAQDoc/Pe
34kR3o9eCREmChNleCKkEl+pBROH1UxN5rNBKL/B93DoKhO+1v6pOIAGAKthW9lJlab231M70U9D
1ov8EW3tNpzwf33IL0XrPrL0W7D6NFNAnmqntt1X/wlVbBqfVtuLDY6VE7PcjURVXwt3NNr8Uj+y
//ydl229MR01fmC26202FunOVjKxz/qWOq32cUiYVIwlECZmWcgmthvKcS/8Ai0ATwxqSW3pb8FQ
d+y0qy4SU7H8b4sPm7C7qytmHtT/swRF7huRrRfl4lsK0okrFtWJqRWN290kaKnWlFowv4lb/Oak
BSJXoUVcYaKRam1hNwOrez+Hvu5w6yi3NEaBhLHcUQR0OpITTP6v80AaYysS/8mtnfFlDELotjOx
W2YpdPXo6tpA6SHK5g6QBvwGYivxLY+11SpxQUCmWkoJ1kVm7uuX5ghhTR42SAVFAWKb0jmhKqjv
dcJGhBw7reY84oDxGE49sf/waAj4i1Cn3u7hAclJGobvHdB6TaAWLCdtSPhHL8Pj0GH+nxLXEiwA
VLzr39+QvE+GyR/aXccBLzaK0asDQUnBS0SpMCowOpAplNIWuNF2eTgxybkpIPl7lpkqUeeECF2j
ICVNrpMEUB4Ehf7pOT7NzKPpsAnOU+7gA4Kn0CnqlhqnKLXu38nY046EGmlSoa8gfeSSMDEInFgn
O3U0me7cb8qlpsq/qtpUUpzH7SlAhNY3TmibFGR74CK+a5KNVXRM9PqanP1ak1Tx1xEgDZKJLkGl
Dsn5u/SkKnbKUmb3+erax6YEw4P/8WEE0Yt5f4Ias7dbyTrsL28LH3vkZOKpj23E3FnYwKW7hM4D
8Pm+SX3QP/C6uFNcFGYBNFnhByfvbWD9FRkOv7cC9D1yXoDtDjJtLmPvyTx+RPyKc9vMV3h2R1o8
QbH/Ldc1v7g428FDuntgMB1+dX227ccMIOA1lcjiZsmK8M6gyQ/mYaOCrYdX9Kwv/5LSRhxRS8vc
R9Pgf3Qu7KCcMDNQBu0kS7ouq3xVBedfA/tIruhfJyfR55qsmjDiuWaCxio/GEZ4KFfCroxTKWYB
hWZv/w1eHKiYq58+vqm00btz2V0WGqZBWQPN8TrkCwy6j2M/imdS61I3OFiRGNfrLI4E7k2J05+s
aVpi2VvqmhQaUb1O8rr/zbbyFCrJHGqwNvYVOF7vfSUAEFpix1GO9OQQ4ut6V1Coxvit2cA0j9QE
hmYGNitJcWOZN3F/TaXq0e6h2/7SUOxHLz2q1/bskn6+Xr7YGkUFzEsmwco1LLleWDZcHBGj3ycH
Hadypz/8TBOlvZlthqjWliFJmOyMm8OvlzZb39L+hQ+VrTebb6dVi/gnJO/uiYiHMXx+zO7LrpoE
gsE7os4cWkAlA81Bvh6SM1XJEDYFrE1Y/CCcjN/8icBjHaNHp0Wx2XbzEhlXe9pLd0oegWK5Zhcf
WwKDdrYwp3sD1fDH+APBBIlzdEMM2FsAUOhzDuji74MXChSxGaZYdlBqQo15rfDuncv2BNMitWNo
Gdewkv1eIWFG5+IQApXuEDRWQ4w4IfSj2ml2n2jwLbnaZAwPwzFG8Q02a722BkuhkFeBkFtUNykM
GkOIOT9099tw9+VfDDil676NWweIl11O3rR1eeaTseoDgVOdz/UWEfDCiTFWh3e7GTAR7bIaifPD
lNogzcNmeqMqbBciTTef0Z17gwmVk6jc8tjZEaizZXlk/Ghr5Oc1d3Q/JfbJo92wetOx+Af1+sbt
LkRRfKxlvOs8CJ+ANcdngyBC2zMH2LefmT5dcZKUS2D3zjYpQqJskr7NF0hzDZMYc5XU5ZDH6qwR
sPjXqmB3jgyFkg/JiszlrGJE2u3IMxOwx1Ac9mprH1uEdwx6Lvd3IR3SP2SqxB9J9PPMTtFm67us
ceRd1LnpSJl5qDWUMkC1wEUtqYdFbKBBi937R/YPriJrOvstTlcH/7AmqKQQHt4Va3TxAlU4WuXU
SSENqnbBCuev9yM+yjp1NXWmAWkZPBvuPzSJYk39NZECft1cdCte8Ml2VO1jCVwdaDy7bNwoPs1H
oWoIf04oiolbVU9H7dyu5VCA2UxYp03x0rPC5eCisGyNXG32SOfvUW/szOcVwnP3oeh+6z55NyTs
D0PuX0fdSXyhEdhQ9itastzwhsycsIWHD7Jufy70HpIlTi48E03E87Tmy/Mev0Cm+P9Gxf5e05j9
3RMuFyVE7hnepbh0B5+iGBt8FHLtDbAErMhCllw5U1WGJXWLQP79akGhXPJPL/z0I/WEhqO0QFvq
OS+iKriNTochhArnkucE+hHvR+F5sWwGVeVIpLEmV5Pt2tHkXdzb8HFjYd48kkkR4H+KxxIQ55QM
q5ZdErFzErlajyk+N3YdhsoXu+EntfmNFvJbGsTYr4Dl/YSmXqo9iqpmzcKGlYKZHZM7CcypdAs7
TGQ4GDYEH6p0wNwnaqPrGhKNolnmIl3umBHGA/o7YqAjYKp4rjblPKNcRehBOmx+GMXCo0yWiUU7
EqKe1GcR4Khct+DWmBXO6ZPNjdg/v5sjFQH1RZvJov004zWlYuBBGK1WXVFaugjrF4kXR8S2rPjQ
g+pD1ID2PkcjA1Qbnp9NoFPmgSqpglYGlOJappDYtluvwt54bnl+NtNAh14TS6wJLdFwbc/iQEJa
NDVh+IEin08SzPMfdbn5P9stY6XaBkmrDWxL1Y6ouTOnoWkH8gj7h79n41ePPocbusj0CPy+sTLE
yH0Du+Xi2SF6aYQDS9R74vYEiwe1U1jvBc06fflldUotxlDQNBO2CdTymdiZJD1JzmG3YoFPHV26
wsY3R+giLZ6Cgu9YFEly6yUa+CSrxfFImSwbM+8Jf0Jv1mrMefeDD8bvU7rXzf2irt6pW8aeaq1e
kA6TlKSbqmoe6Kp6X2RxtwMoIZuR0ZZsXA7SepFSX+mi+5vJnflNrBCkS9sJKUa8No3bFmvAJ0yX
R72r5GG+5Yl3gdlwwyyH9UvjBUtESh6Ou//RtOmWRBB59ZG+uVSWonTKZbK/mgubU6RmAofW7ba/
pi7REh8HJwrILZDhfmy8qXqomTLMHJ5MdX5hVYdg091BX5DAnlS9+meFHsCTXRGLdOxDk8mSvpN9
JCnmbX47bgVFp8fVEYxSlnwFaXHzlxaUw/gkIyhWfQlNZdRP/6lxY/EUH5sGo4opmNtTuJpELbx5
wpAIqhTBKFzxbqUVgYtIHgVqLeO9MEwYp+i5lzIMxavqeAYeEEka6G92cnTovOTt8pxSgqW2wbTI
DEhw5ChVCQiXmeir2MwTgijTCv5nCeAvMJJcMAGXhI4H5U1UkRkiJqW61V6PwF+FO0P5O7l0Ygm4
512qlCEQ748dERqcHCdS+5a3THgVkA16MkxTLjbeKVq2aDR6tyrqg5mlW4Wt2EqlBkPTjbdL8iub
5gdGkBo0C/rpUQqs0mD9rQ8wCA62ssEJDdoVxDCC3xRm015tF8eO7gW2RA20Soz+oWiDvBETkPJ1
Hi7WoEp++dxyZYI1QaMTB8jtAhE9klwQJzvRBUWjCN5ZKzkt9i79ykDssqEabU1X9vJEihommzzo
T37Dfh85+YuZK1YWlRVOr1f77ON5VXfP3/LOXcCN3yy07KHcDQved9wd0JZg5VpmXlIxIjylH5vG
8o8gCozge+FoEi2FpvYqiVvPpzhZ44jxyNFNMTIO2ilyauHTsT8/cq14weyfeqDn8gIQO9ZFCH3I
mmk8mtiQz3PAst/bXMsYF3KCGvbP8eXig4KoKvTpixGGRQ/Mhqvn1PwU0Eg/lgfRLgk3J8H+NsXf
HdxEgm0a+xePYTdkkavuZYp27ijA2xzaiD7wvR1zd4lN1nD9N/N4lw+AZgzWT65l1VPhOMjkv7wF
elwwG2Sdn4Hsbw6Zez3FgGWkkaxY1QzEa/q/nswoElhY5ONHv0r2ymA7y06Qb9XaRkoyJG+HmvBT
mmi+Y55VIEisXCh2EmzYWmqFBNigFMvwLVwW1VuGae3xLJ6nI6eLF6lH1PH4+WxLtBHwh8tvYXXI
WSAABUCOapb69gRhBr6Kj+VsqXtbgKIqnqqXQdlBIwgMaDlLTnSk14SW/wn4z8bLVIELjwK6eQK8
rwCZQ/9tlVod3XRbPMbmBAP6cDkKPjsUS6qrLby9Uf3VSpEmgaEcSuzuGaG+JuWVPYgspxtQTQPK
6DFwKlTRBsSJ3wObab317X/Cuff9oVhxhT58mCMBES2zA/N2kUdt+fA9PprHPQJJc0TBC7FYy9Qd
EAzegF0XMG3ClLGi+Ez+GT9uHnFs8ALj2s3HKP0GrOdAxx43DQxb9b27lG2SmxEDa3JMHvfvgSIU
YDsPaeyD+fXF47DUso8FmQ/MltTHxeHM0lH9t3pzmSMk5JUElGeLGVky24/OXJsvElsbVFgIbSDP
nUITm2KVvy6TES08mSWPJUy+//otKyNGLwkpIIY1l1J70l1bCCiCQ0a7pQUB9BMaOiXYFpuPBkNM
6ZtCINMZ6iNuaQ4a/P4AOuuglgc4Ao16g8WJ8Gp4bw2jdMNj6JoQkF0QG7TPlJIFPD2m9/EBgOkb
fIC/rCqD9nr9dql5K6vtas5gLKBtnS5YX4F/DkmpZoAkhq+RIATGjFIveiNtW4HZJ7dCcD0CSJv9
SwLmscPoTmOA/IgCIGEfFV7VFKtasmvNYkv7Cu/qQmkJJ0RP8cXJY0NjriqGlS8xftk95Mj+oBj/
Uyyhw99kAtaNEjiL00tL9XokIiRO0cFJjzFYVT5LYc5xLmysjQqU+fvO0HsU1npapTEs/6G0vdkm
ktcXZ6CmoabLMSDQWWnc9ADO5eU+r5CFcaLuZZOW3xqsnHLYEcB0NMC96GAGPwVVW2R5RMVef/1D
WdBwvPHN5RF4vsEm0eSLPTpWVlAw9BAYRoIDzV1Bp5Mf6GU/TJ2q03nTNThzx9RnHEdB4gV16J55
CG805ZKIpqxgxbeyb0qZ3K0e+QuJXIyYFl8Ws/OxDSjJlEOnPSlxfDVELrgb2I1xb7B5QdmiZjqG
IW2qVrFRFiIgff+HEE1RystN3xiSKwr9U2UULtp04l3cGsCgevGAg4kFuIgNnoTGoiOTft8Cdx16
iYyqTUBOuf5d9Br4OF9usSObCSZ2DgehEZ8BLoQ2w6UemqnRzkvSCt5GW+BMPVYj8OTmj0Agp5U+
ir+v0mYdQ8obZAdNgFLjo4tdfjxGHW9HqyAC1qCmFJ7LOHlzWsCJmTnww6Nqce/AP5QrYSp/JzWd
xnRFRVg+iQOnA532H46hplfExfSnuSks256mirwrVkWs3kN6MPMbZNQFOIrHHflm+FnetWkzmDMq
SPTBHUyKEzz0RuLLeEKdW1E0CG2rnOlvxSsuSImUkR3qrr+cBolzyUV5twaVEp2HnQJdTtW3k+SY
PlGk4EFN+RfDWwWLbosJR4e2Xx+ZQIyUZ+mVfhU+yM+5jWFv5Sf3xW1ExlN00e+rSLsztjgMijuY
tDRE2lSMr+sv6PT18MxJFKdhM5//bW4lTigyJVd0hbhYa11pbreB7UniiwGw48EwkszF8feRybPx
OObnWG8DrOJcnHC85iu2gtEg1EB/cs1vho9qug+MPYwEGYkFPBzHb2llnPVe6EHi/HN7LpvzcZee
s+/Wn3hjIWnEhlIWeRejNOhXsn5JlfA7Cw/gqUtyyx3/JRghc1Q8bsZG5cm/6oeV0Q25/VxAhhPK
L9Fn5BBptx+rGM+kA0DCowbdoZ3KvjtVFoaCywWu+Wc0OY2wvYHOcoWwLlzrPSPNRPmFqSck1igk
hAaVK/RYBMbSVgNs6JssXEYVXk3VUVdESatzH+DU0xEKftwLhlg/5iJGSDMSdVfTUDSgTGSRQFQR
7+2db3VxbxlHjlQiAbK4Z9BLMvu5XQCXKvKpXppATqT2OSK5GsbZnmKw0uySOJFwlnTEc0NcFagw
KI0YZW/bvY+R09FNa9/umn8EAM/kV0k83nJ0XbppEZ7hYpyHyx0Rz5UaTBZC9Z10Tpn75TPhyYMi
YJwlsG5G5isKRJR6lH06CVC4EvM1ruGJPhu6z6VXvXyrOmTI2ksmqarXOr35+cglFvEP3G2/7VLb
WgPbau42oghdY+xCS8O1QdFvN1T0Qor5SNNasVL7KsdkLpCLkuxhht0a83ro40vgQlWI1ncL3lVQ
48f7QOIBAqVCDbUPKZmOxR7Jm4+mQBoYIvNwWLeDzxRc9Cdo/c4zii200A9zVhanAgmIA0C5sMRJ
LfEKBNTjFlWkQ++QJuMnfVtQR565rv3c8Z8KJmEChjQgaEVEV03Q9pAvTAXhI1No1mUlvhrQloXy
5812Hjp8PGAaontCZfLnde2Cfo6TwtxpW/N352e+C0cHohB2acm+W4nj7dbS9H6h/nFDEgAf7zaD
E33XYDn24GWeBAk26n3v7QCuT9a3+hDEKIiepuDeT9oNGWXYitLVBbvL4R2AWQ/AZUWJg0BV/OO4
jbyaAG5umtKpDx7gaORrf52XCqBpPIBQ8X18gb75i6DdCqfOg1vpR9ODZrXk9umGjaCWV1CgYW9H
oEntaxRl/Q4X4vh/pfYmY8yDOJl8I4YxQYna4030U/1PCpnYC4aNtXoCPYzSRcNbxkv5eRwd9ywr
tiumbTiaJa0QrTrx4SkiJlQ8HXWn+qF3idssXtOfcj7Jij0g9QTH4WtjPNHdWZ8xaF+46ih6jnyu
YEWgs2NgtnfR8o1t9XnVfa0xGwD+GIuZj8ZA8PDljTvq+cjpQcdJ6TtDp6/ZBLmIUy/+OAb85prr
/zojzH881JJ3azXeQ/OVpFE5TX+ye63ECcz/sCP67MacPSdh6YhJ9+KmU5BJmC9wBmes8kD8jmHS
MqmBzgwgm9vedQc9t56i7VuH26G2SCSt7D8YIOWeGH/8YQydrrcdqiucYEuaukowr4YbwoyP6+TV
bzono0nWzf40QcvVO8M23mwuktQyQUy8tvMEJmLdKIJwuwqr0vg9higyoV6mbEUJMHOAlXOyvQcD
0251faOjXvyd1mkvujP4BsRsgt5fII+v1/YwVuZc1D+mG5ABrdeGiS2jkH04OTYF67XBcOdJnhM0
jtzRG1l9SAQB4Mh/h9/v471i+3/GK0zDhXX4Ly6l3iIdceTgd5MSwGrOPDoExxDFirK+5+I3Txev
DKJAQYPnuaiOysfVLQSnY5BahlSps+rZtY24HuPRyZhqS4AowHhU7jTotI40RSfaYmavE1yCwOzy
q7FZdSfyuqGvsrmNlEj2e7O+hTor5jyTtKTkkZbVOcUwrVcUQLETAXG4rYPALdbNWVil4LZCVdLP
5OjAnNreVMaGpg4TKAdDZ+k6LHSleY7lTlFVWgKMApW0r7amEKJQ0EaSp19+G48/JFkF6Gq31q6r
7kZc+8X2KZXy/YzfVj2XhJb/a2X2Z9JDs+3Dl5plr3c4Fz1r+QnxPIxmoQ5BJuqFrX+zO7Z8FI4h
wBYTEMbWAZvUygOsqHFDQ+ds5Pjp38ZZ2hwBOJc5dOhdG+SyfEceIXuuaM9XqRpGmDAjkFzqZlpB
ENYCD2WbZfIW9vWir0Cp2fZtg6xoDDXNNzZF/1ELv+KPMapYdm73ERlj0qozKkkQNGy8ek0SY50S
DlOit+cTqccWWHHU2rlrgHWy1JsvGNc3sj0EOl/OdPff73ol2gZfqTdC8W2zfGwe9Vphg8EY1wbW
VB3vHm03vfa5ePwguqGLLFp+CBplYlGo3rHMp6sme7AdMBqbyKK9xYg/CFK1GMGZA7VfAvtxVSzM
bZMhAzGvO59MVeq1jmj9Jm8skiqfxZtN+WwFpgDT5W4+AR4w8jzG0ds0BRC5DMoACJ1iqw3yKAFO
t0A3dy1CZDeSwF5NAosQchP4X/d9vBWYRf1szybyjkwayQ8yjJwYYasVhKGd8fVw7TNVylZyZ5rX
CJvUaUPEv9b3shP/UdBUs1UEwHRetqol15OxQIxriMlRW8RVriNKMAui4TzFAGV/lS2v86dy7K+4
TUl0eeK2hW5vMdM8ssk03fY13wbmprb+Ouj47IRaTW5bUsK9ozTfDuIozKDh0e6/EapuIwRUY0IE
XQ6gSzxz1oP/NIVFeD3lEHuHk3mBnL7cLZAOeiMNDKI3XxnTupnlbVhhbchcHaXsItJQwkP1MFFX
p0CWHR5b9HV8OY+2PGQUlokhLXYIf49Mc5CGc4KXnChi4ZS3Km9anKJwVK5oUJgkTBVIj0kRZYXc
Agc/TD0ssQ==
`protect end_protected
